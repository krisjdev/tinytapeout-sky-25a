module tt_um_openfpga22 (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire net245;
 wire _0002_;
 wire net252;
 wire _0004_;
 wire net242;
 wire _0006_;
 wire net243;
 wire _0008_;
 wire net237;
 wire _0010_;
 wire net238;
 wire _0012_;
 wire net239;
 wire _0014_;
 wire net240;
 wire _0016_;
 wire net246;
 wire _0018_;
 wire net241;
 wire _0020_;
 wire net251;
 wire _0022_;
 wire net247;
 wire _0024_;
 wire net248;
 wire _0026_;
 wire net249;
 wire _0028_;
 wire net244;
 wire _0030_;
 wire net250;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire net253;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire net282;
 wire _0189_;
 wire _0190_;
 wire net276;
 wire _0192_;
 wire _0193_;
 wire net274;
 wire net332;
 wire net256;
 wire _0197_;
 wire _0198_;
 wire net272;
 wire net261;
 wire net366;
 wire _0202_;
 wire net378;
 wire net330;
 wire net422;
 wire net309;
 wire net392;
 wire net368;
 wire net338;
 wire net354;
 wire net417;
 wire net400;
 wire net323;
 wire net290;
 wire net292;
 wire net346;
 wire net266;
 wire net375;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire net409;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire net285;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire net286;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire net283;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire net284;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire net426;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire net299;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire net254;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire net280;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire net419;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire net302;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire net333;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire net403;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire net376;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire net420;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire net296;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire net421;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire net401;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire net423;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire net344;
 wire _0862_;
 wire net379;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire net313;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire net358;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire net359;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire net314;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire net360;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire net315;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire net319;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire net300;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire net343;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire net404;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire net428;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire net405;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire net380;
 wire _1229_;
 wire net393;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire net316;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire net361;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire net317;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire net362;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire net310;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire net355;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire net363;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire net311;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire net312;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire net356;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire net357;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire net406;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire net407;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire net427;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire clknet_0_net40;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.ccff_head ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.ccff_tail ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__0__1_ccff_tail ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.ccff_head ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.ccff_tail ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__1__1_ccff_tail ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.ccff_head ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.ccff_tail ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_0.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_3.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_4.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_5.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_6.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_7.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_ccff_tail ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.ccff_head ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.ccff_head ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.ccff_head ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_0__1_.ccff_head ;
 wire \dut_0.U0_formal_verification.cby_0__1_.ccff_tail ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_ccff_tail ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_0__2_.ccff_head ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__1_.ccff_tail ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__1__1_ccff_tail ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.ccff_tail ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_2.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_3.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_4.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_5.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_6.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_7.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_ccff_tail ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_ ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_0_ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.RST ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_0_ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \dut_0.U0_formal_verification.grid_io_top_1_ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.ccff_tail ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_right_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__0_.mem_top_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.ccff_head ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_14.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_right_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_0__2_.mem_right_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__0_.mem_top_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_left_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__0_.mem_top_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_left_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_3_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_2_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.D ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_17.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_0_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_1_.Q ;
 wire \dut_0.U0_formal_verification.sb_2__2_.mem_left_track_9.DFF_0_.Q ;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net234;
 wire net235;
 wire net236;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net255;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net273;
 wire net275;
 wire net277;
 wire net278;
 wire net279;
 wire net281;
 wire net287;
 wire net288;
 wire net289;
 wire net291;
 wire net293;
 wire net294;
 wire net295;
 wire net297;
 wire net298;
 wire net301;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net318;
 wire net320;
 wire net321;
 wire net322;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net331;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net345;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net364;
 wire net365;
 wire net367;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net377;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net402;
 wire net408;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net418;
 wire net424;
 wire net425;
 wire clknet_1_0__leaf_net40;
 wire clknet_1_1__leaf_net40;
 wire clknet_0_net39;
 wire clknet_1_0__leaf_net39;
 wire clknet_1_1__leaf_net39;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire clknet_0__0698_;
 wire clknet_1_0__leaf__0698_;
 wire clknet_1_1__leaf__0698_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire clknet_0__0757_;
 wire clknet_1_0__leaf__0757_;
 wire clknet_1_1__leaf__0757_;
 wire clknet_0__0820_;
 wire clknet_1_0__leaf__0820_;
 wire clknet_1_1__leaf__0820_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__1134_;
 wire clknet_1_0__leaf__1134_;
 wire clknet_1_1__leaf__1134_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0__1214_;
 wire clknet_1_0__leaf__1214_;
 wire clknet_1_1__leaf__1214_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire clknet_0_net50;
 wire clknet_1_0__leaf_net50;
 wire clknet_1_1__leaf_net50;
 wire clknet_0_net49;
 wire clknet_1_0__leaf_net49;
 wire clknet_1_1__leaf_net49;
 wire clknet_0__1199_;
 wire clknet_1_0__leaf__1199_;
 wire clknet_1_1__leaf__1199_;
 wire clknet_0__1178_;
 wire clknet_1_0__leaf__1178_;
 wire clknet_1_1__leaf__1178_;
 wire clknet_0__1149_;
 wire clknet_1_0__leaf__1149_;
 wire clknet_1_1__leaf__1149_;
 wire clknet_0__1118_;
 wire clknet_1_0__leaf__1118_;
 wire clknet_1_1__leaf__1118_;
 wire clknet_0__1108_;
 wire clknet_1_0__leaf__1108_;
 wire clknet_1_1__leaf__1108_;
 wire clknet_0__1563_;
 wire clknet_1_0__leaf__1563_;
 wire clknet_1_1__leaf__1563_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire clknet_0__1553_;
 wire clknet_1_0__leaf__1553_;
 wire clknet_1_1__leaf__1553_;
 wire clknet_0__1574_;
 wire clknet_1_0__leaf__1574_;
 wire clknet_1_1__leaf__1574_;
 wire clknet_0__1589_;
 wire clknet_1_0__leaf__1589_;
 wire clknet_1_1__leaf__1589_;
 wire clknet_0__1607_;
 wire clknet_1_0__leaf__1607_;
 wire clknet_1_1__leaf__1607_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0_net53;
 wire clknet_1_0__leaf_net53;
 wire clknet_1_1__leaf_net53;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire clknet_0__0527_;
 wire clknet_1_0__leaf__0527_;
 wire clknet_1_1__leaf__0527_;
 wire clknet_0__0529_;
 wire clknet_1_0__leaf__0529_;
 wire clknet_1_1__leaf__0529_;
 wire clknet_0__0532_;
 wire clknet_1_0__leaf__0532_;
 wire clknet_1_1__leaf__0532_;
 wire clknet_0__1168_;
 wire clknet_1_0__leaf__1168_;
 wire clknet_1_1__leaf__1168_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__1435_;
 wire clknet_1_0__leaf__1435_;
 wire clknet_1_1__leaf__1435_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0__1408_;
 wire clknet_1_0__leaf__1408_;
 wire clknet_1_1__leaf__1408_;
 wire clknet_0__1699_;
 wire clknet_1_0__leaf__1699_;
 wire clknet_1_1__leaf__1699_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0__1759_;
 wire clknet_1_0__leaf__1759_;
 wire clknet_1_1__leaf__1759_;
 wire clknet_0__1749_;
 wire clknet_1_0__leaf__1749_;
 wire clknet_1_1__leaf__1749_;
 wire clknet_0__0192_;
 wire clknet_1_0__leaf__0192_;
 wire clknet_1_1__leaf__0192_;
 wire clknet_0__1770_;
 wire clknet_1_0__leaf__1770_;
 wire clknet_1_1__leaf__1770_;
 wire clknet_0__1238_;
 wire clknet_1_0__leaf__1238_;
 wire clknet_1_1__leaf__1238_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire clknet_0__1393_;
 wire clknet_1_0__leaf__1393_;
 wire clknet_1_1__leaf__1393_;
 wire clknet_0__1395_;
 wire clknet_1_0__leaf__1395_;
 wire clknet_1_1__leaf__1395_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__1482_;
 wire clknet_1_0__leaf__1482_;
 wire clknet_1_1__leaf__1482_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0__1494_;
 wire clknet_1_0__leaf__1494_;
 wire clknet_1_1__leaf__1494_;
 wire clknet_0__1470_;
 wire clknet_1_0__leaf__1470_;
 wire clknet_1_1__leaf__1470_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0__1336_;
 wire clknet_1_0__leaf__1336_;
 wire clknet_1_1__leaf__1336_;
 wire clknet_0__1359_;
 wire clknet_1_0__leaf__1359_;
 wire clknet_1_1__leaf__1359_;
 wire clknet_0__1256_;
 wire clknet_1_0__leaf__1256_;
 wire clknet_1_1__leaf__1256_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0_net19;
 wire clknet_1_0__leaf_net19;
 wire clknet_1_1__leaf_net19;
 wire clknet_0__1420_;
 wire clknet_1_0__leaf__1420_;
 wire clknet_1_1__leaf__1420_;
 wire clknet_0_net18;
 wire clknet_1_0__leaf_net18;
 wire clknet_1_1__leaf_net18;
 wire clknet_0__1689_;
 wire clknet_1_0__leaf__1689_;
 wire clknet_1_1__leaf__1689_;
 wire clknet_0__1712_;
 wire clknet_1_0__leaf__1712_;
 wire clknet_1_1__leaf__1712_;
 wire clknet_0__1729_;
 wire clknet_1_0__leaf__1729_;
 wire clknet_1_1__leaf__1729_;
 wire clknet_0__0987_;
 wire clknet_1_0__leaf__0987_;
 wire clknet_1_1__leaf__0987_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0_net16;
 wire clknet_1_0__leaf_net16;
 wire clknet_1_1__leaf_net16;
 wire clknet_0__0534_;
 wire clknet_1_0__leaf__0534_;
 wire clknet_1_1__leaf__0534_;
 wire clknet_0__0539_;
 wire clknet_1_0__leaf__0539_;
 wire clknet_1_1__leaf__0539_;
 wire clknet_0__0558_;
 wire clknet_1_0__leaf__0558_;
 wire clknet_1_1__leaf__0558_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__1188_;
 wire clknet_1_0__leaf__1188_;
 wire clknet_1_1__leaf__1188_;
 wire clknet_0__1648_;
 wire clknet_1_0__leaf__1648_;
 wire clknet_1_1__leaf__1648_;
 wire clknet_0__1617_;
 wire clknet_1_0__leaf__1617_;
 wire clknet_1_1__leaf__1617_;
 wire clknet_0__1627_;
 wire clknet_1_0__leaf__1627_;
 wire clknet_1_1__leaf__1627_;
 wire clknet_0__1231_;
 wire clknet_1_0__leaf__1231_;
 wire clknet_1_1__leaf__1231_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire clknet_0__0849_;
 wire clknet_1_0__leaf__0849_;
 wire clknet_1_1__leaf__0849_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire clknet_0__1054_;
 wire clknet_1_0__leaf__1054_;
 wire clknet_1_1__leaf__1054_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ;
 wire clknet_0__0639_;
 wire clknet_1_0__leaf__0639_;
 wire clknet_1_1__leaf__0639_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__0642_;
 wire clknet_1_0__leaf__0642_;
 wire clknet_1_1__leaf__0642_;
 wire clknet_0__0646_;
 wire clknet_1_0__leaf__0646_;
 wire clknet_1_1__leaf__0646_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__0914_;
 wire clknet_1_0__leaf__0914_;
 wire clknet_1_1__leaf__0914_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire clknet_0__0524_;
 wire clknet_1_0__leaf__0524_;
 wire clknet_1_1__leaf__0524_;
 wire clknet_0__0526_;
 wire clknet_1_0__leaf__0526_;
 wire clknet_1_1__leaf__0526_;
 wire clknet_0__0528_;
 wire clknet_1_0__leaf__0528_;
 wire clknet_1_1__leaf__0528_;
 wire clknet_0__0611_;
 wire clknet_1_0__leaf__0611_;
 wire clknet_1_1__leaf__0611_;
 wire clknet_0__1072_;
 wire clknet_1_0__leaf__1072_;
 wire clknet_1_1__leaf__1072_;
 wire clknet_0__1077_;
 wire clknet_1_0__leaf__1077_;
 wire clknet_1_1__leaf__1077_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire clknet_0__0598_;
 wire clknet_1_0__leaf__0598_;
 wire clknet_1_1__leaf__0598_;
 wire clknet_0__0600_;
 wire clknet_1_0__leaf__0600_;
 wire clknet_1_1__leaf__0600_;
 wire clknet_0__0771_;
 wire clknet_1_0__leaf__0771_;
 wire clknet_1_1__leaf__0771_;
 wire clknet_0__0791_;
 wire clknet_1_0__leaf__0791_;
 wire clknet_1_1__leaf__0791_;
 wire clknet_0__0794_;
 wire clknet_1_0__leaf__0794_;
 wire clknet_1_1__leaf__0794_;
 wire clknet_0__0805_;
 wire clknet_1_0__leaf__0805_;
 wire clknet_1_1__leaf__0805_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire clknet_0__1346_;
 wire clknet_1_0__leaf__1346_;
 wire clknet_1_1__leaf__1346_;
 wire clknet_0__1280_;
 wire clknet_1_0__leaf__1280_;
 wire clknet_1_1__leaf__1280_;
 wire clknet_0__1266_;
 wire clknet_1_0__leaf__1266_;
 wire clknet_1_1__leaf__1266_;
 wire clknet_0__0938_;
 wire clknet_1_0__leaf__0938_;
 wire clknet_1_1__leaf__0938_;
 wire clknet_0__0924_;
 wire clknet_1_0__leaf__0924_;
 wire clknet_1_1__leaf__0924_;
 wire clknet_0__0879_;
 wire clknet_1_0__leaf__0879_;
 wire clknet_1_1__leaf__0879_;
 wire clknet_0__0881_;
 wire clknet_1_0__leaf__0881_;
 wire clknet_1_1__leaf__0881_;
 wire clknet_0__0883_;
 wire clknet_1_0__leaf__0883_;
 wire clknet_1_1__leaf__0883_;
 wire clknet_0__1091_;
 wire clknet_1_0__leaf__1091_;
 wire clknet_1_1__leaf__1091_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ;
 wire clknet_0__0744_;
 wire clknet_1_0__leaf__0744_;
 wire clknet_1_1__leaf__0744_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire clknet_0__0742_;
 wire clknet_1_0__leaf__0742_;
 wire clknet_1_1__leaf__0742_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ;
 wire clknet_0__0553_;
 wire clknet_1_0__leaf__0553_;
 wire clknet_1_1__leaf__0553_;
 wire clknet_0__0554_;
 wire clknet_1_0__leaf__0554_;
 wire clknet_1_1__leaf__0554_;
 wire clknet_0__0785_;
 wire clknet_1_0__leaf__0785_;
 wire clknet_1_1__leaf__0785_;
 wire clknet_0__0829_;
 wire clknet_1_0__leaf__0829_;
 wire clknet_1_1__leaf__0829_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__0831_;
 wire clknet_1_0__leaf__0831_;
 wire clknet_1_1__leaf__0831_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ;
 wire clknet_0__1049_;
 wire clknet_1_0__leaf__1049_;
 wire clknet_1_1__leaf__1049_;
 wire clknet_0__1061_;
 wire clknet_1_0__leaf__1061_;
 wire clknet_1_1__leaf__1061_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire clknet_0__0223_;
 wire clknet_1_0__leaf__0223_;
 wire clknet_1_1__leaf__0223_;
 wire clknet_0__0789_;
 wire clknet_1_0__leaf__0789_;
 wire clknet_1_1__leaf__0789_;
 wire clknet_0__0790_;
 wire clknet_1_0__leaf__0790_;
 wire clknet_1_1__leaf__0790_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire clknet_0__0895_;
 wire clknet_1_0__leaf__0895_;
 wire clknet_1_1__leaf__0895_;
 wire clknet_0__0897_;
 wire clknet_1_0__leaf__0897_;
 wire clknet_1_1__leaf__0897_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__0977_;
 wire clknet_1_0__leaf__0977_;
 wire clknet_1_1__leaf__0977_;
 wire clknet_0__1000_;
 wire clknet_1_0__leaf__1000_;
 wire clknet_1_1__leaf__1000_;
 wire clknet_0__1314_;
 wire clknet_1_0__leaf__1314_;
 wire clknet_1_1__leaf__1314_;
 wire clknet_0__1316_;
 wire clknet_1_0__leaf__1316_;
 wire clknet_1_1__leaf__1316_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ;
 wire clknet_0__0846_;
 wire clknet_1_0__leaf__0846_;
 wire clknet_1_1__leaf__0846_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__0723_;
 wire clknet_1_0__leaf__0723_;
 wire clknet_1_1__leaf__0723_;
 wire clknet_0_net33;
 wire clknet_1_0__leaf_net33;
 wire clknet_1_1__leaf_net33;
 wire clknet_0__1033_;
 wire clknet_1_0__leaf__1033_;
 wire clknet_1_1__leaf__1033_;
 wire clknet_0__1035_;
 wire clknet_1_0__leaf__1035_;
 wire clknet_1_1__leaf__1035_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__0445_;
 wire clknet_1_0__leaf__0445_;
 wire clknet_1_1__leaf__0445_;
 wire clknet_0__0426_;
 wire clknet_1_0__leaf__0426_;
 wire clknet_1_1__leaf__0426_;
 wire clknet_0__0378_;
 wire clknet_1_0__leaf__0378_;
 wire clknet_1_1__leaf__0378_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire clknet_0__0359_;
 wire clknet_1_0__leaf__0359_;
 wire clknet_1_1__leaf__0359_;
 wire clknet_0__0345_;
 wire clknet_1_0__leaf__0345_;
 wire clknet_1_1__leaf__0345_;
 wire clknet_0__0333_;
 wire clknet_1_0__leaf__0333_;
 wire clknet_1_1__leaf__0333_;
 wire clknet_0__0292_;
 wire clknet_1_0__leaf__0292_;
 wire clknet_1_1__leaf__0292_;
 wire clknet_0__0266_;
 wire clknet_1_0__leaf__0266_;
 wire clknet_1_1__leaf__0266_;
 wire clknet_0__0412_;
 wire clknet_1_0__leaf__0412_;
 wire clknet_1_1__leaf__0412_;
 wire clknet_0__0511_;
 wire clknet_1_0__leaf__0511_;
 wire clknet_1_1__leaf__0511_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ;
 wire clknet_0__0311_;
 wire clknet_1_0__leaf__0311_;
 wire clknet_1_1__leaf__0311_;
 wire clknet_0__0479_;
 wire clknet_1_0__leaf__0479_;
 wire clknet_1_1__leaf__0479_;
 wire clknet_0__0493_;
 wire clknet_1_0__leaf__0493_;
 wire clknet_1_1__leaf__0493_;
 wire clknet_0__0467_;
 wire clknet_1_0__leaf__0467_;
 wire clknet_1_1__leaf__0467_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__0868_;
 wire clknet_1_0__leaf__0868_;
 wire clknet_1_1__leaf__0868_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire clknet_0__0530_;
 wire clknet_1_0__leaf__0530_;
 wire clknet_1_1__leaf__0530_;
 wire clknet_0__0531_;
 wire clknet_1_0__leaf__0531_;
 wire clknet_1_1__leaf__0531_;
 wire clknet_0__0623_;
 wire clknet_1_0__leaf__0623_;
 wire clknet_1_1__leaf__0623_;
 wire clknet_0__0624_;
 wire clknet_1_0__leaf__0624_;
 wire clknet_1_1__leaf__0624_;
 wire clknet_0__0860_;
 wire clknet_1_0__leaf__0860_;
 wire clknet_1_1__leaf__0860_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__0633_;
 wire clknet_1_0__leaf__0633_;
 wire clknet_1_1__leaf__0633_;
 wire clknet_0__0634_;
 wire clknet_1_0__leaf__0634_;
 wire clknet_1_1__leaf__0634_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire clknet_0__0226_;
 wire clknet_1_0__leaf__0226_;
 wire clknet_1_1__leaf__0226_;
 wire clknet_0__0245_;
 wire clknet_1_0__leaf__0245_;
 wire clknet_1_1__leaf__0245_;
 wire clknet_0__0249_;
 wire clknet_1_0__leaf__0249_;
 wire clknet_1_1__leaf__0249_;
 wire clknet_0__0252_;
 wire clknet_1_0__leaf__0252_;
 wire clknet_1_1__leaf__0252_;
 wire clknet_0__0619_;
 wire clknet_1_0__leaf__0619_;
 wire clknet_1_1__leaf__0619_;
 wire clknet_0__0622_;
 wire clknet_1_0__leaf__0622_;
 wire clknet_1_1__leaf__0622_;
 wire clknet_0__0621_;
 wire clknet_1_0__leaf__0621_;
 wire clknet_1_1__leaf__0621_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ;
 wire clknet_0_net35;
 wire clknet_1_0__leaf_net35;
 wire clknet_1_1__leaf_net35;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire clknet_0__0246_;
 wire clknet_1_0__leaf__0246_;
 wire clknet_1_1__leaf__0246_;
 wire clknet_0__0248_;
 wire clknet_1_0__leaf__0248_;
 wire clknet_1_1__leaf__0248_;
 wire clknet_0__0602_;
 wire clknet_1_0__leaf__0602_;
 wire clknet_1_1__leaf__0602_;
 wire clknet_0__0613_;
 wire clknet_1_0__leaf__0613_;
 wire clknet_1_1__leaf__0613_;
 wire clknet_0__0603_;
 wire clknet_1_0__leaf__0603_;
 wire clknet_1_1__leaf__0603_;
 wire clknet_0__1102_;
 wire clknet_1_0__leaf__1102_;
 wire clknet_1_1__leaf__1102_;
 wire clknet_0_net22;
 wire clknet_1_0__leaf_net22;
 wire clknet_1_1__leaf_net22;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire clknet_0__0247_;
 wire clknet_1_0__leaf__0247_;
 wire clknet_1_1__leaf__0247_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire clknet_0__1095_;
 wire clknet_1_0__leaf__1095_;
 wire clknet_1_1__leaf__1095_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire clknet_0__0792_;
 wire clknet_1_0__leaf__0792_;
 wire clknet_1_1__leaf__0792_;
 wire clknet_0__0793_;
 wire clknet_1_0__leaf__0793_;
 wire clknet_1_1__leaf__0793_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ;
 wire clknet_0__0681_;
 wire clknet_1_0__leaf__0681_;
 wire clknet_1_1__leaf__0681_;
 wire clknet_0__0730_;
 wire clknet_1_0__leaf__0730_;
 wire clknet_1_1__leaf__0730_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire clknet_0__0250_;
 wire clknet_1_0__leaf__0250_;
 wire clknet_1_1__leaf__0250_;
 wire clknet_0__0251_;
 wire clknet_1_0__leaf__0251_;
 wire clknet_1_1__leaf__0251_;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ;
 wire clknet_0__0236_;
 wire clknet_1_0__leaf__0236_;
 wire clknet_1_1__leaf__0236_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire clknet_0__0738_;
 wire clknet_1_0__leaf__0738_;
 wire clknet_1_1__leaf__0738_;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ;
 wire clknet_0__0811_;
 wire clknet_1_0__leaf__0811_;
 wire clknet_1_1__leaf__0811_;
 wire clknet_0__0816_;
 wire clknet_1_0__leaf__0816_;
 wire clknet_1_1__leaf__0816_;
 wire clknet_0__0889_;
 wire clknet_1_0__leaf__0889_;
 wire clknet_1_1__leaf__0889_;
 wire clknet_0_net28;
 wire clknet_1_0__leaf_net28;
 wire clknet_1_1__leaf_net28;
 wire clknet_0_net27;
 wire clknet_1_0__leaf_net27;
 wire clknet_1_1__leaf_net27;
 wire clknet_0__0813_;
 wire clknet_1_0__leaf__0813_;
 wire clknet_1_1__leaf__0813_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ;
 wire clknet_0__0812_;
 wire clknet_1_0__leaf__0812_;
 wire clknet_1_1__leaf__0812_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire clknet_0__0592_;
 wire clknet_1_0__leaf__0592_;
 wire clknet_1_1__leaf__0592_;
 wire clknet_0__0594_;
 wire clknet_1_0__leaf__0594_;
 wire clknet_1_1__leaf__0594_;
 wire clknet_0__0597_;
 wire clknet_1_0__leaf__0597_;
 wire clknet_1_1__leaf__0597_;
 wire clknet_0__0599_;
 wire clknet_1_0__leaf__0599_;
 wire clknet_1_1__leaf__0599_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire clknet_0__0570_;
 wire clknet_1_0__leaf__0570_;
 wire clknet_1_1__leaf__0570_;
 wire clknet_0__0588_;
 wire clknet_1_0__leaf__0588_;
 wire clknet_1_1__leaf__0588_;
 wire clknet_0__0591_;
 wire clknet_1_0__leaf__0591_;
 wire clknet_1_1__leaf__0591_;
 wire clknet_0__0593_;
 wire clknet_1_0__leaf__0593_;
 wire clknet_1_1__leaf__0593_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire clknet_0__0650_;
 wire clknet_1_0__leaf__0650_;
 wire clknet_1_1__leaf__0650_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire clknet_0__0775_;
 wire clknet_1_0__leaf__0775_;
 wire clknet_1_1__leaf__0775_;
 wire clknet_0__0535_;
 wire clknet_1_0__leaf__0535_;
 wire clknet_1_1__leaf__0535_;
 wire clknet_0__0542_;
 wire clknet_1_0__leaf__0542_;
 wire clknet_1_1__leaf__0542_;
 wire clknet_0__0545_;
 wire clknet_1_0__leaf__0545_;
 wire clknet_1_1__leaf__0545_;
 wire clknet_0__0548_;
 wire clknet_1_0__leaf__0548_;
 wire clknet_1_1__leaf__0548_;
 wire clknet_0__0551_;
 wire clknet_1_0__leaf__0551_;
 wire clknet_1_1__leaf__0551_;
 wire clknet_0__0555_;
 wire clknet_1_0__leaf__0555_;
 wire clknet_1_1__leaf__0555_;
 wire clknet_0__0550_;
 wire clknet_1_0__leaf__0550_;
 wire clknet_1_1__leaf__0550_;
 wire clknet_0__0702_;
 wire clknet_1_0__leaf__0702_;
 wire clknet_1_1__leaf__0702_;
 wire clknet_0__0704_;
 wire clknet_1_0__leaf__0704_;
 wire clknet_1_1__leaf__0704_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire clknet_0__0665_;
 wire clknet_1_0__leaf__0665_;
 wire clknet_1_1__leaf__0665_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire clknet_0__0667_;
 wire clknet_1_0__leaf__0667_;
 wire clknet_1_1__leaf__0667_;
 wire clknet_0__0669_;
 wire clknet_1_0__leaf__0669_;
 wire clknet_1_1__leaf__0669_;
 wire clknet_0__0795_;
 wire clknet_1_0__leaf__0795_;
 wire clknet_1_1__leaf__0795_;
 wire clknet_0__0796_;
 wire clknet_1_0__leaf__0796_;
 wire clknet_1_1__leaf__0796_;
 wire clknet_0__0671_;
 wire clknet_1_0__leaf__0671_;
 wire clknet_1_1__leaf__0671_;
 wire clknet_0__0675_;
 wire clknet_1_0__leaf__0675_;
 wire clknet_1_1__leaf__0675_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire clknet_0__0668_;
 wire clknet_1_0__leaf__0668_;
 wire clknet_1_1__leaf__0668_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire clknet_0__0567_;
 wire clknet_1_0__leaf__0567_;
 wire clknet_1_1__leaf__0567_;
 wire clknet_0__0569_;
 wire clknet_1_0__leaf__0569_;
 wire clknet_1_1__leaf__0569_;
 wire clknet_0__0572_;
 wire clknet_1_0__leaf__0572_;
 wire clknet_1_1__leaf__0572_;
 wire clknet_0__0574_;
 wire clknet_1_0__leaf__0574_;
 wire clknet_1_1__leaf__0574_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire clknet_0__0571_;
 wire clknet_1_0__leaf__0571_;
 wire clknet_1_1__leaf__0571_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire clknet_0__0546_;
 wire clknet_1_0__leaf__0546_;
 wire clknet_1_1__leaf__0546_;
 wire clknet_0__0547_;
 wire clknet_1_0__leaf__0547_;
 wire clknet_1_1__leaf__0547_;
 wire clknet_0__0568_;
 wire clknet_1_0__leaf__0568_;
 wire clknet_1_1__leaf__0568_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire clknet_0__0230_;
 wire clknet_1_0__leaf__0230_;
 wire clknet_1_1__leaf__0230_;
 wire clknet_0__0255_;
 wire clknet_1_0__leaf__0255_;
 wire clknet_1_1__leaf__0255_;
 wire clknet_0__0523_;
 wire clknet_1_0__leaf__0523_;
 wire clknet_1_1__leaf__0523_;
 wire clknet_0__0525_;
 wire clknet_1_0__leaf__0525_;
 wire clknet_1_1__leaf__0525_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire clknet_0__0543_;
 wire clknet_1_0__leaf__0543_;
 wire clknet_1_1__leaf__0543_;
 wire clknet_0__0544_;
 wire clknet_1_0__leaf__0544_;
 wire clknet_1_1__leaf__0544_;
 wire clknet_0__0688_;
 wire clknet_1_0__leaf__0688_;
 wire clknet_1_1__leaf__0688_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ;
 wire clknet_0__0764_;
 wire clknet_1_0__leaf__0764_;
 wire clknet_1_1__leaf__0764_;
 wire clknet_0__0766_;
 wire clknet_1_0__leaf__0766_;
 wire clknet_1_1__leaf__0766_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ;
 wire clknet_0__0578_;
 wire clknet_1_0__leaf__0578_;
 wire clknet_1_1__leaf__0578_;
 wire clknet_0__0677_;
 wire clknet_1_0__leaf__0677_;
 wire clknet_1_1__leaf__0677_;
 wire clknet_0__0700_;
 wire clknet_1_0__leaf__0700_;
 wire clknet_1_1__leaf__0700_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__0679_;
 wire clknet_1_0__leaf__0679_;
 wire clknet_1_1__leaf__0679_;
 wire clknet_0__0714_;
 wire clknet_1_0__leaf__0714_;
 wire clknet_1_1__leaf__0714_;
 wire clknet_0__0718_;
 wire clknet_1_0__leaf__0718_;
 wire clknet_1_1__leaf__0718_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire clknet_0__0256_;
 wire clknet_1_0__leaf__0256_;
 wire clknet_1_1__leaf__0256_;
 wire clknet_0__0257_;
 wire clknet_1_0__leaf__0257_;
 wire clknet_1_1__leaf__0257_;
 wire clknet_0__0259_;
 wire clknet_1_0__leaf__0259_;
 wire clknet_1_1__leaf__0259_;
 wire clknet_0__0261_;
 wire clknet_1_0__leaf__0261_;
 wire clknet_1_1__leaf__0261_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ;
 wire clknet_0__0653_;
 wire clknet_1_0__leaf__0653_;
 wire clknet_1_1__leaf__0653_;
 wire clknet_0__0655_;
 wire clknet_1_0__leaf__0655_;
 wire clknet_1_1__leaf__0655_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire clknet_0__0626_;
 wire clknet_1_0__leaf__0626_;
 wire clknet_1_1__leaf__0626_;
 wire clknet_0__0628_;
 wire clknet_1_0__leaf__0628_;
 wire clknet_1_1__leaf__0628_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ;
 wire clknet_0__0648_;
 wire clknet_1_0__leaf__0648_;
 wire clknet_1_1__leaf__0648_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire clknet_0__0253_;
 wire clknet_1_0__leaf__0253_;
 wire clknet_1_1__leaf__0253_;
 wire clknet_0__0254_;
 wire clknet_1_0__leaf__0254_;
 wire clknet_1_1__leaf__0254_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire clknet_0__0661_;
 wire clknet_1_0__leaf__0661_;
 wire clknet_1_1__leaf__0661_;
 wire clknet_0__0899_;
 wire clknet_1_0__leaf__0899_;
 wire clknet_1_1__leaf__0899_;
 wire clknet_0__0901_;
 wire clknet_1_0__leaf__0901_;
 wire clknet_1_1__leaf__0901_;
 wire clknet_0__0900_;
 wire clknet_1_0__leaf__0900_;
 wire clknet_1_1__leaf__0900_;
 wire clknet_0__0663_;
 wire clknet_1_0__leaf__0663_;
 wire clknet_1_1__leaf__0663_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire clknet_0__0709_;
 wire clknet_1_0__leaf__0709_;
 wire clknet_1_1__leaf__0709_;
 wire clknet_0__0710_;
 wire clknet_1_0__leaf__0710_;
 wire clknet_1_1__leaf__0710_;
 wire clknet_0__0711_;
 wire clknet_1_0__leaf__0711_;
 wire clknet_1_1__leaf__0711_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ;
 wire clknet_0__0219_;
 wire clknet_1_0__leaf__0219_;
 wire clknet_1_1__leaf__0219_;
 wire clknet_0__0222_;
 wire clknet_1_0__leaf__0222_;
 wire clknet_1_1__leaf__0222_;
 wire clknet_0__0225_;
 wire clknet_1_0__leaf__0225_;
 wire clknet_1_1__leaf__0225_;
 wire clknet_0__0228_;
 wire clknet_1_0__leaf__0228_;
 wire clknet_1_1__leaf__0228_;
 wire clknet_0__0233_;
 wire clknet_1_0__leaf__0233_;
 wire clknet_1_1__leaf__0233_;
 wire clknet_0__0227_;
 wire clknet_1_0__leaf__0227_;
 wire clknet_1_1__leaf__0227_;
 wire clknet_0__0224_;
 wire clknet_1_0__leaf__0224_;
 wire clknet_1_1__leaf__0224_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire clknet_0__0563_;
 wire clknet_1_0__leaf__0563_;
 wire clknet_1_1__leaf__0563_;
 wire clknet_0__0566_;
 wire clknet_1_0__leaf__0566_;
 wire clknet_1_1__leaf__0566_;
 wire clknet_0__0565_;
 wire clknet_1_0__leaf__0565_;
 wire clknet_1_1__leaf__0565_;
 wire clknet_0__0564_;
 wire clknet_1_0__leaf__0564_;
 wire clknet_1_1__leaf__0564_;
 wire clknet_0__0221_;
 wire clknet_1_0__leaf__0221_;
 wire clknet_1_1__leaf__0221_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ;
 wire clknet_0__0559_;
 wire clknet_1_0__leaf__0559_;
 wire clknet_1_1__leaf__0559_;
 wire clknet_0__0562_;
 wire clknet_1_0__leaf__0562_;
 wire clknet_1_1__leaf__0562_;
 wire clknet_0__0561_;
 wire clknet_1_0__leaf__0561_;
 wire clknet_1_1__leaf__0561_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ;
 wire clknet_0__0607_;
 wire clknet_1_0__leaf__0607_;
 wire clknet_1_1__leaf__0607_;
 wire clknet_0__0609_;
 wire clknet_1_0__leaf__0609_;
 wire clknet_1_1__leaf__0609_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ;
 wire clknet_0__0589_;
 wire clknet_1_0__leaf__0589_;
 wire clknet_1_1__leaf__0589_;
 wire clknet_0__0590_;
 wire clknet_1_0__leaf__0590_;
 wire clknet_1_1__leaf__0590_;
 wire clknet_0__0232_;
 wire clknet_1_0__leaf__0232_;
 wire clknet_1_1__leaf__0232_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ;
 wire clknet_0__0620_;
 wire clknet_1_0__leaf__0620_;
 wire clknet_1_1__leaf__0620_;
 wire clknet_0__0537_;
 wire clknet_1_0__leaf__0537_;
 wire clknet_1_1__leaf__0537_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ;
 wire clknet_0__0596_;
 wire clknet_1_0__leaf__0596_;
 wire clknet_1_1__leaf__0596_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ;
 wire clknet_0__0595_;
 wire clknet_1_0__leaf__0595_;
 wire clknet_1_1__leaf__0595_;
 wire \clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ;
 wire clknet_0__0231_;
 wire clknet_1_0__leaf__0231_;
 wire clknet_1_1__leaf__0231_;
 wire \clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ;
 wire clknet_0__0560_;
 wire clknet_1_0__leaf__0560_;
 wire clknet_1_1__leaf__0560_;
 wire clknet_0__0536_;
 wire clknet_1_0__leaf__0536_;
 wire clknet_1_1__leaf__0536_;
 wire clknet_0__0202_;
 wire clknet_1_0__leaf__0202_;
 wire clknet_1_1__leaf__0202_;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__0197_;
 wire clknet_1_0__leaf__0197_;
 wire clknet_1_1__leaf__0197_;
 wire clknet_0__0586_;
 wire clknet_1_0__leaf__0586_;
 wire clknet_1_1__leaf__0586_;
 wire clknet_0__0549_;
 wire clknet_1_0__leaf__0549_;
 wire clknet_1_1__leaf__0549_;
 wire clknet_0__0615_;
 wire clknet_1_0__leaf__0615_;
 wire clknet_1_1__leaf__0615_;
 wire clknet_0__0617_;
 wire clknet_1_0__leaf__0617_;
 wire clknet_1_1__leaf__0617_;
 wire clknet_0__0193_;
 wire clknet_1_0__leaf__0193_;
 wire clknet_1_1__leaf__0193_;
 wire clknet_0_net31;
 wire clknet_1_0__leaf_net31;
 wire clknet_1_1__leaf_net31;
 wire clknet_0_net29;
 wire clknet_1_0__leaf_net29;
 wire clknet_1_1__leaf_net29;
 wire clknet_0_net23;
 wire clknet_1_0__leaf_net23;
 wire clknet_1_1__leaf_net23;
 wire \clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire clknet_0__0220_;
 wire clknet_1_0__leaf__0220_;
 wire clknet_1_1__leaf__0220_;
 wire clknet_0_net52;
 wire clknet_1_0__leaf_net52;
 wire clknet_1_1__leaf_net52;

 sky130_fd_sc_hd__o21a_2 _2173_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_0_.Q ),
    .A2(net377),
    .B1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1800_));
 sky130_fd_sc_hd__o21ai_2 _2174_ (.A1(_0138_),
    .A2(clknet_1_0__leaf__0675_),
    .B1(_1800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_1 _2175_ (.A1(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(net279),
    .B1(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1801_));
 sky130_fd_sc_hd__a21o_1 _2176_ (.A1(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(net38),
    .B1(_1801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _2177_ (.A0(clknet_1_1__leaf__0596_),
    .A1(clknet_1_1__leaf__1238_),
    .S(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1802_));
 sky130_fd_sc_hd__nand2_2 _2178_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_1_.Q ),
    .B(_1802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _2179_ (.A0(net353),
    .A1(clknet_1_0__leaf__0879_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1803_));
 sky130_fd_sc_hd__nand2_2 _2180_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_1_.Q ),
    .B(_1803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o211a_2 _2181_ (.A1(_0139_),
    .A2(clknet_1_1__leaf__0785_),
    .B1(_0140_),
    .C1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1804_));
 sky130_fd_sc_hd__a21bo_2 _2182_ (.A1(_0139_),
    .A2(clknet_1_1__leaf__0650_),
    .B1_N(_1804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1805_));
 sky130_fd_sc_hd__nand2_1 _2183_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1806_));
 sky130_fd_sc_hd__o211a_1 _2184_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .B1(_1806_),
    .C1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1807_));
 sky130_fd_sc_hd__a21oi_2 _2185_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0805_),
    .B1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1808_));
 sky130_fd_sc_hd__o21a_2 _2186_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0704_),
    .B1(_1808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1809_));
 sky130_fd_sc_hd__o31a_1 _2187_ (.A1(_0140_),
    .A2(_1807_),
    .A3(_1809_),
    .B1(_1805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(clknet_1_1__leaf__0796_),
    .A1(clknet_1_0__leaf__1049_),
    .S(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1810_));
 sky130_fd_sc_hd__or3b_2 _2189_ (.A(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_2_.Q ),
    .B(_1810_),
    .C_N(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1811_));
 sky130_fd_sc_hd__mux4_2 _2190_ (.A0(clknet_1_1__leaf__0233_),
    .A1(clknet_1_0__leaf__0846_),
    .A2(net365),
    .A3(clknet_1_0__leaf__1072_),
    .S0(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1812_));
 sky130_fd_sc_hd__a21boi_2 _2191_ (.A1(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_2_.Q ),
    .A2(_1812_),
    .B1_N(_1811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _2192_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1813_));
 sky130_fd_sc_hd__o2111a_2 _2193_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0881_),
    .B1(_1813_),
    .C1(_0144_),
    .D1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1814_));
 sky130_fd_sc_hd__a21bo_2 _2194_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0550_),
    .B1_N(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1815_));
 sky130_fd_sc_hd__a21o_2 _2195_ (.A1(_0143_),
    .A2(clknet_1_0__leaf__0897_),
    .B1(_1815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1816_));
 sky130_fd_sc_hd__nor2_2 _2196_ (.A(_0143_),
    .B(clknet_1_0__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1817_));
 sky130_fd_sc_hd__a211o_2 _2197_ (.A1(_0143_),
    .A2(clknet_1_0__leaf__0793_),
    .B1(_1817_),
    .C1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1818_));
 sky130_fd_sc_hd__a31oi_2 _2198_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_2_.Q ),
    .A2(_1816_),
    .A3(_1818_),
    .B1(_1814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _2199_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1819_));
 sky130_fd_sc_hd__o2111a_2 _2200_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0534_),
    .B1(_1819_),
    .C1(_0145_),
    .D1(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1820_));
 sky130_fd_sc_hd__mux2_1 _2201_ (.A0(clknet_1_1__leaf__0626_),
    .A1(clknet_1_1__leaf__0564_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(clknet_1_0__leaf__0653_),
    .A1(clknet_1_1__leaf__0224_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(_1822_),
    .A1(_1821_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1823_));
 sky130_fd_sc_hd__a21oi_4 _2204_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_2_.Q ),
    .A2(_1823_),
    .B1(_1820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _2205_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1824_));
 sky130_fd_sc_hd__mux4_2 _2206_ (.A0(net329),
    .A1(net291),
    .A2(net265),
    .A3(net289),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1825_));
 sky130_fd_sc_hd__o211a_1 _2207_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_0_.Q ),
    .A2(clknet_1_1__leaf_net35),
    .B1(_1824_),
    .C1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1826_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(_1826_),
    .A1(_1825_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2209_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1827_));
 sky130_fd_sc_hd__nand2_1 _2210_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1828_));
 sky130_fd_sc_hd__o2111a_1 _2211_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0757_),
    .B1(_1828_),
    .C1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_1_.Q ),
    .D1(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1829_));
 sky130_fd_sc_hd__o21bai_1 _2212_ (.A1(_0161_),
    .A2(_1827_),
    .B1_N(_1829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2_1 _2213_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1830_));
 sky130_fd_sc_hd__o2111a_1 _2214_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0757_),
    .B1(_1830_),
    .C1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_1_.Q ),
    .D1(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(clknet_1_1__leaf__0571_),
    .A1(clknet_1_0__leaf__0711_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_1 _2216_ (.A0(clknet_1_0__leaf__0247_),
    .A1(clknet_1_1__leaf__0663_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _2217_ (.A0(_1832_),
    .A1(_1833_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1834_));
 sky130_fd_sc_hd__a21o_1 _2218_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_2_.Q ),
    .A2(_1834_),
    .B1(_1831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2219_ (.A0(net271),
    .A1(net337),
    .A2(clknet_1_0__leaf__0547_),
    .A3(clknet_1_0__leaf__0528_),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1835_));
 sky130_fd_sc_hd__and2b_1 _2220_ (.A_N(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _2221_ (.A0(clknet_1_1__leaf__0571_),
    .A1(clknet_1_1__leaf__0711_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1837_));
 sky130_fd_sc_hd__a22o_1 _2222_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_2_.Q ),
    .A2(_1835_),
    .B1(_1836_),
    .B2(_1837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2223_ (.A0(clknet_1_1__leaf_net35),
    .A1(net260),
    .A2(net328),
    .A3(net264),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1838_));
 sky130_fd_sc_hd__and2b_1 _2224_ (.A_N(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _2225_ (.A0(net270),
    .A1(clknet_1_0__leaf__0547_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1840_));
 sky130_fd_sc_hd__a22o_2 _2226_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_2_.Q ),
    .A2(_1838_),
    .B1(_1839_),
    .B2(_1840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2227_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1841_));
 sky130_fd_sc_hd__o21ai_1 _2228_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf_net35),
    .B1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1842_));
 sky130_fd_sc_hd__a211o_2 _2229_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .B1(_1842_),
    .C1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1843_));
 sky130_fd_sc_hd__o21ai_2 _2230_ (.A1(_0163_),
    .A2(_1841_),
    .B1(_1843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2_1 _2231_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1844_));
 sky130_fd_sc_hd__o2111a_1 _2232_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0757_),
    .B1(_1844_),
    .C1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_1_.Q ),
    .D1(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1845_));
 sky130_fd_sc_hd__mux4_2 _2233_ (.A0(net345),
    .A1(clknet_1_0__leaf__0247_),
    .A2(net331),
    .A3(clknet_1_0__leaf__0663_),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1846_));
 sky130_fd_sc_hd__a21o_1 _2234_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_2_.Q ),
    .A2(_1846_),
    .B1(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2235_ (.A0(clknet_1_0__leaf__0247_),
    .A1(clknet_1_0__leaf__0663_),
    .A2(net336),
    .A3(clknet_1_0__leaf__0528_),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1847_));
 sky130_fd_sc_hd__and2b_1 _2236_ (.A_N(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_1 _2237_ (.A0(clknet_1_0__leaf__0571_),
    .A1(clknet_1_0__leaf__0711_),
    .S(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1849_));
 sky130_fd_sc_hd__a22o_1 _2238_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_2_.Q ),
    .A2(_1847_),
    .B1(_1848_),
    .B2(_1849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2239_ (.A0(net335),
    .A1(net288),
    .A2(net327),
    .A3(clknet_1_0__leaf__0868_),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1850_));
 sky130_fd_sc_hd__or2_1 _2240_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_0_.Q ),
    .B(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1851_));
 sky130_fd_sc_hd__a21oi_2 _2241_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .B1(\dut_0.U0_formal_verification.cbx_1__0__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1852_));
 sky130_fd_sc_hd__a32o_2 _2242_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_1_.Q ),
    .A2(_1851_),
    .A3(_1852_),
    .B1(\dut_0.U0_formal_verification.cbx_1__0__1_ccff_tail ),
    .B2(_1850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2243_ (.A0(clknet_1_1__leaf_net35),
    .A1(net326),
    .A2(clknet_1_1__leaf__1095_),
    .A3(clknet_1_0__leaf__0868_),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1853_));
 sky130_fd_sc_hd__nand2_2 _2244_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1854_));
 sky130_fd_sc_hd__o211a_2 _2245_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0599_),
    .B1(_0165_),
    .C1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1855_));
 sky130_fd_sc_hd__a22o_2 _2246_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_2_.Q ),
    .A2(_1853_),
    .B1(_1854_),
    .B2(_1855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2_2 _2247_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1856_));
 sky130_fd_sc_hd__o211a_2 _2248_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0599_),
    .B1(_0166_),
    .C1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1857_));
 sky130_fd_sc_hd__mux4_2 _2249_ (.A0(clknet_1_1__leaf__0671_),
    .A1(clknet_1_0__leaf__0714_),
    .A2(clknet_1_1__leaf__0547_),
    .A3(clknet_1_1__leaf__0528_),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1858_));
 sky130_fd_sc_hd__a22o_2 _2250_ (.A1(_1856_),
    .A2(_1857_),
    .B1(_1858_),
    .B2(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2251_ (.A0(clknet_1_0__leaf__0572_),
    .A1(clknet_1_1__leaf__0248_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1859_));
 sky130_fd_sc_hd__nor2_1 _2252_ (.A(_0167_),
    .B(_1859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1860_));
 sky130_fd_sc_hd__mux2_1 _2253_ (.A0(clknet_1_0__leaf__0671_),
    .A1(clknet_1_0__leaf__0547_),
    .S(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1861_));
 sky130_fd_sc_hd__a31o_1 _2254_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_1_.Q ),
    .A2(_0167_),
    .A3(_1861_),
    .B1(_1860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2255_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1862_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(clknet_1_1__leaf__0572_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .S(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1863_));
 sky130_fd_sc_hd__or3b_2 _2257_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_2_.Q ),
    .B(_1863_),
    .C_N(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1864_));
 sky130_fd_sc_hd__o21ai_1 _2258_ (.A1(_0168_),
    .A2(_1862_),
    .B1(_1864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2259_ (.A0(clknet_1_1__leaf_net35),
    .A1(net325),
    .A2(clknet_1_1__leaf__1095_),
    .A3(clknet_1_0__leaf__0868_),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1865_));
 sky130_fd_sc_hd__nand2_2 _2260_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1866_));
 sky130_fd_sc_hd__o211a_2 _2261_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(net268),
    .B1(_1866_),
    .C1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_1 _2262_ (.A0(_1867_),
    .A1(_1865_),
    .S(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2_2 _2263_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1868_));
 sky130_fd_sc_hd__o211a_2 _2264_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0599_),
    .B1(_0169_),
    .C1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1869_));
 sky130_fd_sc_hd__mux4_2 _2265_ (.A0(clknet_1_1__leaf_net35),
    .A1(clknet_1_1__leaf__0714_),
    .A2(clknet_1_1__leaf__1095_),
    .A3(clknet_1_1__leaf__0528_),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1870_));
 sky130_fd_sc_hd__a22o_2 _2266_ (.A1(_1868_),
    .A2(_1869_),
    .B1(_1870_),
    .B2(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ ));
 sky130_fd_sc_hd__and2b_1 _2267_ (.A_N(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1871_));
 sky130_fd_sc_hd__mux2_1 _2268_ (.A0(clknet_1_1__leaf__0671_),
    .A1(clknet_1_1__leaf__0547_),
    .S(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1872_));
 sky130_fd_sc_hd__mux4_2 _2269_ (.A0(clknet_1_1__leaf__0714_),
    .A1(clknet_1_1__leaf__0528_),
    .A2(clknet_1_1__leaf__0247_),
    .A3(net263),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1873_));
 sky130_fd_sc_hd__a22o_2 _2270_ (.A1(_1871_),
    .A2(_1872_),
    .B1(_1873_),
    .B2(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2271_ (.A0(net308),
    .A1(net416),
    .A2(clknet_1_0__leaf__0224_),
    .A3(clknet_1_0__leaf__0564_),
    .S0(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1874_));
 sky130_fd_sc_hd__and2b_1 _2272_ (.A_N(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1875_));
 sky130_fd_sc_hd__mux2_1 _2273_ (.A0(clknet_1_0__leaf__0257_),
    .A1(clknet_1_0__leaf__1316_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1876_));
 sky130_fd_sc_hd__a22o_1 _2274_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_2_.Q ),
    .A2(_1874_),
    .B1(_1875_),
    .B2(_1876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_7.out ));
 sky130_fd_sc_hd__mux2_1 _2275_ (.A0(net307),
    .A1(clknet_1_0__leaf__0224_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1877_));
 sky130_fd_sc_hd__mux2_1 _2276_ (.A0(clknet_1_0__leaf__0702_),
    .A1(clknet_1_0__leaf__0677_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1878_));
 sky130_fd_sc_hd__o21ai_2 _2277_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .B1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1879_));
 sky130_fd_sc_hd__a21o_2 _2278_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0665_),
    .B1(_1879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1880_));
 sky130_fd_sc_hd__o211a_1 _2279_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .A2(_1878_),
    .B1(_1880_),
    .C1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1881_));
 sky130_fd_sc_hd__a31o_1 _2280_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .A2(_0170_),
    .A3(_1877_),
    .B1(_1881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_6.out ));
 sky130_fd_sc_hd__mux4_1 _2281_ (.A0(clknet_1_0__leaf__1393_),
    .A1(clknet_1_0__leaf__0829_),
    .A2(clknet_1_0__leaf__0254_),
    .A3(clknet_1_0__leaf__0593_),
    .S0(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _2282_ (.A0(clknet_1_0__leaf__0702_),
    .A1(clknet_1_0__leaf__0677_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1883_));
 sky130_fd_sc_hd__and3b_1 _2283_ (.A_N(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_2_.Q ),
    .B(_1883_),
    .C(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1884_));
 sky130_fd_sc_hd__a21o_1 _2284_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_2_.Q ),
    .A2(_1882_),
    .B1(_1884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_5.out ));
 sky130_fd_sc_hd__mux4_1 _2285_ (.A0(clknet_1_0__leaf__0537_),
    .A1(clknet_1_0__leaf__1393_),
    .A2(clknet_1_0__leaf__0648_),
    .A3(clknet_1_0__leaf__0254_),
    .S0(_0171_),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1885_));
 sky130_fd_sc_hd__nor2_2 _2286_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1886_));
 sky130_fd_sc_hd__a211o_2 _2287_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__1035_),
    .B1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_2_.Q ),
    .C1(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1887_));
 sky130_fd_sc_hd__a2bb2o_1 _2288_ (.A1_N(_1886_),
    .A2_N(_1887_),
    .B1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_2_.Q ),
    .B2(_1885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_4.out ));
 sky130_fd_sc_hd__mux4_2 _2289_ (.A0(clknet_1_0__leaf__0537_),
    .A1(clknet_1_1__leaf__0648_),
    .A2(net415),
    .A3(clknet_1_0__leaf__0564_),
    .S0(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1888_));
 sky130_fd_sc_hd__and2b_1 _2290_ (.A_N(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1889_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(clknet_1_0__leaf__0257_),
    .A1(clknet_1_1__leaf__1316_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1890_));
 sky130_fd_sc_hd__a22o_1 _2292_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .A2(_1888_),
    .B1(_1889_),
    .B2(_1890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_3.out ));
 sky130_fd_sc_hd__mux4_2 _2293_ (.A0(net414),
    .A1(clknet_1_0__leaf__0564_),
    .A2(net352),
    .A3(clknet_1_0__leaf__0665_),
    .S0(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1891_));
 sky130_fd_sc_hd__and2b_1 _2294_ (.A_N(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1892_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(net306),
    .A1(clknet_1_0__leaf__0224_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1893_));
 sky130_fd_sc_hd__a22o_2 _2296_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_2_.Q ),
    .A2(_1891_),
    .B1(_1892_),
    .B2(_1893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.out ));
 sky130_fd_sc_hd__mux4_2 _2297_ (.A0(net351),
    .A1(clknet_1_0__leaf__0665_),
    .A2(clknet_1_0__leaf__0829_),
    .A3(clknet_1_0__leaf__0593_),
    .S0(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _2298_ (.A0(clknet_1_0__leaf__0702_),
    .A1(clknet_1_0__leaf__0677_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1895_));
 sky130_fd_sc_hd__and3b_1 _2299_ (.A_N(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_2_.Q ),
    .B(_1895_),
    .C(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1896_));
 sky130_fd_sc_hd__a21o_1 _2300_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_2_.Q ),
    .A2(_1894_),
    .B1(_1896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.out ));
 sky130_fd_sc_hd__mux4_2 _2301_ (.A0(clknet_1_1__leaf__1393_),
    .A1(clknet_1_0__leaf__0829_),
    .A2(clknet_1_0__leaf__0254_),
    .A3(clknet_1_0__leaf__0593_),
    .S0(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1897_));
 sky130_fd_sc_hd__nand2_2 _2302_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1898_));
 sky130_fd_sc_hd__o2111a_2 _2303_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0811_),
    .B1(_1898_),
    .C1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_1_.Q ),
    .D1(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1899_));
 sky130_fd_sc_hd__a21o_2 _2304_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_2_.Q ),
    .A2(_1897_),
    .B1(_1899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_0.out ));
 sky130_fd_sc_hd__nand2b_1 _2305_ (.A_N(clknet_1_1__leaf__0677_),
    .B(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1900_));
 sky130_fd_sc_hd__mux4_2 _2306_ (.A0(clknet_1_1__leaf__0653_),
    .A1(clknet_1_1__leaf__0537_),
    .A2(clknet_1_1__leaf__0224_),
    .A3(clknet_1_1__leaf__0665_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1901_));
 sky130_fd_sc_hd__o211a_2 _2307_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0257_),
    .B1(_1900_),
    .C1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1902_));
 sky130_fd_sc_hd__mux2_1 _2308_ (.A0(_1902_),
    .A1(_1901_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2309_ (.A0(net305),
    .A1(net413),
    .A2(clknet_1_0__leaf__0254_),
    .A3(clknet_1_0__leaf__0593_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1903_));
 sky130_fd_sc_hd__nand2b_1 _2310_ (.A_N(clknet_1_0__leaf__0677_),
    .B(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1904_));
 sky130_fd_sc_hd__o211a_2 _2311_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0257_),
    .B1(_1904_),
    .C1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _2312_ (.A0(_1905_),
    .A1(_1903_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2313_ (.A0(clknet_1_1__leaf__0702_),
    .A1(clknet_1_0__leaf__0895_),
    .A2(net350),
    .A3(clknet_1_0__leaf__0879_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _2314_ (.A0(net304),
    .A1(clknet_1_1__leaf__0254_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1907_));
 sky130_fd_sc_hd__and3b_2 _2315_ (.A_N(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_2_.Q ),
    .B(_1907_),
    .C(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1908_));
 sky130_fd_sc_hd__a21o_2 _2316_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_2_.Q ),
    .A2(_1906_),
    .B1(_1908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2317_ (.A0(clknet_1_1__leaf__0702_),
    .A1(clknet_1_0__leaf__0895_),
    .A2(clknet_1_1__leaf__0626_),
    .A3(clknet_1_1__leaf__0564_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1909_));
 sky130_fd_sc_hd__nand2_2 _2318_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1910_));
 sky130_fd_sc_hd__o211a_1 _2319_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0534_),
    .B1(_0173_),
    .C1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1911_));
 sky130_fd_sc_hd__a22o_1 _2320_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_2_.Q ),
    .A2(_1909_),
    .B1(_1910_),
    .B2(_1911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2321_ (.A0(clknet_1_0__leaf__0626_),
    .A1(clknet_1_1__leaf__0564_),
    .A2(clknet_1_1__leaf__0537_),
    .A3(clknet_1_1__leaf__0665_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1912_));
 sky130_fd_sc_hd__and2b_1 _2322_ (.A_N(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _2323_ (.A0(clknet_1_0__leaf__0653_),
    .A1(clknet_1_1__leaf__0224_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1914_));
 sky130_fd_sc_hd__a22o_2 _2324_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .A2(_1912_),
    .B1(_1913_),
    .B2(_1914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2325_ (.A0(clknet_1_1__leaf__0537_),
    .A1(clknet_1_1__leaf__0665_),
    .A2(net412),
    .A3(clknet_1_1__leaf__0593_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1915_));
 sky130_fd_sc_hd__nand2b_1 _2326_ (.A_N(clknet_1_1__leaf__0677_),
    .B(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1916_));
 sky130_fd_sc_hd__o211a_2 _2327_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0257_),
    .B1(_1916_),
    .C1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1917_));
 sky130_fd_sc_hd__mux2_1 _2328_ (.A0(_1917_),
    .A1(_1915_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2329_ (.A0(net411),
    .A1(clknet_1_1__leaf__0593_),
    .A2(net349),
    .A3(clknet_1_0__leaf__0879_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1918_));
 sky130_fd_sc_hd__mux2_1 _2330_ (.A0(net303),
    .A1(clknet_1_1__leaf__0254_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1919_));
 sky130_fd_sc_hd__and3b_2 _2331_ (.A_N(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_2_.Q ),
    .B(_1919_),
    .C(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1920_));
 sky130_fd_sc_hd__a21o_2 _2332_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_2_.Q ),
    .A2(_1918_),
    .B1(_1920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2333_ (.A0(clknet_1_1__leaf__0702_),
    .A1(clknet_1_1__leaf__0895_),
    .A2(net348),
    .A3(clknet_1_1__leaf__0879_),
    .S0(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1921_));
 sky130_fd_sc_hd__nand2_2 _2334_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1922_));
 sky130_fd_sc_hd__o211a_1 _2335_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0534_),
    .B1(_0174_),
    .C1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1923_));
 sky130_fd_sc_hd__a22o_2 _2336_ (.A1(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_2_.Q ),
    .A2(_1921_),
    .B1(_1922_),
    .B2(_1923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2337_ (.A0(clknet_1_0__leaf__0730_),
    .A1(clknet_1_0__leaf__0698_),
    .A2(clknet_1_1__leaf__0561_),
    .A3(clknet_1_1__leaf__0221_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1924_));
 sky130_fd_sc_hd__and2b_1 _2338_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.ccff_tail ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _2339_ (.A0(clknet_1_0__leaf__0742_),
    .A1(net295),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1926_));
 sky130_fd_sc_hd__a22o_1 _2340_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.ccff_tail ),
    .A2(_1924_),
    .B1(_1925_),
    .B2(_1926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2341_ (.A0(clknet_1_1__leaf__0607_),
    .A1(clknet_1_1__leaf__0738_),
    .A2(clknet_1_1__leaf__0820_),
    .A3(clknet_1_0__leaf__0764_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1927_));
 sky130_fd_sc_hd__and2b_1 _2342_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1928_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(clknet_1_0__leaf__0742_),
    .A1(net294),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1929_));
 sky130_fd_sc_hd__a22o_1 _2344_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_2_.Q ),
    .A2(_1927_),
    .B1(_1928_),
    .B2(_1929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2345_ (.A0(clknet_1_1__leaf__0709_),
    .A1(clknet_1_1__leaf__0661_),
    .A2(clknet_1_1__leaf__0590_),
    .A3(clknet_1_1__leaf__0251_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1930_));
 sky130_fd_sc_hd__and2b_1 _2346_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1931_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(clknet_1_1__leaf__0607_),
    .A1(clknet_1_0__leaf__0820_),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1932_));
 sky130_fd_sc_hd__a22o_1 _2348_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_2_.Q ),
    .A2(_1930_),
    .B1(_1931_),
    .B2(_1932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2349_ (.A0(clknet_1_1__leaf__0544_),
    .A1(clknet_1_0__leaf__0586_),
    .A2(clknet_1_1__leaf__0525_),
    .A3(clknet_1_1__leaf__0578_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1933_));
 sky130_fd_sc_hd__and2b_1 _2350_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1934_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(clknet_1_0__leaf__0709_),
    .A1(clknet_1_1__leaf__0590_),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1935_));
 sky130_fd_sc_hd__a22o_2 _2352_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_2_.Q ),
    .A2(_1933_),
    .B1(_1934_),
    .B2(_1935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2353_ (.A0(clknet_1_0__leaf__0730_),
    .A1(clknet_1_0__leaf__0698_),
    .A2(clknet_1_1__leaf__0561_),
    .A3(clknet_1_1__leaf__0221_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(clknet_1_1__leaf__0544_),
    .A1(clknet_1_0__leaf__0586_),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1937_));
 sky130_fd_sc_hd__and3b_2 _2355_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_2_.Q ),
    .B(_1937_),
    .C(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1938_));
 sky130_fd_sc_hd__a21o_2 _2356_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_2_.Q ),
    .A2(_1936_),
    .B1(_1938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2357_ (.A0(clknet_1_0__leaf__0730_),
    .A1(clknet_1_1__leaf__0738_),
    .A2(clknet_1_1__leaf__0561_),
    .A3(clknet_1_1__leaf__0764_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1939_));
 sky130_fd_sc_hd__and2b_1 _2358_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1940_));
 sky130_fd_sc_hd__mux2_1 _2359_ (.A0(clknet_1_0__leaf__0742_),
    .A1(net293),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1941_));
 sky130_fd_sc_hd__a22o_2 _2360_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_2_.Q ),
    .A2(_1939_),
    .B1(_1940_),
    .B2(_1941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2361_ (.A0(clknet_1_1__leaf__0738_),
    .A1(clknet_1_0__leaf__0764_),
    .A2(clknet_1_1__leaf__0661_),
    .A3(clknet_1_1__leaf__0251_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1942_));
 sky130_fd_sc_hd__and2b_1 _2362_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1943_));
 sky130_fd_sc_hd__mux2_1 _2363_ (.A0(clknet_1_1__leaf__0607_),
    .A1(clknet_1_1__leaf__0820_),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1944_));
 sky130_fd_sc_hd__a22o_2 _2364_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_2_.Q ),
    .A2(_1942_),
    .B1(_1943_),
    .B2(_1944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2365_ (.A0(clknet_1_1__leaf__0661_),
    .A1(clknet_1_1__leaf__0525_),
    .A2(clknet_1_1__leaf__0251_),
    .A3(clknet_1_1__leaf__0578_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1945_));
 sky130_fd_sc_hd__and2b_1 _2366_ (.A_N(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1946_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(clknet_1_1__leaf__0709_),
    .A1(clknet_1_1__leaf__0590_),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1947_));
 sky130_fd_sc_hd__a22o_2 _2368_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_2_.Q ),
    .A2(_1945_),
    .B1(_1946_),
    .B2(_1947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux2_1 _2369_ (.A0(clknet_1_0__leaf__0525_),
    .A1(clknet_1_0__leaf__1314_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1948_));
 sky130_fd_sc_hd__mux2_1 _2370_ (.A0(clknet_1_0__leaf__0544_),
    .A1(clknet_1_0__leaf__0646_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1949_));
 sky130_fd_sc_hd__mux2_1 _2371_ (.A0(_1949_),
    .A1(_1948_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1950_));
 sky130_fd_sc_hd__nand2_2 _2372_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1951_));
 sky130_fd_sc_hd__o2111a_2 _2373_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0813_),
    .B1(_1951_),
    .C1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_1_.Q ),
    .D1(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1952_));
 sky130_fd_sc_hd__a21o_2 _2374_ (.A1(\dut_0.U0_formal_verification.cby_0__1__1_ccff_tail ),
    .A2(_1950_),
    .B1(_1952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2375_ (.A0(clknet_1_0__leaf__0831_),
    .A1(clknet_1_1__leaf__1395_),
    .A2(clknet_1_0__leaf__0590_),
    .A3(clknet_1_0__leaf__0251_),
    .S0(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1953_));
 sky130_fd_sc_hd__nand2_2 _2376_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1954_));
 sky130_fd_sc_hd__o2111a_2 _2377_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0813_),
    .B1(_1954_),
    .C1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_1_.Q ),
    .D1(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1955_));
 sky130_fd_sc_hd__a21o_2 _2378_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_2_.Q ),
    .A2(_1953_),
    .B1(_1955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_ ));
 sky130_fd_sc_hd__and2b_1 _2379_ (.A_N(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1956_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(clknet_1_1__leaf__0831_),
    .A1(clknet_1_1__leaf__0590_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1957_));
 sky130_fd_sc_hd__mux4_2 _2381_ (.A0(clknet_1_0__leaf__0607_),
    .A1(clknet_1_0__leaf__0738_),
    .A2(clknet_1_1__leaf__0586_),
    .A3(clknet_1_0__leaf__0578_),
    .S0(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1958_));
 sky130_fd_sc_hd__a22o_2 _2382_ (.A1(_1956_),
    .A2(_1957_),
    .B1(_1958_),
    .B2(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2b_2 _2383_ (.A_N(clknet_1_0__leaf__0586_),
    .B(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1959_));
 sky130_fd_sc_hd__mux4_2 _2384_ (.A0(clknet_1_0__leaf__0709_),
    .A1(clknet_1_0__leaf__0661_),
    .A2(clknet_1_0__leaf__0561_),
    .A3(clknet_1_0__leaf__0221_),
    .S0(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1960_));
 sky130_fd_sc_hd__o211a_2 _2385_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0607_),
    .B1(_1959_),
    .C1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(_1961_),
    .A1(_1960_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(clknet_1_0__leaf__0525_),
    .A1(clknet_1_1__leaf__1314_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1962_));
 sky130_fd_sc_hd__mux2_1 _2388_ (.A0(clknet_1_0__leaf__0544_),
    .A1(clknet_1_0__leaf__0646_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(_1963_),
    .A1(_1962_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1964_));
 sky130_fd_sc_hd__nand2b_2 _2390_ (.A_N(clknet_1_0__leaf__0561_),
    .B(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1965_));
 sky130_fd_sc_hd__o211a_2 _2391_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0709_),
    .B1(_1965_),
    .C1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1966_));
 sky130_fd_sc_hd__mux2_1 _2392_ (.A0(_1966_),
    .A1(_1964_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2393_ (.A0(clknet_1_0__leaf__0544_),
    .A1(clknet_1_0__leaf__0646_),
    .A2(clknet_1_0__leaf__1395_),
    .A3(clknet_1_0__leaf__0251_),
    .S0(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1967_));
 sky130_fd_sc_hd__nand2_2 _2394_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1968_));
 sky130_fd_sc_hd__o2111a_2 _2395_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0813_),
    .B1(_1968_),
    .C1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_1_.Q ),
    .D1(_0177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1969_));
 sky130_fd_sc_hd__a21o_2 _2396_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_2_.Q ),
    .A2(_1967_),
    .B1(_1969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2397_ (.A0(clknet_1_0__leaf__1395_),
    .A1(clknet_1_0__leaf__0738_),
    .A2(clknet_1_0__leaf__0251_),
    .A3(clknet_1_1__leaf__0578_),
    .S0(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1970_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(clknet_1_0__leaf__0831_),
    .A1(clknet_1_0__leaf__0590_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1971_));
 sky130_fd_sc_hd__and3b_2 _2399_ (.A_N(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_2_.Q ),
    .B(_1971_),
    .C(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1972_));
 sky130_fd_sc_hd__a21o_2 _2400_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_2_.Q ),
    .A2(_1970_),
    .B1(_1972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2401_ (.A0(clknet_1_0__leaf__0738_),
    .A1(clknet_1_0__leaf__0661_),
    .A2(clknet_1_1__leaf__0578_),
    .A3(clknet_1_0__leaf__0221_),
    .S0(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1973_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(clknet_1_1__leaf__0607_),
    .A1(clknet_1_0__leaf__0586_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1974_));
 sky130_fd_sc_hd__and3b_2 _2403_ (.A_N(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_2_.Q ),
    .B(_1974_),
    .C(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1975_));
 sky130_fd_sc_hd__a21o_2 _2404_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_2_.Q ),
    .A2(_1973_),
    .B1(_1975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2_2 _2405_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1976_));
 sky130_fd_sc_hd__or2_1 _2406_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1977_));
 sky130_fd_sc_hd__a31o_1 _2407_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_2_.Q ),
    .A2(_1976_),
    .A3(_1977_),
    .B1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1978_));
 sky130_fd_sc_hd__o211a_2 _2408_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0669_),
    .B1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_2_.Q ),
    .C1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1979_));
 sky130_fd_sc_hd__a21bo_2 _2409_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0550_),
    .B1_N(_1979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1980_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(clknet_1_1__leaf__0227_),
    .A1(clknet_1_0__leaf__0615_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1981_));
 sky130_fd_sc_hd__o211a_1 _2411_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_2_.Q ),
    .A2(_1981_),
    .B1(_1980_),
    .C1(_1978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_7.out ));
 sky130_fd_sc_hd__mux4_2 _2412_ (.A0(clknet_1_1__leaf__0621_),
    .A1(clknet_1_1__leaf__0596_),
    .A2(net322),
    .A3(net399),
    .S0(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1982_));
 sky130_fd_sc_hd__nand2_2 _2413_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1983_));
 sky130_fd_sc_hd__o211a_1 _2414_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0679_),
    .B1(_0178_),
    .C1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1984_));
 sky130_fd_sc_hd__a22o_2 _2415_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_2_.Q ),
    .A2(_1982_),
    .B1(_1983_),
    .B2(_1984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_6.out ));
 sky130_fd_sc_hd__mux4_1 _2416_ (.A0(clknet_1_1__leaf__1054_),
    .A1(clknet_1_1__leaf__0849_),
    .A2(clknet_1_1__leaf__0232_),
    .A3(net374),
    .S0(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_2 _2417_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1986_));
 sky130_fd_sc_hd__o2111a_2 _2418_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0621_),
    .B1(_1986_),
    .C1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_1_.Q ),
    .D1(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1987_));
 sky130_fd_sc_hd__a21o_1 _2419_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_2_.Q ),
    .A2(_1985_),
    .B1(_1987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_5.out ));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(clknet_1_1__leaf__0568_),
    .A1(clknet_1_1__leaf__0639_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1988_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(clknet_1_1__leaf__1054_),
    .A1(clknet_1_1__leaf__0232_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1989_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(_1988_),
    .A1(_1989_),
    .S(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1990_));
 sky130_fd_sc_hd__nor2_2 _2423_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1991_));
 sky130_fd_sc_hd__a211o_1 _2424_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0553_),
    .B1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_2_.Q ),
    .C1(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1992_));
 sky130_fd_sc_hd__a2bb2o_1 _2425_ (.A1_N(_1991_),
    .A2_N(_1992_),
    .B1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_2_.Q ),
    .B2(_1990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_4.out ));
 sky130_fd_sc_hd__mux4_2 _2426_ (.A0(clknet_1_1__leaf__0568_),
    .A1(clknet_1_0__leaf__0639_),
    .A2(clknet_1_1__leaf__0668_),
    .A3(clknet_1_1__leaf__0550_),
    .S0(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1993_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(clknet_1_1__leaf__0227_),
    .A1(clknet_1_1__leaf__0615_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1994_));
 sky130_fd_sc_hd__and3b_2 _2428_ (.A_N(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_2_.Q ),
    .B(_1994_),
    .C(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1995_));
 sky130_fd_sc_hd__a21o_2 _2429_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_2_.Q ),
    .A2(_1993_),
    .B1(_1995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_3.out ));
 sky130_fd_sc_hd__mux4_2 _2430_ (.A0(clknet_1_1__leaf__0668_),
    .A1(clknet_1_1__leaf__0596_),
    .A2(clknet_1_1__leaf__0550_),
    .A3(net398),
    .S0(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1996_));
 sky130_fd_sc_hd__nand2_2 _2431_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1997_));
 sky130_fd_sc_hd__o211a_1 _2432_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0679_),
    .B1(_0181_),
    .C1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1998_));
 sky130_fd_sc_hd__a22o_2 _2433_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_2_.Q ),
    .A2(_1996_),
    .B1(_1997_),
    .B2(_1998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_2.out ));
 sky130_fd_sc_hd__mux4_2 _2434_ (.A0(clknet_1_1__leaf__0596_),
    .A1(clknet_1_1__leaf__0849_),
    .A2(net397),
    .A3(net373),
    .S0(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1999_));
 sky130_fd_sc_hd__nand2_2 _2435_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2000_));
 sky130_fd_sc_hd__o2111a_2 _2436_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0621_),
    .B1(_2000_),
    .C1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_1_.Q ),
    .D1(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2001_));
 sky130_fd_sc_hd__a21o_2 _2437_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_2_.Q ),
    .A2(_1999_),
    .B1(_2001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.out ));
 sky130_fd_sc_hd__mux4_2 _2438_ (.A0(clknet_1_0__leaf__1054_),
    .A1(clknet_1_0__leaf__0849_),
    .A2(clknet_1_1__leaf__0232_),
    .A3(net372),
    .S0(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2002_));
 sky130_fd_sc_hd__nand2_1 _2439_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2003_));
 sky130_fd_sc_hd__o2111a_2 _2440_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__1077_),
    .B1(_2003_),
    .C1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_1_.Q ),
    .D1(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2004_));
 sky130_fd_sc_hd__a21o_2 _2441_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_2_.Q ),
    .A2(_2002_),
    .B1(_2004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.out ));
 sky130_fd_sc_hd__mux4_2 _2442_ (.A0(clknet_1_0__leaf__0227_),
    .A1(clknet_1_0__leaf__0568_),
    .A2(net321),
    .A3(net396),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2005_));
 sky130_fd_sc_hd__nand2_2 _2443_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2006_));
 sky130_fd_sc_hd__o2111a_2 _2444_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0793_),
    .B1(_2006_),
    .C1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_1_.Q ),
    .D1(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2007_));
 sky130_fd_sc_hd__a21o_2 _2445_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_2_.Q ),
    .A2(_2005_),
    .B1(_2007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2446_ (.A0(clknet_1_1__leaf__0679_),
    .A1(clknet_1_0__leaf__0668_),
    .A2(clknet_1_0__leaf__0232_),
    .A3(net371),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2008_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(clknet_1_0__leaf__0228_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .S(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2009_));
 sky130_fd_sc_hd__or3b_2 _2448_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_2_.Q ),
    .B(_2009_),
    .C_N(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2010_));
 sky130_fd_sc_hd__a21bo_2 _2449_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_2_.Q ),
    .A2(_2008_),
    .B1_N(_2010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_1 _2450_ (.A0(clknet_1_0__leaf__0621_),
    .A1(clknet_1_0__leaf__1061_),
    .A2(clknet_1_0__leaf__0596_),
    .A3(clknet_1_0__leaf__1238_),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2011_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(clknet_1_0__leaf__0679_),
    .A1(clknet_1_0__leaf__0232_),
    .S(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2012_));
 sky130_fd_sc_hd__and3b_2 _2452_ (.A_N(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_2_.Q ),
    .B(_2012_),
    .C(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2013_));
 sky130_fd_sc_hd__a21o_1 _2453_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_2_.Q ),
    .A2(_2011_),
    .B1(_2013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2454_ (.A0(clknet_1_0__leaf__0621_),
    .A1(clknet_1_0__leaf__0897_),
    .A2(clknet_1_1__leaf__1061_),
    .A3(clknet_1_0__leaf__0550_),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2014_));
 sky130_fd_sc_hd__nand2_2 _2455_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2015_));
 sky130_fd_sc_hd__o2111a_2 _2456_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0881_),
    .B1(_2015_),
    .C1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_1_.Q ),
    .D1(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2016_));
 sky130_fd_sc_hd__a21o_2 _2457_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_2_.Q ),
    .A2(_2014_),
    .B1(_2016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2458_ (.A0(clknet_1_1__leaf__0897_),
    .A1(clknet_1_0__leaf__0568_),
    .A2(clknet_1_0__leaf__0550_),
    .A3(net395),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2017_));
 sky130_fd_sc_hd__nand2_2 _2459_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2018_));
 sky130_fd_sc_hd__o2111a_2 _2460_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0793_),
    .B1(_2018_),
    .C1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_1_.Q ),
    .D1(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2019_));
 sky130_fd_sc_hd__a21o_2 _2461_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_2_.Q ),
    .A2(_2017_),
    .B1(_2019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2462_ (.A0(clknet_1_0__leaf__0568_),
    .A1(clknet_1_0__leaf__0668_),
    .A2(net394),
    .A3(net370),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2020_));
 sky130_fd_sc_hd__mux2_1 _2463_ (.A0(clknet_1_1__leaf__0228_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .S(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2021_));
 sky130_fd_sc_hd__or3b_2 _2464_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_2_.Q ),
    .B(_2021_),
    .C_N(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2022_));
 sky130_fd_sc_hd__a21bo_2 _2465_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_2_.Q ),
    .A2(_2020_),
    .B1_N(_2022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2466_ (.A0(clknet_1_0__leaf__0668_),
    .A1(clknet_1_1__leaf__0596_),
    .A2(net369),
    .A3(clknet_1_1__leaf__1238_),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2023_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(clknet_1_1__leaf__0679_),
    .A1(clknet_1_0__leaf__0232_),
    .S(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2024_));
 sky130_fd_sc_hd__and3b_2 _2468_ (.A_N(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_2_.Q ),
    .B(_2024_),
    .C(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2025_));
 sky130_fd_sc_hd__a21o_2 _2469_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_2_.Q ),
    .A2(_2023_),
    .B1(_2025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_ ));
 sky130_fd_sc_hd__mux4_2 _2470_ (.A0(clknet_1_0__leaf__0621_),
    .A1(clknet_1_1__leaf__1061_),
    .A2(clknet_1_0__leaf__0596_),
    .A3(clknet_1_1__leaf__1238_),
    .S0(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2026_));
 sky130_fd_sc_hd__nand2_2 _2471_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2027_));
 sky130_fd_sc_hd__o2111a_2 _2472_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0881_),
    .B1(_2027_),
    .C1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_1_.Q ),
    .D1(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2028_));
 sky130_fd_sc_hd__a21o_2 _2473_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_2_.Q ),
    .A2(_2026_),
    .B1(_2028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_ ));
 sky130_fd_sc_hd__nand2_1 _2474_ (.A(net221),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0028_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(net219),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0026_));
 sky130_fd_sc_hd__nand2_1 _2476_ (.A(net219),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2_1 _2477_ (.A(net219),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0022_));
 sky130_fd_sc_hd__nand2_1 _2478_ (.A(net220),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0020_));
 sky130_fd_sc_hd__nand2_1 _2479_ (.A(net219),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _2480_ (.A(net219),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0016_));
 sky130_fd_sc_hd__nand2_1 _2481_ (.A(net222),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2_1 _2482_ (.A(net222),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0012_));
 sky130_fd_sc_hd__nand2_1 _2483_ (.A(net222),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _2484_ (.A(net222),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_1 _2485_ (.A(net221),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_1 _2486_ (.A(net220),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_1 _2487_ (.A(net220),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _2488_ (.A(net221),
    .B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0000_));
 sky130_fd_sc_hd__clkbuf_1 _2489_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _2490_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _2492_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2061_));
 sky130_fd_sc_hd__clkbuf_1 _2493_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_1 _2494_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2059_));
 sky130_fd_sc_hd__clkbuf_1 _2495_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _2496_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _2497_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2048_));
 sky130_fd_sc_hd__clkbuf_1 _2498_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _2499_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _2501_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2043_));
 sky130_fd_sc_hd__clkbuf_1 _2503_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2034_));
 sky130_fd_sc_hd__clkbuf_1 _2504_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2033_));
 sky130_fd_sc_hd__clkbuf_1 _2505_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _2506_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2031_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2030_));
 sky130_fd_sc_hd__clkbuf_1 _2508_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _2509_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2156_));
 sky130_fd_sc_hd__clkbuf_1 _2510_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2147_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_1 _2512_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2145_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2144_));
 sky130_fd_sc_hd__clkbuf_1 _2514_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2143_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2142_));
 sky130_fd_sc_hd__clkbuf_1 _2516_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2141_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2132_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2131_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2130_));
 sky130_fd_sc_hd__buf_1 _2520_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2129_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _2522_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2127_));
 sky130_fd_sc_hd__buf_1 _2523_ (.A(\dut_0.U0_formal_verification.grid_io_right_1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2126_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _2525_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2116_));
 sky130_fd_sc_hd__clkbuf_1 _2526_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2115_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_1 _2528_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2113_));
 sky130_fd_sc_hd__clkbuf_1 _2529_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2112_));
 sky130_fd_sc_hd__clkbuf_1 _2530_ (.A(\dut_0.U0_formal_verification.grid_io_right_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2111_));
 sky130_fd_sc_hd__clkbuf_1 _2531_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2102_));
 sky130_fd_sc_hd__clkbuf_1 _2532_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2101_));
 sky130_fd_sc_hd__clkbuf_1 _2533_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_1 _2534_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2099_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2098_));
 sky130_fd_sc_hd__clkbuf_1 _2536_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2097_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(\dut_0.U0_formal_verification.grid_io_top_1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2096_));
 sky130_fd_sc_hd__clkbuf_1 _2538_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2088_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2087_));
 sky130_fd_sc_hd__clkbuf_1 _2540_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _2541_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2085_));
 sky130_fd_sc_hd__clkbuf_1 _2542_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2084_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_1 _2544_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_1 _2545_ (.A(\dut_0.U0_formal_verification.grid_io_top_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2081_));
 sky130_fd_sc_hd__clkbuf_1 _2546_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _2548_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2148_));
 sky130_fd_sc_hd__clkbuf_1 _2550_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2118_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2103_));
 sky130_fd_sc_hd__inv_2 _2644__17 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _2555__7 (.A(clknet_1_1__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _2566__8 (.A(clknet_1_0__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _2557__2 (.A(clknet_1_0__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _2558__3 (.A(clknet_1_0__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _2559__4 (.A(clknet_1_0__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _2561__5 (.A(clknet_1_1__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _2563__11 (.A(clknet_1_0__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _2554__6 (.A(clknet_1_1__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _2553__16 (.A(clknet_1_1__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _2564__12 (.A(clknet_1_0__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _2565__13 (.A(clknet_1_0__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _2567__14 (.A(clknet_1_0__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _2789__9 (.A(clknet_1_1__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _2562__15 (.A(clknet_1_1__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _2568_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2072_));
 sky130_fd_sc_hd__inv_2 _2569_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2071_));
 sky130_fd_sc_hd__inv_2 _2570_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2070_));
 sky130_fd_sc_hd__inv_2 _2571_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2069_));
 sky130_fd_sc_hd__inv_2 _2572_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2068_));
 sky130_fd_sc_hd__inv_2 _2573_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2067_));
 sky130_fd_sc_hd__inv_2 _2574_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2066_));
 sky130_fd_sc_hd__inv_2 _2575_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2057_));
 sky130_fd_sc_hd__inv_2 _2576_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2056_));
 sky130_fd_sc_hd__inv_2 _2577_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2055_));
 sky130_fd_sc_hd__inv_2 _2578_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2054_));
 sky130_fd_sc_hd__inv_2 _2579_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2053_));
 sky130_fd_sc_hd__inv_2 _2580_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2052_));
 sky130_fd_sc_hd__inv_2 _2581_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2051_));
 sky130_fd_sc_hd__inv_2 _2582_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2042_));
 sky130_fd_sc_hd__inv_2 _2583_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2041_));
 sky130_fd_sc_hd__inv_2 _2584_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2040_));
 sky130_fd_sc_hd__inv_2 _2585_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2039_));
 sky130_fd_sc_hd__inv_2 _2586_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2038_));
 sky130_fd_sc_hd__inv_2 _2587_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2037_));
 sky130_fd_sc_hd__inv_2 _2588_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2036_));
 sky130_fd_sc_hd__inv_2 _2589_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2155_));
 sky130_fd_sc_hd__inv_2 _2590_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2154_));
 sky130_fd_sc_hd__inv_2 _2591_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2153_));
 sky130_fd_sc_hd__inv_2 _2592_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2152_));
 sky130_fd_sc_hd__inv_2 _2593_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2151_));
 sky130_fd_sc_hd__inv_2 _2594_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2150_));
 sky130_fd_sc_hd__inv_2 _2595_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2149_));
 sky130_fd_sc_hd__inv_2 _2596_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2140_));
 sky130_fd_sc_hd__inv_2 _2597_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2139_));
 sky130_fd_sc_hd__inv_2 _2598_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2138_));
 sky130_fd_sc_hd__inv_2 _2599_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2137_));
 sky130_fd_sc_hd__inv_2 _2600_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2136_));
 sky130_fd_sc_hd__inv_2 _2601_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2135_));
 sky130_fd_sc_hd__inv_2 _2602_ (.A(\dut_0.U0_formal_verification.grid_io_right_1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2134_));
 sky130_fd_sc_hd__inv_2 _2603_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2125_));
 sky130_fd_sc_hd__inv_2 _2604_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2124_));
 sky130_fd_sc_hd__inv_2 _2605_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2123_));
 sky130_fd_sc_hd__inv_2 _2606_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2122_));
 sky130_fd_sc_hd__inv_2 _2607_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2121_));
 sky130_fd_sc_hd__inv_2 _2608_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2120_));
 sky130_fd_sc_hd__inv_2 _2609_ (.A(\dut_0.U0_formal_verification.grid_io_right_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2119_));
 sky130_fd_sc_hd__inv_2 _2610_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2110_));
 sky130_fd_sc_hd__inv_2 _2611_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2109_));
 sky130_fd_sc_hd__inv_2 _2612_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2108_));
 sky130_fd_sc_hd__inv_2 _2613_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2107_));
 sky130_fd_sc_hd__inv_2 _2614_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2106_));
 sky130_fd_sc_hd__inv_2 _2615_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2105_));
 sky130_fd_sc_hd__inv_2 _2616_ (.A(\dut_0.U0_formal_verification.grid_io_top_1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2104_));
 sky130_fd_sc_hd__inv_2 _2617_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2095_));
 sky130_fd_sc_hd__inv_2 _2618_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2094_));
 sky130_fd_sc_hd__inv_2 _2619_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2093_));
 sky130_fd_sc_hd__inv_2 _2620_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2092_));
 sky130_fd_sc_hd__inv_2 _2621_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2091_));
 sky130_fd_sc_hd__inv_2 _2622_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2090_));
 sky130_fd_sc_hd__inv_2 _2623_ (.A(\dut_0.U0_formal_verification.grid_io_top_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2089_));
 sky130_fd_sc_hd__inv_2 _2624_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2080_));
 sky130_fd_sc_hd__inv_2 _2625_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2079_));
 sky130_fd_sc_hd__inv_2 _2626_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2078_));
 sky130_fd_sc_hd__inv_2 _2627_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2077_));
 sky130_fd_sc_hd__inv_2 _2628_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2076_));
 sky130_fd_sc_hd__inv_2 _2629_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2075_));
 sky130_fd_sc_hd__inv_2 _2630_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2074_));
 sky130_fd_sc_hd__inv_2 _2631_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _2632_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _2633_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _2634_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _2635_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _2636_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _2637_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _2638_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _2639_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _2640_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _2641_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _2642_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _2643_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _3191__18 (.A(clknet_1_0__leaf__0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _2645_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _2646_ (.A(\dut_0.U0_formal_verification.cby_1__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _2647_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _2648_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _2649_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _2650_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _2651_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _2652_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _2653_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _2654_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _2655_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _2656_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _2657_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _2658_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _2659_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _2660_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _2661_ (.A(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _2662_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _2663_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _2664_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _2665_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _2666_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _2667_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _2668_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _2669_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _2670_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _2671_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _2672_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _2673_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _2674_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _2675_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _2676_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _2677_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _2678_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _2679_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _2680_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _2681_ (.A(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _2682_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _2683_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _2684_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _2685_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _2686_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _2687_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _2688_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _2689_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _2690_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _2691_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _2692_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _2693_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _2694_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _2695_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _2696_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _2697_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _2698_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _2699_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _2700_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _2701_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _2702_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _2703_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _2704_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _2705_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _2706_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _2707_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _2708_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _2709_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _2710_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _2711_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _2712_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _2713_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _2714_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _2715_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _2716_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _2717_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _2718_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _2719_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _2720_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _2721_ (.A(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _2722_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _2723_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _2724_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _2725_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _2726_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _2727_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _2728_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _2729_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _2730_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _2731_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _2732_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _2733_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _2734_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _2735_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _2736_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _2737_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _2738_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _2739_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _2740_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _2741_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _2742_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _2743_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _2744_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _2745_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _2746_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _2747_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _2748_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _2749_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _2750_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _2751_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _2752_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _2753_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _2754_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _2755_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _2756_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _2757_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _2758_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _2759_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _2760_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _2761_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _2762_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _2763_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _2764_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _2765_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _2766_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _2767_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _2768_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _2769_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _2770_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _2771_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _2772_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _2773_ (.A(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _2774_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _2775_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _2776_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _2777_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _2778_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _2779_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _2780_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _2781_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _2782_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _2783_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _2784_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _2785_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _2786_ (.A(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _2787_ (.A(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.RST ));
 sky130_fd_sc_hd__inv_2 _2788_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2073_));
 sky130_fd_sc_hd__inv_2 _2560__10 (.A(clknet_1_0__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _3011__47 (.A(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _2791_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _2792_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _3257__41 (.A(clknet_1_1__leaf__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _2794_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _2795_ (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _2793__39 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _3286__97 (.A(clknet_1_0__leaf__0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _2802__21 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _2799_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _2800_ (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _2796__37 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _2819__26 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _2810__131 (.A(clknet_1_0__leaf_net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _2804_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _3487__143 (.A(_0862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _2797__95 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _3465__187 (.A(_0842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _3978__74 (.A(_1326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _3874__157 (.A(_1229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _2820__133 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _3741__103 (.A(clknet_1_0__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _3985__119 (.A(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _3270__182 (.A(clknet_1_1__leaf__0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _3436__165 (.A(_0817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _2806__88 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _2817__55 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _3360__57 (.A(clknet_1_0__leaf__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _2812__111 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _2801__31 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _3335__140 (.A(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net375));
 sky130_fd_sc_hd__nand2_1 _2821_ (.A(net219),
    .B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2b_2 _2822_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0219_));
 sky130_fd_sc_hd__nand2b_2 _2823_ (.A_N(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0220_));
 sky130_fd_sc_hd__and3_2 _2824_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0219_),
    .C(clknet_1_0__leaf__0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__a31o_2 _2825_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0219_),
    .A3(clknet_1_1__leaf__0220_),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__o21a_4 _2826_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .A2(_0038_),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__and2_2 _2827_ (.A(clknet_1_0__leaf__0222_),
    .B(clknet_1_0__leaf__0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_2 _2828_ (.A1(clknet_1_1__leaf__0222_),
    .A2(clknet_1_1__leaf__0223_),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__nand2b_2 _2829_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0226_));
 sky130_fd_sc_hd__and3_2 _2830_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0225_),
    .C(clknet_1_1__leaf__0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__nand3_2 _2831_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0225_),
    .C(clknet_1_0__leaf__0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_2 _2832_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_9.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2b_2 _2833_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2b_2 _2834_ (.A_N(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_8.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0231_));
 sky130_fd_sc_hd__and3_2 _2835_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.D ),
    .B(clknet_1_0__leaf__0230_),
    .C(clknet_1_1__leaf__0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__o211a_2 _2836_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_9.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0232_),
    .B1(_0229_),
    .C1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__inv_2 _2813__174 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net409));
 sky130_fd_sc_hd__o21ai_2 _2838_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0233_),
    .B1(\dut_0.U0_formal_verification.cbx_1__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0235_));
 sky130_fd_sc_hd__a21o_2 _2839_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .B1(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__o21ai_2 _2840_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .A2(net390),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0237_));
 sky130_fd_sc_hd__a21o_2 _2841_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(net41),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__o211a_2 _2843_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .A2(_0239_),
    .B1(_0238_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__nand2_1 _2844_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0241_));
 sky130_fd_sc_hd__or2_1 _2845_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__a31o_1 _2846_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .A2(_0241_),
    .A3(_0242_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__nor2_2 _2847_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .B(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0244_));
 sky130_fd_sc_hd__a31o_2 _2848_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0225_),
    .A3(clknet_1_0__leaf__0226_),
    .B1(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__or2_2 _2849_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__and3_2 _2850_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0245_),
    .C(clknet_1_1__leaf__0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__nand3_2 _2851_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0245_),
    .C(clknet_1_0__leaf__0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0248_));
 sky130_fd_sc_hd__a31o_2 _2852_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0245_),
    .A3(clknet_1_0__leaf__0246_),
    .B1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__nand2b_2 _2853_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0250_));
 sky130_fd_sc_hd__and3_2 _2854_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0249_),
    .C(clknet_1_1__leaf__0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__a31o_2 _2855_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0249_),
    .A3(clknet_1_0__leaf__0250_),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__nand2b_1 _2856_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0253_));
 sky130_fd_sc_hd__and3_4 _2857_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.D ),
    .B(clknet_1_0__leaf__0252_),
    .C(clknet_1_0__leaf__0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__a31o_2 _2858_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.D ),
    .A2(clknet_1_1__leaf__0230_),
    .A3(clknet_1_0__leaf__0231_),
    .B1(_0041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__or2_2 _2859_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__and3_2 _2860_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0255_),
    .C(clknet_1_0__leaf__0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(clknet_1_1__leaf__0254_),
    .A1(clknet_1_1__leaf__0257_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__nand2_2 _2862_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_1_.Q ),
    .B(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0259_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(clknet_1_1__leaf__0259_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .S(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__or2_2 _2864_ (.A(_0049_),
    .B(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__mux4_2 _2865_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__nand2b_2 _2866_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .B(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0263_));
 sky130_fd_sc_hd__mux4_1 _2867_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_1 _2868_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .B(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0265_));
 sky130_fd_sc_hd__a32o_2 _2869_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .A2(_0263_),
    .A3(_0265_),
    .B1(_0243_),
    .B2(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0236_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_2 _2871_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .B(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0268_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(net41),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__inv_2 _2942__50 (.A(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net285));
 sky130_fd_sc_hd__o211a_2 _2874_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .A2(net284),
    .B1(_0268_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__nand2_1 _2875_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0272_));
 sky130_fd_sc_hd__o2111a_1 _2876_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .A2(net45),
    .B1(_0272_),
    .C1(_0036_),
    .D1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__mux4_2 _2877_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_2 _2878_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .B(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0275_));
 sky130_fd_sc_hd__mux4_2 _2879_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__o21ai_2 _2880_ (.A1(_0036_),
    .A2(_0276_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0277_));
 sky130_fd_sc_hd__o32a_2 _2881_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .A2(_0271_),
    .A3(_0273_),
    .B1(_0275_),
    .B2(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__o21ai_2 _2883_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .A2(net391),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0280_));
 sky130_fd_sc_hd__a21o_2 _2884_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(net41),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__o211a_2 _2886_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .A2(_0282_),
    .B1(_0281_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _2887_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0284_));
 sky130_fd_sc_hd__or2_1 _2888_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__a31o_1 _2889_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .A2(_0284_),
    .A3(_0285_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_2 _2890_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .B(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0287_));
 sky130_fd_sc_hd__mux4_2 _2891_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__nand2b_2 _2892_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0289_));
 sky130_fd_sc_hd__mux4_2 _2893_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_2 _2894_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .B(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0291_));
 sky130_fd_sc_hd__a32o_2 _2895_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .A2(_0289_),
    .A3(_0291_),
    .B1(_0286_),
    .B2(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(_0279_),
    .A1(_0293_),
    .S(clknet_1_0__leaf__0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__nand2b_1 _2898_ (.A_N(_0294_),
    .B(clknet_1_0__leaf__0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0295_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(_0296_),
    .A1(_0297_),
    .S(clknet_1_0__leaf__0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_2 _2902_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .A2(net384),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0299_));
 sky130_fd_sc_hd__a21o_2 _2903_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0236_),
    .B1(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(net41),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_2 _2905_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .A2(_0301_),
    .B1(_0300_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _2906_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0303_));
 sky130_fd_sc_hd__or2_1 _2907_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__a31o_1 _2908_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .A2(_0303_),
    .A3(_0304_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__nor2_2 _2909_ (.A(\dut_0.U0_formal_verification.grid_clb_0_ccff_tail ),
    .B(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0306_));
 sky130_fd_sc_hd__mux4_2 _2910_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__nand2b_2 _2911_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .B(_0307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0308_));
 sky130_fd_sc_hd__mux4_2 _2912_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_2 _2913_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .B(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0310_));
 sky130_fd_sc_hd__a32o_2 _2914_ (.A1(\dut_0.U0_formal_verification.grid_clb_0_ccff_tail ),
    .A2(_0308_),
    .A3(_0310_),
    .B1(_0305_),
    .B2(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__o21ba_2 _2915_ (.A1(clknet_1_0__leaf__0292_),
    .A2(_0298_),
    .B1_N(clknet_1_1__leaf__0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2917_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(_0313_),
    .A1(_0314_),
    .S(clknet_1_1__leaf__0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(_0317_),
    .A1(_0316_),
    .S(clknet_1_1__leaf__0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_0318_),
    .A1(_0315_),
    .S(clknet_1_1__leaf__0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_1 _2923_ (.A1(_0295_),
    .A2(_0312_),
    .B1(_0319_),
    .B2(clknet_1_0__leaf__0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _2924_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_2 _2925_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .B(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _2926_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .A2(net389),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0321_));
 sky130_fd_sc_hd__a21o_2 _2927_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(net41),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__o211a_2 _2929_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .A2(_0323_),
    .B1(_0322_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _2930_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0325_));
 sky130_fd_sc_hd__or2_1 _2931_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__a31o_1 _2932_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .A2(_0325_),
    .A3(_0326_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_2 _2933_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .B(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0328_));
 sky130_fd_sc_hd__mux4_2 _2934_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__nand2b_2 _2935_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .B(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0330_));
 sky130_fd_sc_hd__mux4_2 _2936_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_2 _2937_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .B(_0331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0332_));
 sky130_fd_sc_hd__a32o_1 _2938_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .A2(_0330_),
    .A3(_0332_),
    .B1(_0327_),
    .B2(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0236_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_2 _2940_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .B(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0335_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(net41),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__inv_2 _2816__51 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net286));
 sky130_fd_sc_hd__o211a_2 _2943_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .A2(net285),
    .B1(_0335_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__nand2_1 _2944_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0339_));
 sky130_fd_sc_hd__o2111a_1 _2945_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .A2(net46),
    .B1(_0339_),
    .C1(_0035_),
    .D1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__mux4_2 _2946_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_2 _2947_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .B(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0342_));
 sky130_fd_sc_hd__mux4_2 _2948_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net48),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__o21ai_2 _2949_ (.A1(_0035_),
    .A2(_0343_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0344_));
 sky130_fd_sc_hd__o32a_2 _2950_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .A2(_0338_),
    .A3(_0340_),
    .B1(_0342_),
    .B2(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__o21ai_2 _2952_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(net388),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0347_));
 sky130_fd_sc_hd__a21o_2 _2953_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(net41),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__o211a_2 _2955_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .A2(_0349_),
    .B1(_0348_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _2956_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0351_));
 sky130_fd_sc_hd__or2_1 _2957_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__a31o_1 _2958_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .A2(_0351_),
    .A3(_0352_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__nor2_2 _2959_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .B(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0354_));
 sky130_fd_sc_hd__mux4_2 _2960_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__nand2b_2 _2961_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .B(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0356_));
 sky130_fd_sc_hd__mux4_2 _2962_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net48),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_2 _2963_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .B(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0358_));
 sky130_fd_sc_hd__a32o_2 _2964_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .A2(_0356_),
    .A3(_0358_),
    .B1(_0353_),
    .B2(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_0346_),
    .A1(_0360_),
    .S(clknet_1_0__leaf__0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__nand2b_1 _2967_ (.A_N(_0361_),
    .B(clknet_1_0__leaf__0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0362_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_0__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_0__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(_0363_),
    .A1(_0364_),
    .S(clknet_1_0__leaf__0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__o21ai_2 _2971_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .A2(net387),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0366_));
 sky130_fd_sc_hd__a21o_2 _2972_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(net42),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__o211a_2 _2974_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .A2(_0368_),
    .B1(_0367_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__nand2_1 _2975_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0370_));
 sky130_fd_sc_hd__or2_1 _2976_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__a31o_1 _2977_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .A2(_0370_),
    .A3(_0371_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__nor2_2 _2978_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .B(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0373_));
 sky130_fd_sc_hd__mux4_2 _2979_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__nand2b_2 _2980_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .B(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0375_));
 sky130_fd_sc_hd__mux4_2 _2981_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net48),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__nand2_2 _2982_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .B(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0377_));
 sky130_fd_sc_hd__a32o_2 _2983_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .A2(_0375_),
    .A3(_0377_),
    .B1(_0372_),
    .B2(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__o21ba_2 _2984_ (.A1(clknet_1_0__leaf__0359_),
    .A2(_0365_),
    .B1_N(clknet_1_0__leaf__0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(_0380_),
    .A1(_0381_),
    .S(clknet_1_1__leaf__0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_1__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_1__leaf__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(_0384_),
    .A1(_0383_),
    .S(clknet_1_1__leaf__0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(_0385_),
    .A1(_0382_),
    .S(clknet_1_1__leaf__0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__a22o_1 _2992_ (.A1(_0362_),
    .A2(_0379_),
    .B1(_0386_),
    .B2(clknet_1_1__leaf__0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_2 _2994_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .B(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _2995_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .A2(net380),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0388_));
 sky130_fd_sc_hd__a21o_2 _2996_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0236_),
    .B1(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(net41),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__o211a_2 _2998_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .A2(_0390_),
    .B1(_0389_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_1 _2999_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0392_));
 sky130_fd_sc_hd__or2_1 _3000_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__a31o_1 _3001_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .A2(_0392_),
    .A3(_0393_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__nor2_2 _3002_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .B(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0395_));
 sky130_fd_sc_hd__mux4_2 _3003_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__nand2b_2 _3004_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .B(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0397_));
 sky130_fd_sc_hd__mux4_2 _3005_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net48),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_2 _3006_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .B(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0399_));
 sky130_fd_sc_hd__a32o_2 _3007_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .A2(_0397_),
    .A3(_0399_),
    .B1(_0394_),
    .B2(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0236_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_2 _3009_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .B(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0402_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(net42),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__inv_2 _3080__48 (.A(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net283));
 sky130_fd_sc_hd__o211a_2 _3012_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .A2(net282),
    .B1(_0402_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_1 _3013_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0406_));
 sky130_fd_sc_hd__o2111a_1 _3014_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .A2(net45),
    .B1(_0406_),
    .C1(_0034_),
    .D1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_2 _3015_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_2 _3016_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .B(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0409_));
 sky130_fd_sc_hd__mux4_2 _3017_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__o21ai_2 _3018_ (.A1(_0034_),
    .A2(_0410_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0411_));
 sky130_fd_sc_hd__o32a_2 _3019_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .A2(_0405_),
    .A3(_0407_),
    .B1(_0409_),
    .B2(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__o21ai_2 _3021_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .A2(net385),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0414_));
 sky130_fd_sc_hd__a21o_2 _3022_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(net41),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__o211a_2 _3024_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .A2(_0416_),
    .B1(_0415_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _3025_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _3026_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__a31o_1 _3027_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .A2(_0418_),
    .A3(_0419_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_2 _3028_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0421_));
 sky130_fd_sc_hd__mux4_2 _3029_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__nand2b_2 _3030_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .B(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0423_));
 sky130_fd_sc_hd__mux4_2 _3031_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net48),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_2 _3032_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .B(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0425_));
 sky130_fd_sc_hd__a32o_1 _3033_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .A2(_0423_),
    .A3(_0425_),
    .B1(_0420_),
    .B2(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3035_ (.A0(_0413_),
    .A1(_0427_),
    .S(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__nand2b_1 _3036_ (.A_N(_0428_),
    .B(clknet_1_0__leaf__0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0429_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_1__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(_0430_),
    .A1(_0431_),
    .S(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__o21ai_2 _3040_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .A2(net386),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0433_));
 sky130_fd_sc_hd__a21o_2 _3041_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0236_),
    .B1(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(net41),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__o211a_2 _3043_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .A2(_0435_),
    .B1(_0434_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0437_));
 sky130_fd_sc_hd__or2_1 _3045_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__a31o_1 _3046_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .A2(_0437_),
    .A3(_0438_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__nor2_2 _3047_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .B(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0440_));
 sky130_fd_sc_hd__mux4_2 _3048_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0261_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0441_));
 sky130_fd_sc_hd__nand2b_2 _3049_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0442_));
 sky130_fd_sc_hd__mux4_2 _3050_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net48),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_2 _3051_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .B(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0444_));
 sky130_fd_sc_hd__a32o_2 _3052_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .A2(_0442_),
    .A3(_0444_),
    .B1(_0439_),
    .B2(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__o21ba_2 _3053_ (.A1(clknet_1_1__leaf__0426_),
    .A2(_0432_),
    .B1_N(clknet_1_0__leaf__0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(_0447_),
    .A1(_0448_),
    .S(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_0__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(_0451_),
    .A1(_0450_),
    .S(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(_0452_),
    .A1(_0449_),
    .S(clknet_1_0__leaf__0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _3061_ (.A1(_0429_),
    .A2(_0446_),
    .B1(_0453_),
    .B2(clknet_1_1__leaf__0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_4 _3063_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .B(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _3064_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(net383),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0455_));
 sky130_fd_sc_hd__a21o_2 _3065_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0236_),
    .B1(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(net42),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0457_));
 sky130_fd_sc_hd__o211a_2 _3067_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .A2(_0457_),
    .B1(_0456_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0458_));
 sky130_fd_sc_hd__nand2_1 _3068_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0459_));
 sky130_fd_sc_hd__or2_1 _3069_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0460_));
 sky130_fd_sc_hd__a31o_1 _3070_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .A2(_0459_),
    .A3(_0460_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0461_));
 sky130_fd_sc_hd__nor2_2 _3071_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .B(_0458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0462_));
 sky130_fd_sc_hd__mux4_2 _3072_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0463_));
 sky130_fd_sc_hd__nand2b_2 _3073_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .B(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0464_));
 sky130_fd_sc_hd__mux4_2 _3074_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0465_));
 sky130_fd_sc_hd__nand2_2 _3075_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .B(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0466_));
 sky130_fd_sc_hd__a32o_2 _3076_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .A2(_0464_),
    .A3(_0466_),
    .B1(_0461_),
    .B2(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0236_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_2 _3078_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .B(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0469_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(net42),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0470_));
 sky130_fd_sc_hd__inv_2 _2873__49 (.A(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net284));
 sky130_fd_sc_hd__o211a_2 _3081_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .A2(net283),
    .B1(_0469_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_1 _3082_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0473_));
 sky130_fd_sc_hd__o2111a_1 _3083_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .A2(net45),
    .B1(_0473_),
    .C1(_0032_),
    .D1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0474_));
 sky130_fd_sc_hd__mux4_2 _3084_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_2 _3085_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .B(_0475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0476_));
 sky130_fd_sc_hd__mux4_2 _3086_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0477_));
 sky130_fd_sc_hd__o21ai_2 _3087_ (.A1(_0032_),
    .A2(_0477_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0478_));
 sky130_fd_sc_hd__o32a_2 _3088_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .A2(_0472_),
    .A3(_0474_),
    .B1(_0476_),
    .B2(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0480_));
 sky130_fd_sc_hd__o21ai_2 _3090_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(net382),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0481_));
 sky130_fd_sc_hd__a21o_2 _3091_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0236_),
    .B1(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(net42),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0483_));
 sky130_fd_sc_hd__o211a_2 _3093_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .A2(_0483_),
    .B1(_0482_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0484_));
 sky130_fd_sc_hd__nand2_1 _3094_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0485_));
 sky130_fd_sc_hd__o211a_1 _3095_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(net45),
    .B1(_0485_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0486_));
 sky130_fd_sc_hd__or2_1 _3096_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .B(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0487_));
 sky130_fd_sc_hd__nor2_2 _3097_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .B(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0488_));
 sky130_fd_sc_hd__mux4_2 _3098_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0489_));
 sky130_fd_sc_hd__nand2b_2 _3099_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .B(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0490_));
 sky130_fd_sc_hd__mux4_2 _3100_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_2 _3101_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .B(_0491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0492_));
 sky130_fd_sc_hd__a32o_2 _3102_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .A2(_0490_),
    .A3(_0492_),
    .B1(_0487_),
    .B2(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(_0480_),
    .A1(_0494_),
    .S(clknet_1_1__leaf__0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0495_));
 sky130_fd_sc_hd__nand2b_2 _3105_ (.A_N(_0495_),
    .B(clknet_1_0__leaf__0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0496_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_1__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(_0497_),
    .A1(_0498_),
    .S(clknet_1_1__leaf__0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_2 _3109_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0500_));
 sky130_fd_sc_hd__o211a_2 _3110_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .A2(net381),
    .B1(_0500_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(net42),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0502_));
 sky130_fd_sc_hd__o21ai_2 _3112_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .A2(_0502_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _3113_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0504_));
 sky130_fd_sc_hd__o211a_1 _3114_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .A2(net45),
    .B1(_0504_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0505_));
 sky130_fd_sc_hd__o221a_2 _3115_ (.A1(_0501_),
    .A2(_0503_),
    .B1(_0505_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .C1(_0033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0506_));
 sky130_fd_sc_hd__mux4_2 _3116_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0261_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0507_));
 sky130_fd_sc_hd__nand2b_2 _3117_ (.A_N(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .B(_0507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0508_));
 sky130_fd_sc_hd__mux4_2 _3118_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(net47),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_2 _3119_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .B(_0509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0510_));
 sky130_fd_sc_hd__a31o_2 _3120_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .A2(_0508_),
    .A3(_0510_),
    .B1(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0511_));
 sky130_fd_sc_hd__o21ba_2 _3121_ (.A1(clknet_1_1__leaf__0493_),
    .A2(_0499_),
    .B1_N(clknet_1_1__leaf__0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _3124_ (.A0(_0513_),
    .A1(_0514_),
    .S(clknet_1_0__leaf__0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_0__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(_0517_),
    .A1(_0516_),
    .S(clknet_1_0__leaf__0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(_0518_),
    .A1(_0515_),
    .S(clknet_1_0__leaf__0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_2 _3129_ (.A1(_0496_),
    .A2(_0512_),
    .B1(_0519_),
    .B2(clknet_1_0__leaf__0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_2 _3131_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .B(_0520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0521_));
 sky130_fd_sc_hd__or2_2 _3133_ (.A(_0037_),
    .B(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0522_));
 sky130_fd_sc_hd__a31o_2 _3134_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0255_),
    .A3(clknet_1_1__leaf__0256_),
    .B1(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_2 _3135_ (.A(_0042_),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0524_));
 sky130_fd_sc_hd__and3_2 _3136_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0523_),
    .C(clknet_1_0__leaf__0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0525_));
 sky130_fd_sc_hd__a31o_2 _3137_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0523_),
    .A3(clknet_1_1__leaf__0524_),
    .B1(_0043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0526_));
 sky130_fd_sc_hd__or2_1 _3138_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0527_));
 sky130_fd_sc_hd__and3_2 _3139_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0526_),
    .C(clknet_1_1__leaf__0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0528_));
 sky130_fd_sc_hd__a31o_2 _3140_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0526_),
    .A3(clknet_1_0__leaf__0527_),
    .B1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0529_));
 sky130_fd_sc_hd__nand2b_1 _3141_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0530_));
 sky130_fd_sc_hd__and3_1 _3142_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0529_),
    .C(clknet_1_0__leaf__0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0531_));
 sky130_fd_sc_hd__nand3_2 _3143_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0529_),
    .C(clknet_1_1__leaf__0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _3144_ (.A(_0044_),
    .B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0533_));
 sky130_fd_sc_hd__o211a_2 _3145_ (.A1(_0044_),
    .A2(clknet_1_0__leaf__0531_),
    .B1(_0533_),
    .C1(\dut_0.U0_formal_verification.cbx_2__2_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0534_));
 sky130_fd_sc_hd__or2_2 _3146_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_2 _3147_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0536_));
 sky130_fd_sc_hd__and3_2 _3148_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0535_),
    .C(clknet_1_0__leaf__0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0537_));
 sky130_fd_sc_hd__nand2b_2 _3149_ (.A_N(clknet_1_1__leaf__0537_),
    .B(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0538_));
 sky130_fd_sc_hd__o211a_2 _3150_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0534_),
    .B1(_0538_),
    .C1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0539_));
 sky130_fd_sc_hd__inv_2 _4311__191 (.A(_1641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net426));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(net425),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0541_));
 sky130_fd_sc_hd__a31o_2 _3153_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0535_),
    .A3(clknet_1_1__leaf__0536_),
    .B1(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0542_));
 sky130_fd_sc_hd__o21a_2 _3154_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_9.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0543_));
 sky130_fd_sc_hd__and2_2 _3155_ (.A(clknet_1_0__leaf__0542_),
    .B(clknet_1_0__leaf__0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0544_));
 sky130_fd_sc_hd__a21bo_2 _3156_ (.A1(clknet_1_1__leaf__0542_),
    .A2(clknet_1_1__leaf__0543_),
    .B1_N(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0545_));
 sky130_fd_sc_hd__or2_1 _3157_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0546_));
 sky130_fd_sc_hd__and3_2 _3158_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0545_),
    .C(clknet_1_1__leaf__0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0547_));
 sky130_fd_sc_hd__a31o_2 _3159_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0545_),
    .A3(clknet_1_0__leaf__0546_),
    .B1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0548_));
 sky130_fd_sc_hd__nand2b_2 _3160_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0549_));
 sky130_fd_sc_hd__and3_2 _3161_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0548_),
    .C(clknet_1_0__leaf__0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0550_));
 sky130_fd_sc_hd__a31o_2 _3162_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0548_),
    .A3(clknet_1_1__leaf__0549_),
    .B1(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(net287),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_2 _3164_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.D ),
    .B(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _3165_ (.A(_0040_),
    .B(clknet_1_0__leaf__0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0554_));
 sky130_fd_sc_hd__nand3_2 _3166_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0551_),
    .C(clknet_1_1__leaf__0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0555_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(clknet_1_0__leaf__0555_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0556_));
 sky130_fd_sc_hd__mux4_2 _3168_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net408),
    .A2(_0556_),
    .A3(_0541_),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_0522_),
    .A1(_0557_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0558_));
 sky130_fd_sc_hd__nand2b_2 _3170_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2b_1 _3171_ (.A_N(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_8.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0560_));
 sky130_fd_sc_hd__and3_2 _3172_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.D ),
    .B(clknet_1_1__leaf__0559_),
    .C(clknet_1_1__leaf__0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0561_));
 sky130_fd_sc_hd__a31o_2 _3173_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.D ),
    .A2(clknet_1_0__leaf__0559_),
    .A3(clknet_1_0__leaf__0560_),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0562_));
 sky130_fd_sc_hd__nand2b_2 _3174_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0563_));
 sky130_fd_sc_hd__and3_2 _3175_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0562_),
    .C(clknet_1_0__leaf__0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0564_));
 sky130_fd_sc_hd__nand3_2 _3176_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0562_),
    .C(clknet_1_0__leaf__0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0565_));
 sky130_fd_sc_hd__a31o_2 _3177_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0562_),
    .A3(clknet_1_1__leaf__0563_),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0566_));
 sky130_fd_sc_hd__nand2b_2 _3178_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0567_));
 sky130_fd_sc_hd__and3_2 _3179_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0566_),
    .C(clknet_1_0__leaf__0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0568_));
 sky130_fd_sc_hd__a31o_2 _3180_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0566_),
    .A3(clknet_1_1__leaf__0567_),
    .B1(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0569_));
 sky130_fd_sc_hd__or2_2 _3181_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0570_));
 sky130_fd_sc_hd__and3_2 _3182_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0569_),
    .C(clknet_1_0__leaf__0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0571_));
 sky130_fd_sc_hd__nand3_2 _3183_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0569_),
    .C(clknet_1_1__leaf__0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0572_));
 sky130_fd_sc_hd__o21ai_1 _3184_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_8.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0547_),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0573_));
 sky130_fd_sc_hd__a21o_2 _3185_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_8.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0572_),
    .B1(_0573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0574_));
 sky130_fd_sc_hd__inv_2 _3704__64 (.A(_1067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net299));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(clknet_1_1__leaf__0558_),
    .A1(clknet_1_1__leaf__0574_),
    .S(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0576_));
 sky130_fd_sc_hd__or2_2 _3188_ (.A(_0047_),
    .B(_0576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__nand2b_2 _3189_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0577_));
 sky130_fd_sc_hd__o211a_2 _3190_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_0_.Q ),
    .A2(net334),
    .B1(_0577_),
    .C1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0578_));
 sky130_fd_sc_hd__inv_2 _2798__19 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net254));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(clknet_1_1__leaf__0525_),
    .A1(clknet_1_1__leaf__0578_),
    .S(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_2 _3193_ (.A(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_1_.Q ),
    .B(_0580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _3194_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(net324),
    .B1(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0581_));
 sky130_fd_sc_hd__a21o_2 _3195_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .B1(_0581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__nand2_1 _3196_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0582_));
 sky130_fd_sc_hd__o211a_2 _3197_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .A2(net298),
    .B1(_0582_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0583_));
 sky130_fd_sc_hd__a31o_1 _3198_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .A2(_0051_),
    .A3(net281),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0584_));
 sky130_fd_sc_hd__nand2b_2 _3199_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0585_));
 sky130_fd_sc_hd__o211a_2 _3200_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.Q ),
    .A2(net267),
    .B1(_0585_),
    .C1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0586_));
 sky130_fd_sc_hd__a21o_2 _3201_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0586_),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0587_));
 sky130_fd_sc_hd__a31o_2 _3202_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0569_),
    .A3(clknet_1_0__leaf__0570_),
    .B1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0588_));
 sky130_fd_sc_hd__nand2b_1 _3203_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0589_));
 sky130_fd_sc_hd__and3_2 _3204_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0588_),
    .C(clknet_1_0__leaf__0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0590_));
 sky130_fd_sc_hd__a31o_2 _3205_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0588_),
    .A3(clknet_1_1__leaf__0589_),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0591_));
 sky130_fd_sc_hd__nand2b_2 _3206_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0592_));
 sky130_fd_sc_hd__and3_2 _3207_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0591_),
    .C(clknet_1_0__leaf__0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0593_));
 sky130_fd_sc_hd__a31o_2 _3208_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0591_),
    .A3(clknet_1_1__leaf__0592_),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0594_));
 sky130_fd_sc_hd__nand2b_2 _3209_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0595_));
 sky130_fd_sc_hd__and3_2 _3210_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0594_),
    .C(clknet_1_1__leaf__0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0596_));
 sky130_fd_sc_hd__a31o_2 _3211_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0594_),
    .A3(clknet_1_0__leaf__0595_),
    .B1(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0597_));
 sky130_fd_sc_hd__or2_2 _3212_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0598_));
 sky130_fd_sc_hd__and3_2 _3213_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.ccff_head ),
    .B(clknet_1_1__leaf__0597_),
    .C(clknet_1_1__leaf__0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0599_));
 sky130_fd_sc_hd__a41o_2 _3214_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.ccff_head ),
    .A2(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_0_.Q ),
    .A3(clknet_1_0__leaf__0597_),
    .A4(clknet_1_0__leaf__0598_),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(clknet_1_0__leaf__0248_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0601_));
 sky130_fd_sc_hd__nand2_2 _3216_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_1_.Q ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0602_));
 sky130_fd_sc_hd__and2_2 _3217_ (.A(clknet_1_0__leaf__0600_),
    .B(clknet_1_0__leaf__0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_2 _3218_ (.A1(clknet_1_0__leaf__0600_),
    .A2(clknet_1_0__leaf__0602_),
    .B1(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0604_));
 sky130_fd_sc_hd__nand2_2 _3219_ (.A(_0054_),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_2 _3220_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0606_));
 sky130_fd_sc_hd__o211a_2 _3221_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_1_.Q ),
    .C1(_0606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .A1(clknet_1_1__leaf__0607_),
    .S(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0608_));
 sky130_fd_sc_hd__nand2_2 _3223_ (.A(\dut_0.U0_formal_verification.cby_0__1_.ccff_head ),
    .B(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _3224_ (.A(_0055_),
    .B(clknet_1_1__leaf__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0610_));
 sky130_fd_sc_hd__o211a_1 _3225_ (.A1(_0055_),
    .A2(clknet_1_0__leaf__0528_),
    .B1(_0610_),
    .C1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0611_));
 sky130_fd_sc_hd__a31o_1 _3226_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_1_.Q ),
    .A2(_0057_),
    .A3(clknet_1_0__leaf__0611_),
    .B1(\dut_0.U0_formal_verification.cbx_1__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0612_));
 sky130_fd_sc_hd__a31o_1 _3227_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ),
    .A2(_0604_),
    .A3(_0605_),
    .B1(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0613_));
 sky130_fd_sc_hd__nand2b_2 _3228_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0614_));
 sky130_fd_sc_hd__o211a_2 _3229_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_0_.Q ),
    .A2(net262),
    .B1(_0614_),
    .C1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0615_));
 sky130_fd_sc_hd__o21ai_2 _3230_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0615_),
    .B1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0616_));
 sky130_fd_sc_hd__a21o_2 _3231_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .B1(_0616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0617_));
 sky130_fd_sc_hd__nor2_2 _3232_ (.A(_0054_),
    .B(clknet_1_0__leaf__0617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0618_));
 sky130_fd_sc_hd__a31o_2 _3233_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.D ),
    .A2(clknet_1_1__leaf__0252_),
    .A3(clknet_1_1__leaf__0253_),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0619_));
 sky130_fd_sc_hd__nand2b_2 _3234_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0620_));
 sky130_fd_sc_hd__and3_2 _3235_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.D ),
    .B(clknet_1_0__leaf__0619_),
    .C(clknet_1_0__leaf__0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0621_));
 sky130_fd_sc_hd__a31o_2 _3236_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.D ),
    .A2(clknet_1_1__leaf__0619_),
    .A3(clknet_1_1__leaf__0620_),
    .B1(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0622_));
 sky130_fd_sc_hd__o21a_1 _3237_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0531_),
    .B1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0623_));
 sky130_fd_sc_hd__and2_2 _3238_ (.A(clknet_1_1__leaf__0622_),
    .B(clknet_1_0__leaf__0623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0624_));
 sky130_fd_sc_hd__nand2_2 _3239_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0625_));
 sky130_fd_sc_hd__o211a_2 _3240_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .A2(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_1_.Q ),
    .C1(_0625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0626_));
 sky130_fd_sc_hd__o21ai_2 _3241_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0626_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0627_));
 sky130_fd_sc_hd__a21o_2 _3242_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .B1(_0627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0628_));
 sky130_fd_sc_hd__nor2_2 _3243_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0629_));
 sky130_fd_sc_hd__a21o_2 _3244_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .B1(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0630_));
 sky130_fd_sc_hd__o221a_2 _3245_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0628_),
    .B1(_0629_),
    .B2(_0630_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0631_));
 sky130_fd_sc_hd__a211oi_2 _3246_ (.A1(_0054_),
    .A2(clknet_1_0__leaf__0624_),
    .B1(_0618_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0632_));
 sky130_fd_sc_hd__o21ai_2 _3247_ (.A1(_0631_),
    .A2(_0632_),
    .B1(\dut_0.U0_formal_verification.cbx_1__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _3248_ (.A(clknet_1_1__leaf__0613_),
    .B(clknet_1_1__leaf__0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0634_));
 sky130_fd_sc_hd__o21ai_2 _3249_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ),
    .A2(net253),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0635_));
 sky130_fd_sc_hd__a31o_2 _3250_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0613_),
    .A3(clknet_1_0__leaf__0633_),
    .B1(_0635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0636_));
 sky130_fd_sc_hd__a21o_2 _3251_ (.A1(_0587_),
    .A2(_0636_),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0637_));
 sky130_fd_sc_hd__nand2b_2 _3252_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0638_));
 sky130_fd_sc_hd__o211a_2 _3253_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_0_.Q ),
    .A2(net259),
    .B1(_0638_),
    .C1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_2 _3254_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0640_));
 sky130_fd_sc_hd__nor2_4 _3255_ (.A(_0053_),
    .B(_0640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0641_));
 sky130_fd_sc_hd__a31oi_4 _3256_ (.A1(_0053_),
    .A2(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_1_.Q ),
    .A3(clknet_1_0__leaf__0639_),
    .B1(_0641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0642_));
 sky130_fd_sc_hd__inv_2 _2790__45 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net280));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_2 _3259_ (.A0(clknet_1_0__leaf__0233_),
    .A1(net278),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .A3(_0644_),
    .S0(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0645_));
 sky130_fd_sc_hd__o21a_2 _3260_ (.A1(_0059_),
    .A2(_0645_),
    .B1(_0637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0646_));
 sky130_fd_sc_hd__nand2b_1 _3261_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0647_));
 sky130_fd_sc_hd__o211a_1 _3262_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0646_),
    .B1(_0647_),
    .C1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(clknet_1_1__leaf__0648_),
    .A1(clknet_1_0__leaf__0593_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_2 _3264_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_1_.Q ),
    .B(_0649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0650_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(clknet_1_0__leaf__0642_),
    .A1(clknet_1_0__leaf__0650_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_2 _3266_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0652_));
 sky130_fd_sc_hd__o211a_2 _3267_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .A2(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_1_.Q ),
    .C1(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0653_));
 sky130_fd_sc_hd__nand2_2 _3268_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0654_));
 sky130_fd_sc_hd__o211a_2 _3269_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0653_),
    .B1(_0654_),
    .C1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0655_));
 sky130_fd_sc_hd__inv_2 _3340__184 (.A(_0724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net419));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(net418),
    .A1(clknet_1_0__leaf__0259_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0657_));
 sky130_fd_sc_hd__a21o_2 _3272_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .A2(_0657_),
    .B1(_0051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0658_));
 sky130_fd_sc_hd__a21o_2 _3273_ (.A1(_0050_),
    .A2(_0651_),
    .B1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0659_));
 sky130_fd_sc_hd__nand2_2 _3274_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0660_));
 sky130_fd_sc_hd__o211a_2 _3275_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_1_.Q ),
    .C1(_0660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .A1(clknet_1_1__leaf__0661_),
    .S(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0662_));
 sky130_fd_sc_hd__and2_2 _3277_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_1_.Q ),
    .B(_0662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0663_));
 sky130_fd_sc_hd__nand2b_1 _3278_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0664_));
 sky130_fd_sc_hd__o211a_2 _3279_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0586_),
    .B1(_0664_),
    .C1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0665_));
 sky130_fd_sc_hd__inv_2 _2808__67 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net302));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(clknet_1_1__leaf__0665_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0667_));
 sky130_fd_sc_hd__and2_2 _3282_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0668_));
 sky130_fd_sc_hd__nand2_2 _3283_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_2 _3284_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0670_));
 sky130_fd_sc_hd__o211a_2 _3285_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .A2(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_1_.Q ),
    .C1(_0670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0671_));
 sky130_fd_sc_hd__inv_2 _2811__98 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net333));
 sky130_fd_sc_hd__mux4_2 _3287_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .A1(net332),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .A3(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_2 _3288_ (.A(_0052_),
    .B(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0674_));
 sky130_fd_sc_hd__a31o_2 _3289_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_1_.Q ),
    .A2(_0052_),
    .A3(clknet_1_1__leaf__0663_),
    .B1(_0674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0675_));
 sky130_fd_sc_hd__nand2b_1 _3290_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0676_));
 sky130_fd_sc_hd__o211a_4 _3291_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0578_),
    .B1(_0676_),
    .C1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0677_));
 sky130_fd_sc_hd__nand2b_1 _3292_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0678_));
 sky130_fd_sc_hd__o211a_4 _3293_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0677_),
    .B1(_0678_),
    .C1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(net320),
    .A1(clknet_1_0__leaf__0679_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0680_));
 sky130_fd_sc_hd__and2_2 _3295_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_1_.Q ),
    .B(_0680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0681_));
 sky130_fd_sc_hd__inv_2 _3750__168 (.A(_1111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net403));
 sky130_fd_sc_hd__or3_2 _3297_ (.A(_0050_),
    .B(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ),
    .C(net402),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0683_));
 sky130_fd_sc_hd__or3b_2 _3298_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .B(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ),
    .C_N(clknet_1_1__leaf__0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0684_));
 sky130_fd_sc_hd__and3_2 _3299_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.D ),
    .B(_0683_),
    .C(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0685_));
 sky130_fd_sc_hd__o2bb2a_4 _3300_ (.A1_N(_0685_),
    .A2_N(_0659_),
    .B1(_0584_),
    .B2(_0583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(clknet_1_0__leaf__0561_),
    .A1(clknet_1_1__leaf__0544_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0687_));
 sky130_fd_sc_hd__and2_2 _3302_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.D ),
    .B(_0687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_4 _3303_ (.A0(_0686_),
    .A1(clknet_1_1__leaf__0688_),
    .S(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_8 _3304_ (.A(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_1_.Q ),
    .B(_0689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__nand2b_2 _3305_ (.A_N(clknet_1_1__leaf__0525_),
    .B(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0690_));
 sky130_fd_sc_hd__o211a_2 _3306_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0544_),
    .B1(_0690_),
    .C1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0691_));
 sky130_fd_sc_hd__o21ai_2 _3307_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0692_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(clknet_1_0__leaf__0624_),
    .A1(_0686_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0693_));
 sky130_fd_sc_hd__o22a_2 _3309_ (.A1(_0691_),
    .A2(_0692_),
    .B1(_0693_),
    .B2(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0694_));
 sky130_fd_sc_hd__nand2_1 _3310_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0695_));
 sky130_fd_sc_hd__o211a_1 _3311_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ),
    .B1(_0695_),
    .C1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0696_));
 sky130_fd_sc_hd__a31o_1 _3312_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .A2(_0061_),
    .A3(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ),
    .B1(_0696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_2 _3313_ (.A0(_0697_),
    .A1(_0694_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0698_));
 sky130_fd_sc_hd__o21ai_1 _3314_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0677_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0699_));
 sky130_fd_sc_hd__a21o_2 _3315_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .B1(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .A1(clknet_1_0__leaf__0550_),
    .S(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0701_));
 sky130_fd_sc_hd__and2_4 _3317_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.D ),
    .B(_0701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(clknet_1_1__leaf__0224_),
    .A1(clknet_1_1__leaf__0702_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_4 _3319_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.D ),
    .B(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0704_));
 sky130_fd_sc_hd__mux4_2 _3320_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .A1(clknet_1_0__leaf__0700_),
    .A2(clknet_1_1__leaf__0704_),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .A1(net407),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(_0706_),
    .A1(_0705_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_2 _3323_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0708_));
 sky130_fd_sc_hd__o211a_2 _3324_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_1_.Q ),
    .C1(_0708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _3325_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .A1(clknet_1_1__leaf__0709_),
    .S(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0710_));
 sky130_fd_sc_hd__and2_1 _3326_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0711_));
 sky130_fd_sc_hd__a31o_1 _3327_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_1_.Q ),
    .A2(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_1_.Q ),
    .A3(clknet_1_1__leaf__0710_),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .A1(clknet_1_0__leaf__0679_),
    .S(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0713_));
 sky130_fd_sc_hd__and2_2 _3329_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_1_.Q ),
    .B(_0713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_2 _3330_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0715_));
 sky130_fd_sc_hd__o211a_2 _3331_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0714_),
    .B1(_0715_),
    .C1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0716_));
 sky130_fd_sc_hd__o21ai_1 _3332_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_1_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0717_));
 sky130_fd_sc_hd__o21ai_2 _3333_ (.A1(_0716_),
    .A2(_0717_),
    .B1(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0718_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(clknet_1_0__leaf__0718_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0719_));
 sky130_fd_sc_hd__inv_2 _2805__141 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net376));
 sky130_fd_sc_hd__nor2_1 _3336_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_2_.Q ),
    .B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0721_));
 sky130_fd_sc_hd__a221o_2 _3337_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_2_.Q ),
    .A2(net375),
    .B1(_0721_),
    .B2(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0722_));
 sky130_fd_sc_hd__a21bo_2 _3338_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_3_.Q ),
    .A2(_0707_),
    .B1_N(_0722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(clknet_1_1__leaf__0709_),
    .A1(clknet_1_1__leaf__0661_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0724_));
 sky130_fd_sc_hd__inv_2 _3391__185 (.A(_0772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net420));
 sky130_fd_sc_hd__mux4_2 _3341_ (.A0(clknet_1_0__leaf__0617_),
    .A1(net401),
    .A2(net419),
    .A3(clknet_1_0__leaf__0723_),
    .S0(_0060_),
    .S1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0727_));
 sky130_fd_sc_hd__a31o_2 _3343_ (.A1(_0060_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .A3(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_2_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0728_));
 sky130_fd_sc_hd__a21oi_2 _3344_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_1_.Q ),
    .A2(_0727_),
    .B1(_0728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0729_));
 sky130_fd_sc_hd__a21oi_2 _3345_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.D ),
    .A2(_0726_),
    .B1(_0729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0730_));
 sky130_fd_sc_hd__mux4_2 _3346_ (.A0(clknet_1_0__leaf__0730_),
    .A1(clknet_1_1__leaf__0698_),
    .A2(clknet_1_1__leaf__0561_),
    .A3(clknet_1_1__leaf__0221_),
    .S0(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0731_));
 sky130_fd_sc_hd__nand2b_1 _3347_ (.A_N(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ),
    .B(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0732_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0733_));
 sky130_fd_sc_hd__a2bb2oi_1 _3349_ (.A1_N(net252),
    .A2_N(_0732_),
    .B1(_0733_),
    .B2(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0734_));
 sky130_fd_sc_hd__nor2_1 _3350_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0735_));
 sky130_fd_sc_hd__a211o_2 _3351_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0233_),
    .B1(_0735_),
    .C1(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _3352_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .A1(clknet_1_0__leaf__0702_),
    .S(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0737_));
 sky130_fd_sc_hd__and2_2 _3353_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_1_.Q ),
    .B(_0737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0738_));
 sky130_fd_sc_hd__nand2_1 _3354_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ),
    .B(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0739_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(clknet_1_0__leaf__0607_),
    .A1(clknet_1_0__leaf__0738_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0740_));
 sky130_fd_sc_hd__o221a_2 _3356_ (.A1(net277),
    .A2(_0732_),
    .B1(_0739_),
    .B2(_0740_),
    .C1(\dut_0.U0_formal_verification.cby_0__2_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0741_));
 sky130_fd_sc_hd__a2bb2o_2 _3357_ (.A1_N(\dut_0.U0_formal_verification.cby_0__2_.ccff_head ),
    .A2_N(_0734_),
    .B1(_0736_),
    .B2(_0741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0742_));
 sky130_fd_sc_hd__nand2_1 _3358_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_16.DFF_0_.Q ),
    .B(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0743_));
 sky130_fd_sc_hd__o211ai_2 _3359_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_16.DFF_0_.Q ),
    .A2(net290),
    .B1(_0743_),
    .C1(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0744_));
 sky130_fd_sc_hd__inv_2 _3186__61 (.A(clknet_1_0__leaf__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net296));
 sky130_fd_sc_hd__nand2_2 _3361_ (.A(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0746_));
 sky130_fd_sc_hd__o2111a_2 _3362_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0742_),
    .B1(_0746_),
    .C1(_0062_),
    .D1(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0747_));
 sky130_fd_sc_hd__a21oi_2 _3363_ (.A1(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_2_.Q ),
    .A2(_0731_),
    .B1(_0747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__mux4_2 _3364_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0748_));
 sky130_fd_sc_hd__a21o_1 _3365_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0749_));
 sky130_fd_sc_hd__nand3b_1 _3366_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ),
    .C(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0750_));
 sky130_fd_sc_hd__o21ba_1 _3367_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .B1_N(\dut_0.U0_formal_verification.cbx_1__0_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(clknet_1_0__leaf__0558_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(net417),
    .A1(_0752_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_2 _3370_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ),
    .B(_0753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0754_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(clknet_1_0__leaf__0571_),
    .A1(clknet_1_0__leaf__0247_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0755_));
 sky130_fd_sc_hd__o211a_2 _3372_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ),
    .A2(_0755_),
    .B1(_0754_),
    .C1(\dut_0.U0_formal_verification.cbx_1__0_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0756_));
 sky130_fd_sc_hd__a31o_2 _3373_ (.A1(_0749_),
    .A2(_0750_),
    .A3(_0751_),
    .B1(_0756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0757_));
 sky130_fd_sc_hd__nand2_1 _3374_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0758_));
 sky130_fd_sc_hd__o2111a_1 _3375_ (.A1(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0757_),
    .B1(_0758_),
    .C1(_0063_),
    .D1(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0759_));
 sky130_fd_sc_hd__o21ba_2 _3376_ (.A1(_0063_),
    .A2(_0748_),
    .B1_N(_0759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nor2_2 _3377_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0760_));
 sky130_fd_sc_hd__a211o_2 _3378_ (.A1(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .B1(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_2_.Q ),
    .C1(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0761_));
 sky130_fd_sc_hd__mux4_1 _3379_ (.A0(clknet_1_1__leaf__0202_),
    .A1(clknet_1_1__leaf__0603_),
    .A2(net376),
    .A3(clknet_1_0__leaf_net35),
    .S0(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_0_.Q ),
    .S1(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0762_));
 sky130_fd_sc_hd__o2bb2a_2 _3380_ (.A1_N(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_2_.Q ),
    .A2_N(_0762_),
    .B1(_0761_),
    .B2(_0760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2b_2 _3381_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0763_));
 sky130_fd_sc_hd__o211a_2 _3382_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_0_.Q ),
    .A2(net344),
    .B1(_0763_),
    .C1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(clknet_1_1__leaf__0764_),
    .A1(clknet_1_1__leaf__0221_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0765_));
 sky130_fd_sc_hd__and2_2 _3384_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.D ),
    .B(_0765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(clknet_1_1__leaf__0624_),
    .A1(clknet_1_0__leaf__0766_),
    .S(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0767_));
 sky130_fd_sc_hd__and3b_2 _3386_ (.A_N(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_2_.Q ),
    .B(_0767_),
    .C(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0768_));
 sky130_fd_sc_hd__a21o_2 _3387_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0586_),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_2 _3388_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0770_));
 sky130_fd_sc_hd__a311o_2 _3389_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0600_),
    .A3(clknet_1_1__leaf__0602_),
    .B1(_0770_),
    .C1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0772_));
 sky130_fd_sc_hd__inv_2 _2807__186 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net421));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(net17),
    .A1(net420),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_2 _3393_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ),
    .B(_0774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0775_));
 sky130_fd_sc_hd__a21oi_2 _3394_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0766_),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0776_));
 sky130_fd_sc_hd__and2_2 _3395_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .A1(_0777_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0778_));
 sky130_fd_sc_hd__nor2_2 _3397_ (.A(_0776_),
    .B(_0778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0779_));
 sky130_fd_sc_hd__o21ai_2 _3398_ (.A1(_0067_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0780_));
 sky130_fd_sc_hd__a41o_2 _3399_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_1_.Q ),
    .A2(_0067_),
    .A3(clknet_1_0__leaf__0551_),
    .A4(clknet_1_0__leaf__0554_),
    .B1(_0780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0781_));
 sky130_fd_sc_hd__o211a_2 _3400_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0233_),
    .B1(_0781_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0783_));
 sky130_fd_sc_hd__o21ai_2 _3402_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ),
    .A2(_0783_),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0784_));
 sky130_fd_sc_hd__o22a_2 _3403_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.D ),
    .A2(_0779_),
    .B1(_0782_),
    .B2(_0784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0785_));
 sky130_fd_sc_hd__o21ai_2 _3404_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0565_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0786_));
 sky130_fd_sc_hd__a21o_2 _3405_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0785_),
    .B1(_0786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0787_));
 sky130_fd_sc_hd__a31o_2 _3406_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0222_),
    .A3(clknet_1_0__leaf__0223_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0788_));
 sky130_fd_sc_hd__and3b_2 _3407_ (.A_N(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.D ),
    .B(_0787_),
    .C(_0788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0789_));
 sky130_fd_sc_hd__a31oi_2 _3408_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.D ),
    .A2(clknet_1_1__leaf__0771_),
    .A3(clknet_1_1__leaf__0775_),
    .B1(clknet_1_1__leaf__0789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0790_));
 sky130_fd_sc_hd__a311o_2 _3409_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.D ),
    .A2(clknet_1_0__leaf__0771_),
    .A3(clknet_1_0__leaf__0775_),
    .B1(clknet_1_0__leaf__0789_),
    .C1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0791_));
 sky130_fd_sc_hd__nand2b_2 _3410_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0792_));
 sky130_fd_sc_hd__and3_2 _3411_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0791_),
    .C(clknet_1_0__leaf__0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0793_));
 sky130_fd_sc_hd__a31o_2 _3412_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0791_),
    .A3(clknet_1_1__leaf__0792_),
    .B1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0794_));
 sky130_fd_sc_hd__nand2_2 _3413_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_17.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0795_));
 sky130_fd_sc_hd__nand3_2 _3414_ (.A(\dut_0.U0_formal_verification.cbx_2__1_.ccff_head ),
    .B(clknet_1_0__leaf__0794_),
    .C(clknet_1_0__leaf__0795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0796_));
 sky130_fd_sc_hd__a31o_2 _3415_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0622_),
    .A3(clknet_1_1__leaf__0623_),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0797_));
 sky130_fd_sc_hd__a41o_2 _3416_ (.A1(\dut_0.U0_formal_verification.cbx_2__1_.ccff_head ),
    .A2(_0068_),
    .A3(clknet_1_1__leaf__0794_),
    .A4(clknet_1_1__leaf__0795_),
    .B1(_0797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0617_),
    .S(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_2 _3418_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ),
    .A2(_0799_),
    .B1(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0800_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(net258),
    .A1(clknet_1_1__leaf__0603_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0801_));
 sky130_fd_sc_hd__a22o_2 _3420_ (.A1(_0798_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_2 _3422_ (.A(_0066_),
    .B(_0803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0804_));
 sky130_fd_sc_hd__mux2_2 _3423_ (.A0(_0804_),
    .A1(_0802_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(clknet_1_0__leaf__0257_),
    .A1(clknet_1_0__leaf__0537_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0806_));
 sky130_fd_sc_hd__mux4_2 _3425_ (.A0(net330),
    .A1(clknet_1_0__leaf__0675_),
    .A2(clknet_1_0__leaf__0805_),
    .A3(_0806_),
    .S0(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_1 _3427_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_2_.Q ),
    .B(clknet_1_1__leaf_net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0809_));
 sky130_fd_sc_hd__a22o_2 _3428_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_2_.Q ),
    .A2(_0808_),
    .B1(_0809_),
    .B2(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_2 _3429_ (.A0(_0810_),
    .A1(_0807_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0811_));
 sky130_fd_sc_hd__or2_2 _3430_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0812_));
 sky130_fd_sc_hd__o211a_2 _3431_ (.A1(_0069_),
    .A2(clknet_1_1__leaf__0811_),
    .B1(clknet_1_1__leaf__0812_),
    .C1(\dut_0.U0_formal_verification.sb_0__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0813_));
 sky130_fd_sc_hd__o2111a_2 _3432_ (.A1(_0069_),
    .A2(clknet_1_1__leaf__0811_),
    .B1(clknet_1_0__leaf__0812_),
    .C1(\dut_0.U0_formal_verification.sb_0__1_.ccff_head ),
    .D1(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0814_));
 sky130_fd_sc_hd__a21bo_2 _3433_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0738_),
    .B1_N(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0815_));
 sky130_fd_sc_hd__o21ai_2 _3434_ (.A1(_0814_),
    .A2(_0815_),
    .B1(_0769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0816_));
 sky130_fd_sc_hd__mux4_2 _3435_ (.A0(clknet_1_1__leaf__0617_),
    .A1(clknet_1_1__leaf__0642_),
    .A2(clknet_1_1__leaf__0816_),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0817_));
 sky130_fd_sc_hd__inv_2 _3296__166 (.A(clknet_1_0__leaf__0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net401));
 sky130_fd_sc_hd__a21oi_2 _3437_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_2_.Q ),
    .A2(net400),
    .B1(_0768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2b_1 _3438_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0819_));
 sky130_fd_sc_hd__o211a_1 _3439_ (.A1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0757_),
    .B1(_0819_),
    .C1(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0820_));
 sky130_fd_sc_hd__a21o_1 _3440_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0820_),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_2 _3441_ (.A0(clknet_1_0__leaf__0578_),
    .A1(clknet_1_0__leaf__0607_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0822_));
 sky130_fd_sc_hd__o21ai_4 _3442_ (.A1(_0822_),
    .A2(_0151_),
    .B1(_0821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__a21o_1 _3443_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0590_),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0824_));
 sky130_fd_sc_hd__and3b_1 _3445_ (.A_N(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_1_.Q ),
    .B(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_2_.Q ),
    .C(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0825_));
 sky130_fd_sc_hd__a21o_2 _3446_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_1_.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(clknet_1_1__leaf__0702_),
    .A1(net347),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0827_));
 sky130_fd_sc_hd__mux4_2 _3448_ (.A0(clknet_1_0__leaf__0785_),
    .A1(clknet_1_0__leaf__0603_),
    .A2(net297),
    .A3(_0827_),
    .S0(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(_0826_),
    .A1(_0828_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .A1(clknet_1_1__leaf__0829_),
    .S(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0830_));
 sky130_fd_sc_hd__and2_2 _3451_ (.A(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_1_.Q ),
    .B(_0830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(clknet_1_1__leaf__0831_),
    .A1(clknet_1_0__leaf__0661_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0832_));
 sky130_fd_sc_hd__o21ai_4 _3453_ (.A1(_0832_),
    .A2(_0153_),
    .B1(_0823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__o21a_2 _3454_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_8.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0833_));
 sky130_fd_sc_hd__o21ai_4 _3455_ (.A1(_0146_),
    .A2(clknet_1_1__leaf__0738_),
    .B1(_0833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand2b_2 _3456_ (.A_N(clknet_1_0__leaf__0596_),
    .B(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0834_));
 sky130_fd_sc_hd__o21a_2 _3457_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0621_),
    .B1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0835_));
 sky130_fd_sc_hd__a22o_2 _3458_ (.A1(_0112_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .B1(_0834_),
    .B2(_0835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _3459_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(net266),
    .A1(clknet_1_1__leaf__0675_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0838_));
 sky130_fd_sc_hd__mux4_2 _3461_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf__0700_),
    .A2(clknet_1_1__leaf__0704_),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0839_));
 sky130_fd_sc_hd__nand2_2 _3462_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ),
    .B(_0839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0840_));
 sky130_fd_sc_hd__o21a_2 _3463_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ),
    .A2(_0838_),
    .B1(_0840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .A1(clknet_1_1__leaf__0574_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0842_));
 sky130_fd_sc_hd__inv_2 _3151__188 (.A(clknet_1_1__leaf__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net423));
 sky130_fd_sc_hd__nor2_2 _3466_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0844_));
 sky130_fd_sc_hd__a22o_2 _3467_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ),
    .A2(net422),
    .B1(_0844_),
    .B2(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_2 _3468_ (.A0(_0845_),
    .A1(_0841_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(clknet_1_1__leaf__0193_),
    .A1(clknet_1_1__leaf__0846_),
    .S(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0847_));
 sky130_fd_sc_hd__nor2_2 _3470_ (.A(_0112_),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0848_));
 sky130_fd_sc_hd__mux4_2 _3471_ (.A0(_0848_),
    .A1(_0847_),
    .A2(_0837_),
    .A3(_0836_),
    .S0(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0849_));
 sky130_fd_sc_hd__o21a_1 _3472_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.Q ),
    .A2(net367),
    .B1(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0850_));
 sky130_fd_sc_hd__o21ai_2 _3473_ (.A1(_0150_),
    .A2(clknet_1_0__leaf__0849_),
    .B1(_0850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__o21ai_1 _3474_ (.A1(_0148_),
    .A2(clknet_1_1__leaf__0742_),
    .B1(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0851_));
 sky130_fd_sc_hd__a21o_2 _3475_ (.A1(_0148_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .B1(_0851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(clknet_1_0__leaf__0816_),
    .A1(net38),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0852_));
 sky130_fd_sc_hd__a21oi_2 _3477_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0688_),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0853_));
 sky130_fd_sc_hd__a211oi_1 _3478_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ),
    .A2(_0852_),
    .B1(_0853_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2_2 _3479_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0855_));
 sky130_fd_sc_hd__a211o_2 _3480_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0624_),
    .B1(_0855_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0856_));
 sky130_fd_sc_hd__o21ai_2 _3481_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0655_),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0857_));
 sky130_fd_sc_hd__a21o_2 _3482_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0259_),
    .B1(_0857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0858_));
 sky130_fd_sc_hd__o211ai_2 _3483_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0617_),
    .B1(_0858_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0859_));
 sky130_fd_sc_hd__a31o_1 _3484_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_3_.Q ),
    .A2(_0856_),
    .A3(_0859_),
    .B1(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0860_));
 sky130_fd_sc_hd__inv_2 _2818__109 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net344));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(clknet_1_1__leaf__0704_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0862_));
 sky130_fd_sc_hd__inv_2 _3872__144 (.A(_1227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net379));
 sky130_fd_sc_hd__mux4_2 _3488_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .A1(net366),
    .A2(clknet_1_1__leaf__0860_),
    .A3(net378),
    .S0(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(net286),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0865_));
 sky130_fd_sc_hd__nor2_2 _3490_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_2_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0866_));
 sky130_fd_sc_hd__a22o_2 _3491_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_2_.Q ),
    .A2(_0865_),
    .B1(_0866_),
    .B2(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_2 _3492_ (.A0(_0867_),
    .A1(_0864_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0868_));
 sky130_fd_sc_hd__o21ai_2 _3493_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0868_),
    .B1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0869_));
 sky130_fd_sc_hd__a21o_2 _3494_ (.A1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .B1(_0869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__a21o_1 _3495_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_0_.Q ),
    .A2(_0198_),
    .B1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0870_));
 sky130_fd_sc_hd__nand2_2 _3496_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0871_));
 sky130_fd_sc_hd__o211a_2 _3497_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0593_),
    .B1(_0871_),
    .C1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0872_));
 sky130_fd_sc_hd__a31o_1 _3498_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .A2(_0115_),
    .A3(clknet_1_1__leaf__0254_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0873_));
 sky130_fd_sc_hd__or3b_2 _3499_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ),
    .B(clknet_1_0__leaf__0675_),
    .C_N(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .A1(_0875_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0876_));
 sky130_fd_sc_hd__or2_2 _3502_ (.A(_0115_),
    .B(_0876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0877_));
 sky130_fd_sc_hd__o311a_2 _3503_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .A2(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ),
    .A3(clknet_1_1__leaf__0805_),
    .B1(_0874_),
    .C1(_0877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0878_));
 sky130_fd_sc_hd__o22a_2 _3504_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0878_),
    .B2(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0879_));
 sky130_fd_sc_hd__nand2_1 _3505_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_0_.Q ),
    .B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0880_));
 sky130_fd_sc_hd__o211a_2 _3506_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0879_),
    .B1(_0880_),
    .C1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0881_));
 sky130_fd_sc_hd__nand2b_2 _3507_ (.A_N(clknet_1_0__leaf__0568_),
    .B(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0882_));
 sky130_fd_sc_hd__o211a_2 _3508_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0881_),
    .B1(_0882_),
    .C1(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0883_));
 sky130_fd_sc_hd__mux4_1 _3509_ (.A0(clknet_1_0__leaf__0883_),
    .A1(clknet_1_1__leaf__0681_),
    .A2(net276),
    .A3(_0190_),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_0_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(net296),
    .A1(clknet_1_1__leaf__0675_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0885_));
 sky130_fd_sc_hd__nand2_1 _3511_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0886_));
 sky130_fd_sc_hd__o21ai_2 _3512_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0816_),
    .B1(_0886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0887_));
 sky130_fd_sc_hd__and2_2 _3513_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0888_));
 sky130_fd_sc_hd__mux4_2 _3514_ (.A0(_0888_),
    .A1(_0887_),
    .A2(_0885_),
    .A3(_0884_),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0890_));
 sky130_fd_sc_hd__mux4_2 _3516_ (.A0(clknet_1_0__leaf_net35),
    .A1(clknet_1_1__leaf__0889_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .A3(_0890_),
    .S0(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0891_));
 sky130_fd_sc_hd__a21oi_1 _3517_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0677_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0892_));
 sky130_fd_sc_hd__nor2_2 _3518_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0893_));
 sky130_fd_sc_hd__a311o_2 _3519_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ),
    .A2(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_2_.Q ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .B1(_0892_),
    .C1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0894_));
 sky130_fd_sc_hd__a2bb2o_2 _3520_ (.A1_N(_0893_),
    .A2_N(_0894_),
    .B1(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.D ),
    .B2(_0891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0895_));
 sky130_fd_sc_hd__nand2b_2 _3521_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0896_));
 sky130_fd_sc_hd__o211a_2 _3522_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0895_),
    .B1(_0896_),
    .C1(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(clknet_1_1__leaf__0897_),
    .A1(clknet_1_0__leaf__0596_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0898_));
 sky130_fd_sc_hd__o21ai_2 _3524_ (.A1(_0156_),
    .A2(_0898_),
    .B1(_0870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(clknet_1_0__leaf__0661_),
    .A1(clknet_1_0__leaf__0221_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0899_));
 sky130_fd_sc_hd__and2_2 _3526_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0900_));
 sky130_fd_sc_hd__nand2_2 _3527_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_1_.Q ),
    .B(clknet_1_1__leaf__0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_2 _3528_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0902_));
 sky130_fd_sc_hd__a211o_2 _3529_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_0902_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0904_));
 sky130_fd_sc_hd__inv_2 _3555__78 (.A(_0928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net313));
 sky130_fd_sc_hd__a21oi_2 _3532_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .A2(net312),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0906_));
 sky130_fd_sc_hd__mux4_2 _3533_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_0__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0907_));
 sky130_fd_sc_hd__a22o_2 _3534_ (.A1(_0903_),
    .A2(_0906_),
    .B1(_0907_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _3535_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0909_));
 sky130_fd_sc_hd__or3b_2 _3536_ (.A(_0909_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0910_));
 sky130_fd_sc_hd__mux4_2 _3537_ (.A0(clknet_1_0__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0911_));
 sky130_fd_sc_hd__inv_2 _3548__123 (.A(_0921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net358));
 sky130_fd_sc_hd__a21oi_2 _3539_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .A2(net357),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0913_));
 sky130_fd_sc_hd__a22o_2 _3540_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .A2(_0908_),
    .B1(_0910_),
    .B2(_0913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0914_));
 sky130_fd_sc_hd__mux4_2 _3541_ (.A0(clknet_1_0__leaf__0901_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0915_));
 sky130_fd_sc_hd__mux4_2 _3542_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_1__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0916_));
 sky130_fd_sc_hd__or2_2 _3543_ (.A(_0072_),
    .B(_0916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0917_));
 sky130_fd_sc_hd__o211a_2 _3544_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .A2(_0915_),
    .B1(_0917_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0919_));
 sky130_fd_sc_hd__or3_2 _3546_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .B(_0072_),
    .C(_0919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0920_));
 sky130_fd_sc_hd__mux4_2 _3547_ (.A0(clknet_1_1__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0921_));
 sky130_fd_sc_hd__inv_2 _3562__124 (.A(_0935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net359));
 sky130_fd_sc_hd__a21oi_2 _3549_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .A2(net358),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0923_));
 sky130_fd_sc_hd__a21oi_2 _3550_ (.A1(_0920_),
    .A2(_0923_),
    .B1(_0918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0924_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_1__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0925_));
 sky130_fd_sc_hd__nor2_2 _3552_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0926_));
 sky130_fd_sc_hd__a211o_2 _3553_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_0926_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0928_));
 sky130_fd_sc_hd__inv_2 _3570__79 (.A(_0943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net314));
 sky130_fd_sc_hd__a21oi_2 _3556_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .A2(net313),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0930_));
 sky130_fd_sc_hd__mux4_2 _3557_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_0__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0931_));
 sky130_fd_sc_hd__a22o_2 _3558_ (.A1(_0927_),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0933_));
 sky130_fd_sc_hd__or3b_2 _3560_ (.A(_0933_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0934_));
 sky130_fd_sc_hd__mux4_2 _3561_ (.A0(clknet_1_0__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0935_));
 sky130_fd_sc_hd__inv_2 _3911__125 (.A(_1263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net360));
 sky130_fd_sc_hd__a21oi_2 _3563_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .A2(net359),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0937_));
 sky130_fd_sc_hd__a22o_2 _3564_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .A2(_0932_),
    .B1(_0934_),
    .B2(_0937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_1__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(_0925_),
    .A1(_0939_),
    .S(clknet_1_0__leaf__0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_2 _3567_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0941_));
 sky130_fd_sc_hd__a211o_2 _3568_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_0941_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0943_));
 sky130_fd_sc_hd__inv_2 _3895__80 (.A(_1247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net315));
 sky130_fd_sc_hd__a21oi_2 _3571_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .A2(net314),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0945_));
 sky130_fd_sc_hd__mux4_2 _3572_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_1__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0946_));
 sky130_fd_sc_hd__a22o_2 _3573_ (.A1(_0942_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0948_));
 sky130_fd_sc_hd__or3b_2 _3575_ (.A(_0948_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0949_));
 sky130_fd_sc_hd__mux4_2 _3576_ (.A0(clknet_1_1__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0950_));
 sky130_fd_sc_hd__inv_2 _3577_ (.A(_0950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0951_));
 sky130_fd_sc_hd__a21oi_2 _3578_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .A2(_0951_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0952_));
 sky130_fd_sc_hd__a22o_2 _3579_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .A2(_0947_),
    .B1(_0949_),
    .B2(_0952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_1__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_1__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(_0955_),
    .A1(_0954_),
    .S(clknet_1_1__leaf__0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3583_ (.A0(_0956_),
    .A1(_0940_),
    .S(clknet_1_1__leaf__0938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_0__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_0__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(_0958_),
    .A1(_0959_),
    .S(clknet_1_1__leaf__0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _3587_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_0__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_0__leaf__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _3589_ (.A0(_0961_),
    .A1(_0962_),
    .S(clknet_1_0__leaf__0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(_0963_),
    .A1(_0960_),
    .S(clknet_1_0__leaf__0938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _3591_ (.A0(_0957_),
    .A1(_0964_),
    .S(_0953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0965_));
 sky130_fd_sc_hd__nand2_2 _3593_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .B(_0965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux4_2 _3594_ (.A0(net15),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net17),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0966_));
 sky130_fd_sc_hd__and2b_1 _3595_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .B(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0967_));
 sky130_fd_sc_hd__a211o_1 _3596_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .A2(net26),
    .B1(_0133_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0968_));
 sky130_fd_sc_hd__o22a_2 _3597_ (.A1(_0132_),
    .A2(_0966_),
    .B1(_0967_),
    .B2(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _3598_ (.A0(clknet_1_0__leaf_net28),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_2 _3599_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .B(_0970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0971_));
 sky130_fd_sc_hd__mux2_1 _3600_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_2 _3601_ (.A(_0132_),
    .B(_0972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0973_));
 sky130_fd_sc_hd__mux4_1 _3602_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net19),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0974_));
 sky130_fd_sc_hd__nand2_1 _3603_ (.A(_0133_),
    .B(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0975_));
 sky130_fd_sc_hd__o31a_2 _3604_ (.A1(_0133_),
    .A2(_0971_),
    .A3(_0973_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0976_));
 sky130_fd_sc_hd__a2bb2o_2 _3605_ (.A1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .A2_N(_0969_),
    .B1(_0975_),
    .B2(_0976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0977_));
 sky130_fd_sc_hd__mux4_2 _3606_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf_net28),
    .A2(clknet_1_0__leaf_net19),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0978_));
 sky130_fd_sc_hd__and2b_2 _3607_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .B(_0978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0979_));
 sky130_fd_sc_hd__mux4_2 _3608_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0980_));
 sky130_fd_sc_hd__a21bo_2 _3609_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .A2(_0980_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0981_));
 sky130_fd_sc_hd__mux4_2 _3610_ (.A0(net15),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net17),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0982_));
 sky130_fd_sc_hd__and2_2 _3611_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .B(_0982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(net24),
    .A1(net26),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0984_));
 sky130_fd_sc_hd__inv_2 _3613_ (.A(_0984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0985_));
 sky130_fd_sc_hd__a21oi_1 _3614_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .A2(_0985_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0986_));
 sky130_fd_sc_hd__o32a_2 _3615_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .A2(_0983_),
    .A3(_0986_),
    .B1(_0979_),
    .B2(_0981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _3616_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .S(clknet_1_0__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0988_));
 sky130_fd_sc_hd__mux4_2 _3617_ (.A0(net15),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net17),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0989_));
 sky130_fd_sc_hd__and2b_1 _3618_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0990_));
 sky130_fd_sc_hd__a211o_1 _3619_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(net25),
    .B1(_0135_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0991_));
 sky130_fd_sc_hd__o22a_2 _3620_ (.A1(_0134_),
    .A2(_0989_),
    .B1(_0990_),
    .B2(_0991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(clknet_1_0__leaf_net28),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0993_));
 sky130_fd_sc_hd__nor2_2 _3622_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .B(_0993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0994_));
 sky130_fd_sc_hd__mux2_1 _3623_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0995_));
 sky130_fd_sc_hd__nor2_2 _3624_ (.A(_0134_),
    .B(_0995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0996_));
 sky130_fd_sc_hd__mux4_2 _3625_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net19),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0997_));
 sky130_fd_sc_hd__nand2_2 _3626_ (.A(_0135_),
    .B(_0997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0998_));
 sky130_fd_sc_hd__o31a_2 _3627_ (.A1(_0135_),
    .A2(_0994_),
    .A3(_0996_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0999_));
 sky130_fd_sc_hd__a2bb2o_2 _3628_ (.A1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .A2_N(_0992_),
    .B1(_0998_),
    .B2(_0999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .S(clknet_1_0__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _3630_ (.A0(_0988_),
    .A1(_1001_),
    .S(clknet_1_0__leaf__0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1002_));
 sky130_fd_sc_hd__mux4_2 _3631_ (.A0(clknet_1_0__leaf_net28),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1003_));
 sky130_fd_sc_hd__nand2_2 _3632_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .B(_1003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1004_));
 sky130_fd_sc_hd__mux4_2 _3633_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net19),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1005_));
 sky130_fd_sc_hd__nand2b_2 _3634_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .B(_1005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1006_));
 sky130_fd_sc_hd__mux4_2 _3635_ (.A0(net24),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net25),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1007_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf_net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1008_));
 sky130_fd_sc_hd__o211a_1 _3637_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0192_),
    .B1(_1008_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _3638_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .B(_1009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1010_));
 sky130_fd_sc_hd__a211oi_2 _3639_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .A2(_1007_),
    .B1(_1010_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1011_));
 sky130_fd_sc_hd__a31o_2 _3640_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .A2(_1004_),
    .A3(_1006_),
    .B1(_1011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _3641_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .S(clknet_1_1__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _3642_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .S(clknet_1_1__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _3643_ (.A0(_1014_),
    .A1(_1013_),
    .S(clknet_1_1__leaf__0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_1 _3644_ (.A0(_1015_),
    .A1(_1002_),
    .S(clknet_1_1__leaf__1000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .S(clknet_1_1__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _3646_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .S(clknet_1_1__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _3647_ (.A0(_1017_),
    .A1(_1018_),
    .S(clknet_1_1__leaf__0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _3648_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .S(clknet_1_0__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .S(clknet_1_0__leaf__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(_1020_),
    .A1(_1021_),
    .S(clknet_1_0__leaf__0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _3651_ (.A0(_1022_),
    .A1(_1019_),
    .S(clknet_1_0__leaf__1000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(_1016_),
    .A1(_1023_),
    .S(_1012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _3654_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .B(_1024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _3655_ (.A0(clknet_1_0__leaf__0251_),
    .A1(clknet_1_0__leaf__0681_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1025_));
 sky130_fd_sc_hd__a31o_1 _3656_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ),
    .A2(_0080_),
    .A3(clknet_1_0__leaf__0590_),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1026_));
 sky130_fd_sc_hd__a21oi_2 _3657_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ),
    .A2(_1025_),
    .B1(_1026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1027_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(clknet_1_0__leaf__0617_),
    .A1(clknet_1_0__leaf__0723_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1028_));
 sky130_fd_sc_hd__or2_2 _3659_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ),
    .B(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1029_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(clknet_1_0__leaf__0197_),
    .A1(_1030_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1031_));
 sky130_fd_sc_hd__nand2_2 _3662_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ),
    .B(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1032_));
 sky130_fd_sc_hd__a31o_2 _3663_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.D ),
    .A2(_1029_),
    .A3(_1032_),
    .B1(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(clknet_1_1__leaf__1033_),
    .A1(clknet_1_1__leaf_net31),
    .S(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1034_));
 sky130_fd_sc_hd__or2_2 _3665_ (.A(_0084_),
    .B(_1034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1035_));
 sky130_fd_sc_hd__or2_2 _3666_ (.A(_0159_),
    .B(clknet_1_1__leaf__1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf__0565_),
    .S(_0159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_2 _3668_ (.A0(_1036_),
    .A1(_1037_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .A1(clknet_1_1__leaf__0621_),
    .S(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_4 _3670_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.D ),
    .B(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__a21o_2 _3671_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.Q ),
    .A2(net292),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _3672_ (.A0(clknet_1_1__leaf__0251_),
    .A1(clknet_1_0__leaf__0709_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1040_));
 sky130_fd_sc_hd__o21ai_4 _3673_ (.A1(_0152_),
    .A2(_1040_),
    .B1(_1039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ));
 sky130_fd_sc_hd__o21a_1 _3674_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1041_));
 sky130_fd_sc_hd__o21ai_4 _3675_ (.A1(_0147_),
    .A2(clknet_1_1__leaf__0698_),
    .B1(_1041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__nand2_2 _3676_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1042_));
 sky130_fd_sc_hd__o211a_2 _3677_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0688_),
    .B1(_1042_),
    .C1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1043_));
 sky130_fd_sc_hd__nand2b_2 _3678_ (.A_N(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .B(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1044_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .A1(clknet_1_0__leaf__0718_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(_1044_),
    .A1(_1045_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(net424),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1047_));
 sky130_fd_sc_hd__mux4_2 _3682_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .A1(clknet_1_1__leaf__0628_),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .A3(_1047_),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_2 _3683_ (.A0(_1046_),
    .A1(_1048_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1049_));
 sky130_fd_sc_hd__inv_2 _2815__84 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net319));
 sky130_fd_sc_hd__a31o_2 _3685_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ),
    .A2(_0149_),
    .A3(net318),
    .B1(_1043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _3686_ (.A0(clknet_1_0__leaf__0679_),
    .A1(clknet_1_1__leaf__0668_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1052_));
 sky130_fd_sc_hd__mux4_1 _3687_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .A3(_1052_),
    .S0(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_2 _3688_ (.A0(_1051_),
    .A1(_1053_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1054_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .A1(clknet_1_0__leaf__1054_),
    .S(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_2 _3690_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_1_.Q ),
    .B(_1055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_2 _3691_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1056_));
 sky130_fd_sc_hd__o211a_2 _3692_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0688_),
    .B1(_1056_),
    .C1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1057_));
 sky130_fd_sc_hd__a31o_2 _3693_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ),
    .A2(_0157_),
    .A3(net317),
    .B1(_1057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _3694_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1059_));
 sky130_fd_sc_hd__mux4_2 _3695_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .A1(net319),
    .A2(_1059_),
    .A3(net393),
    .S0(_0157_),
    .S1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _3696_ (.A0(_1058_),
    .A1(_1060_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1061_));
 sky130_fd_sc_hd__o21a_2 _3697_ (.A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .A2(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1062_));
 sky130_fd_sc_hd__o21ai_4 _3698_ (.A1(_0158_),
    .A2(clknet_1_0__leaf__1061_),
    .B1(_1062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__and2b_2 _3699_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .B(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1063_));
 sky130_fd_sc_hd__and2_2 _3700_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _3701_ (.A0(clknet_1_0__leaf__0193_),
    .A1(clknet_1_1__leaf__0611_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(_1064_),
    .A1(_1065_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(net26),
    .A1(clknet_1_0__leaf__0650_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1067_));
 sky130_fd_sc_hd__inv_2 _3280__65 (.A(clknet_1_0__leaf__0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net300));
 sky130_fd_sc_hd__nor2_2 _3705_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1069_));
 sky130_fd_sc_hd__a21oi_2 _3706_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0259_),
    .B1(_1069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1070_));
 sky130_fd_sc_hd__mux4_2 _3707_ (.A0(net257),
    .A1(clknet_1_0__leaf__0603_),
    .A2(net299),
    .A3(_1070_),
    .S0(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_2 _3708_ (.A0(_1066_),
    .A1(_1071_),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _3709_ (.A0(net255),
    .A1(clknet_1_1__leaf__1072_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1073_));
 sky130_fd_sc_hd__mux2_1 _3710_ (.A0(_1063_),
    .A1(_1073_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(clknet_1_0__leaf__0227_),
    .A1(clknet_1_1__leaf__0568_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1075_));
 sky130_fd_sc_hd__mux4_2 _3712_ (.A0(net51),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .A3(_1075_),
    .S0(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_2 _3713_ (.A0(_1074_),
    .A1(_1076_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _3714_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .A1(clknet_1_0__leaf__1077_),
    .S(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_2 _3715_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_1_.Q ),
    .B(_1078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__mux2_1 _3716_ (.A0(net261),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1079_));
 sky130_fd_sc_hd__nor2_2 _3717_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_2_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1080_));
 sky130_fd_sc_hd__a22o_2 _3718_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_2_.Q ),
    .A2(_1079_),
    .B1(_1080_),
    .B2(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1081_));
 sky130_fd_sc_hd__a21oi_2 _3719_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0766_),
    .B1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1082_));
 sky130_fd_sc_hd__a31o_2 _3720_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .A2(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .B1(_1082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1083_));
 sky130_fd_sc_hd__a211o_2 _3721_ (.A1(_0114_),
    .A2(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .B1(_1083_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1084_));
 sky130_fd_sc_hd__nor2_1 _3722_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1085_));
 sky130_fd_sc_hd__a211oi_2 _3723_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .A2(clknet_1_0__leaf__0883_),
    .B1(_1085_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1086_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(clknet_1_0__leaf__0704_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_2 _3725_ (.A(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1088_));
 sky130_fd_sc_hd__a211o_2 _3726_ (.A1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0642_),
    .B1(_1088_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1089_));
 sky130_fd_sc_hd__o211a_2 _3727_ (.A1(_0114_),
    .A2(_1087_),
    .B1(_1089_),
    .C1(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1090_));
 sky130_fd_sc_hd__o31a_2 _3728_ (.A1(_0117_),
    .A2(_1086_),
    .A3(_1090_),
    .B1(_1084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1091_));
 sky130_fd_sc_hd__or2_2 _3729_ (.A(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1092_));
 sky130_fd_sc_hd__o21ai_2 _3730_ (.A1(_0119_),
    .A2(clknet_1_1__leaf__1091_),
    .B1(_1092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1093_));
 sky130_fd_sc_hd__mux4_2 _3731_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .A2(clknet_1_1__leaf__0539_),
    .A3(_1093_),
    .S0(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _3732_ (.A0(_1081_),
    .A1(_1094_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(clknet_1_0__leaf__1095_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1096_));
 sky130_fd_sc_hd__nand2_2 _3734_ (.A(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_1_.Q ),
    .B(_1096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__mux4_2 _3735_ (.A0(clknet_1_1__leaf_net49),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net52),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_1 _3736_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .B(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1098_));
 sky130_fd_sc_hd__a211o_1 _3737_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .A2(net20),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .C1(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1099_));
 sky130_fd_sc_hd__o22a_2 _3738_ (.A1(_0101_),
    .A2(_1097_),
    .B1(_1098_),
    .B2(_1099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(clknet_1_0__leaf__0202_),
    .A1(clknet_1_1__leaf__0603_),
    .S(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1101_));
 sky130_fd_sc_hd__and2_2 _3740_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_1_.Q ),
    .B(_1101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1102_));
 sky130_fd_sc_hd__inv_2 _3485__108 (.A(clknet_1_0__leaf__0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net343));
 sky130_fd_sc_hd__mux4_2 _3742_ (.A0(net339),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1104_));
 sky130_fd_sc_hd__mux4_2 _3743_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1105_));
 sky130_fd_sc_hd__a21bo_2 _3744_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .A2(_1105_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1106_));
 sky130_fd_sc_hd__a21o_2 _3745_ (.A1(_0101_),
    .A2(_1104_),
    .B1(_1106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1107_));
 sky130_fd_sc_hd__o21ai_2 _3746_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .A2(_1100_),
    .B1(_1107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1108_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(clknet_1_1__leaf_net49),
    .A1(clknet_1_1__leaf_net52),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1109_));
 sky130_fd_sc_hd__or3_1 _3748_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .B(_0099_),
    .C(_1109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_2 _3749_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net21),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1111_));
 sky130_fd_sc_hd__inv_2 _3824__169 (.A(_1181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net404));
 sky130_fd_sc_hd__a21oi_2 _3751_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .A2(net403),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1113_));
 sky130_fd_sc_hd__mux4_2 _3752_ (.A0(net340),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1114_));
 sky130_fd_sc_hd__mux4_2 _3753_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1115_));
 sky130_fd_sc_hd__or2_2 _3754_ (.A(_0099_),
    .B(_1115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1116_));
 sky130_fd_sc_hd__o211a_2 _3755_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .A2(_1114_),
    .B1(_1116_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1117_));
 sky130_fd_sc_hd__a21oi_2 _3756_ (.A1(_1110_),
    .A2(_1113_),
    .B1(_1117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1118_));
 sky130_fd_sc_hd__mux2_1 _3757_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1119_));
 sky130_fd_sc_hd__mux4_2 _3758_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net20),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1120_));
 sky130_fd_sc_hd__or2_2 _3759_ (.A(_0102_),
    .B(_1120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _3760_ (.A0(clknet_1_1__leaf_net50),
    .A1(clknet_1_1__leaf_net53),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1122_));
 sky130_fd_sc_hd__or3b_1 _3761_ (.A(_1122_),
    .B(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1123_));
 sky130_fd_sc_hd__a21oi_2 _3762_ (.A1(_1121_),
    .A2(_1123_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1124_));
 sky130_fd_sc_hd__or2_1 _3763_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1125_));
 sky130_fd_sc_hd__a21oi_2 _3764_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1126_));
 sky130_fd_sc_hd__mux2_1 _3765_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1127_));
 sky130_fd_sc_hd__inv_2 _4407__193 (.A(_1726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net428));
 sky130_fd_sc_hd__a221o_2 _3767_ (.A1(_1125_),
    .A2(_1126_),
    .B1(net427),
    .B2(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_1 _3768_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _3769_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1131_));
 sky130_fd_sc_hd__o21a_2 _3770_ (.A1(_0102_),
    .A2(_1131_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1132_));
 sky130_fd_sc_hd__o21ai_2 _3771_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .A2(_1130_),
    .B1(_1132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1133_));
 sky130_fd_sc_hd__a31o_2 _3772_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .A2(_1129_),
    .A3(_1133_),
    .B1(_1124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _3774_ (.A0(_1119_),
    .A1(_1135_),
    .S(clknet_1_0__leaf__1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1136_));
 sky130_fd_sc_hd__nand2b_2 _3775_ (.A_N(_1136_),
    .B(clknet_1_0__leaf__1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1137_));
 sky130_fd_sc_hd__mux2_1 _3776_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_1__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(_1138_),
    .A1(_1139_),
    .S(clknet_1_0__leaf__1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1140_));
 sky130_fd_sc_hd__mux4_2 _3779_ (.A0(clknet_1_1__leaf_net49),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net52),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1141_));
 sky130_fd_sc_hd__nor2_1 _3780_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1142_));
 sky130_fd_sc_hd__a211o_1 _3781_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .A2(net21),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .C1(_0103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1143_));
 sky130_fd_sc_hd__o22a_2 _3782_ (.A1(_0104_),
    .A2(_1141_),
    .B1(_1142_),
    .B2(_1143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1144_));
 sky130_fd_sc_hd__mux4_1 _3783_ (.A0(net341),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1145_));
 sky130_fd_sc_hd__mux4_2 _3784_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1146_));
 sky130_fd_sc_hd__a21bo_2 _3785_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .A2(_1146_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1147_));
 sky130_fd_sc_hd__a21o_1 _3786_ (.A1(_0104_),
    .A2(_1145_),
    .B1(_1147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1148_));
 sky130_fd_sc_hd__o21ai_1 _3787_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .A2(_1144_),
    .B1(_1148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1149_));
 sky130_fd_sc_hd__o21ba_1 _3788_ (.A1(clknet_1_0__leaf__1134_),
    .A2(_1140_),
    .B1_N(clknet_1_0__leaf__1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _3789_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(_1151_),
    .A1(_1152_),
    .S(clknet_1_1__leaf__1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _3792_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_0__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _3794_ (.A0(_1155_),
    .A1(_1154_),
    .S(clknet_1_1__leaf__1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1156_));
 sky130_fd_sc_hd__mux2_1 _3795_ (.A0(_1156_),
    .A1(_1153_),
    .S(clknet_1_1__leaf__1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1157_));
 sky130_fd_sc_hd__a22o_1 _3796_ (.A1(_1137_),
    .A2(_1150_),
    .B1(_1157_),
    .B2(clknet_1_1__leaf__1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3797_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1158_));
 sky130_fd_sc_hd__nand2_4 _3798_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .B(_1158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _3799_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .A1(clknet_1_1__leaf__0730_),
    .S(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1159_));
 sky130_fd_sc_hd__nand2_2 _3800_ (.A(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_1_.Q ),
    .B(_1159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__mux2_1 _3801_ (.A0(clknet_1_0__leaf__0846_),
    .A1(clknet_1_1__leaf__0193_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1160_));
 sky130_fd_sc_hd__and2b_2 _3802_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .B(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_2 _3803_ (.A0(_1160_),
    .A1(_1161_),
    .S(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1162_));
 sky130_fd_sc_hd__nor2_2 _3804_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ),
    .B(clknet_1_0__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1163_));
 sky130_fd_sc_hd__a21o_2 _3805_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0550_),
    .B1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _3806_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _3807_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .A1(_1165_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1166_));
 sky130_fd_sc_hd__o221a_2 _3808_ (.A1(_1163_),
    .A2(_1164_),
    .B1(_1166_),
    .B2(_0141_),
    .C1(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1167_));
 sky130_fd_sc_hd__a21oi_4 _3809_ (.A1(_1162_),
    .A2(_0142_),
    .B1(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1168_));
 sky130_fd_sc_hd__o21ai_2 _3810_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .A2(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_0_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1169_));
 sky130_fd_sc_hd__a21o_2 _3811_ (.A1(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__1168_),
    .B1(_1169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__mux4_2 _3812_ (.A0(clknet_1_1__leaf_net49),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net52),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1170_));
 sky130_fd_sc_hd__nor2_1 _3813_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1171_));
 sky130_fd_sc_hd__a211o_1 _3814_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .A2(net21),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .C1(_0093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1172_));
 sky130_fd_sc_hd__o22a_2 _3815_ (.A1(_0094_),
    .A2(_1170_),
    .B1(_1171_),
    .B2(_1172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1173_));
 sky130_fd_sc_hd__mux4_2 _3816_ (.A0(net342),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1174_));
 sky130_fd_sc_hd__mux4_2 _3817_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1175_));
 sky130_fd_sc_hd__a21bo_2 _3818_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .A2(_1175_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1176_));
 sky130_fd_sc_hd__a21o_2 _3819_ (.A1(_0094_),
    .A2(_1174_),
    .B1(_1176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1177_));
 sky130_fd_sc_hd__o21ai_2 _3820_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .A2(_1173_),
    .B1(_1177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1178_));
 sky130_fd_sc_hd__mux2_1 _3821_ (.A0(clknet_1_0__leaf_net49),
    .A1(clknet_1_0__leaf_net52),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1179_));
 sky130_fd_sc_hd__or3_1 _3822_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .B(_0092_),
    .C(_1179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1180_));
 sky130_fd_sc_hd__mux4_2 _3823_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net20),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1181_));
 sky130_fd_sc_hd__inv_2 _4224__170 (.A(_1556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net405));
 sky130_fd_sc_hd__a21oi_2 _3825_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .A2(net404),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1183_));
 sky130_fd_sc_hd__mux4_2 _3826_ (.A0(clknet_1_1__leaf_net22),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1184_));
 sky130_fd_sc_hd__mux4_2 _3827_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1185_));
 sky130_fd_sc_hd__or2_2 _3828_ (.A(_0092_),
    .B(_1185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1186_));
 sky130_fd_sc_hd__o211a_2 _3829_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .A2(_1184_),
    .B1(_1186_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1187_));
 sky130_fd_sc_hd__a21oi_2 _3830_ (.A1(_1180_),
    .A2(_1183_),
    .B1(_1187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1188_));
 sky130_fd_sc_hd__mux2_1 _3831_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1189_));
 sky130_fd_sc_hd__mux4_2 _3832_ (.A0(clknet_1_1__leaf_net49),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net52),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1190_));
 sky130_fd_sc_hd__nor2_1 _3833_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1191_));
 sky130_fd_sc_hd__a211o_1 _3834_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .A2(net21),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .C1(_0095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1192_));
 sky130_fd_sc_hd__o22a_2 _3835_ (.A1(_0096_),
    .A2(_1190_),
    .B1(_1191_),
    .B2(_1192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1193_));
 sky130_fd_sc_hd__nor2_2 _3836_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .B(_1193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1194_));
 sky130_fd_sc_hd__mux4_2 _3837_ (.A0(clknet_1_1__leaf_net22),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1195_));
 sky130_fd_sc_hd__nand2_2 _3838_ (.A(_0096_),
    .B(_1195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1196_));
 sky130_fd_sc_hd__mux4_2 _3839_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1197_));
 sky130_fd_sc_hd__nand2_2 _3840_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .B(_1197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1198_));
 sky130_fd_sc_hd__a31o_2 _3841_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .A2(_1196_),
    .A3(_1198_),
    .B1(_1194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _3842_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _3843_ (.A0(_1189_),
    .A1(_1200_),
    .S(clknet_1_1__leaf__1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1201_));
 sky130_fd_sc_hd__nand2b_2 _3844_ (.A_N(_1201_),
    .B(clknet_1_0__leaf__1199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1202_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1203_));
 sky130_fd_sc_hd__mux2_1 _3846_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_1__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(_1203_),
    .A1(_1204_),
    .S(clknet_1_1__leaf__1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1205_));
 sky130_fd_sc_hd__mux4_2 _3848_ (.A0(clknet_1_1__leaf_net49),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net52),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1206_));
 sky130_fd_sc_hd__nor2_1 _3849_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1207_));
 sky130_fd_sc_hd__a211o_1 _3850_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .A2(net21),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .C1(_0097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1208_));
 sky130_fd_sc_hd__o22a_1 _3851_ (.A1(_0098_),
    .A2(_1206_),
    .B1(_1207_),
    .B2(_1208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1209_));
 sky130_fd_sc_hd__mux4_2 _3852_ (.A0(clknet_1_1__leaf_net22),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1210_));
 sky130_fd_sc_hd__mux4_2 _3853_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1211_));
 sky130_fd_sc_hd__a21bo_2 _3854_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .A2(_1211_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1212_));
 sky130_fd_sc_hd__a21o_2 _3855_ (.A1(_0098_),
    .A2(_1210_),
    .B1(_1212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1213_));
 sky130_fd_sc_hd__o21ai_1 _3856_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .A2(_1209_),
    .B1(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1214_));
 sky130_fd_sc_hd__o21ba_1 _3857_ (.A1(clknet_1_1__leaf__1199_),
    .A2(_1205_),
    .B1_N(clknet_1_1__leaf__1214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _3859_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1217_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(_1216_),
    .A1(_1217_),
    .S(clknet_1_0__leaf__1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_0__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1220_));
 sky130_fd_sc_hd__mux2_1 _3863_ (.A0(_1220_),
    .A1(_1219_),
    .S(clknet_1_0__leaf__1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _3864_ (.A0(_1221_),
    .A1(_1218_),
    .S(clknet_1_0__leaf__1199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1222_));
 sky130_fd_sc_hd__a22o_1 _3865_ (.A1(_1202_),
    .A2(_1215_),
    .B1(_1222_),
    .B2(clknet_1_0__leaf__1214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3866_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1223_));
 sky130_fd_sc_hd__nand2_4 _3867_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .B(_1223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__a21o_1 _3868_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_1_.Q ),
    .A2(clknet_1_1__leaf__0547_),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(clknet_1_1__leaf__0528_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1225_));
 sky130_fd_sc_hd__o21ai_2 _3870_ (.A1(_0118_),
    .A2(_1225_),
    .B1(_1224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1226_));
 sky130_fd_sc_hd__mux2_1 _3871_ (.A0(clknet_1_1__leaf__0558_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1227_));
 sky130_fd_sc_hd__inv_2 _2809__145 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net380));
 sky130_fd_sc_hd__mux4_2 _3873_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .A1(clknet_1_1__leaf__0655_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .A3(net379),
    .S0(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1229_));
 sky130_fd_sc_hd__inv_2 _2814__158 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net393));
 sky130_fd_sc_hd__mux2_1 _3875_ (.A0(_1226_),
    .A1(net392),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1231_));
 sky130_fd_sc_hd__o21ai_2 _3876_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .A2(_0160_),
    .B1(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1232_));
 sky130_fd_sc_hd__a21o_2 _3877_ (.A1(_0160_),
    .A2(clknet_1_0__leaf__1231_),
    .B1(_1232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .A1(clknet_1_1__leaf__0192_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1233_));
 sky130_fd_sc_hd__mux4_1 _3879_ (.A0(clknet_1_1__leaf__0232_),
    .A1(net368),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .A3(_1233_),
    .S0(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _3880_ (.A0(net254),
    .A1(clknet_1_0__leaf__1072_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1235_));
 sky130_fd_sc_hd__or3b_2 _3881_ (.A(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_2_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .C_N(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1236_));
 sky130_fd_sc_hd__a21bo_2 _3882_ (.A1(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_2_.Q ),
    .A2(_1235_),
    .B1_N(_1236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1237_));
 sky130_fd_sc_hd__mux2_2 _3883_ (.A0(_1237_),
    .A1(_1234_),
    .S(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _3884_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .A1(clknet_1_0__leaf__1238_),
    .S(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1239_));
 sky130_fd_sc_hd__nand2_2 _3885_ (.A(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_1_.Q ),
    .B(_1239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__a21oi_1 _3886_ (.A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .A2(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ),
    .B1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1240_));
 sky130_fd_sc_hd__nor2_2 _3887_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1241_));
 sky130_fd_sc_hd__a311o_2 _3888_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ),
    .A2(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_2_.Q ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .B1(_1240_),
    .C1(_1241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _3889_ (.A0(clknet_1_1__leaf__0259_),
    .A1(clknet_1_0__leaf__1091_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1243_));
 sky130_fd_sc_hd__mux4_2 _3890_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .A2(net423),
    .A3(_1243_),
    .S0(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _3891_ (.A0(_1242_),
    .A1(_1244_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__nor2_2 _3892_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1245_));
 sky130_fd_sc_hd__a211o_2 _3893_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1245_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1247_));
 sky130_fd_sc_hd__inv_2 _3918__81 (.A(_1270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net316));
 sky130_fd_sc_hd__a21oi_2 _3896_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .A2(net315),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1249_));
 sky130_fd_sc_hd__mux4_2 _3897_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_0__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1250_));
 sky130_fd_sc_hd__a22o_2 _3898_ (.A1(_1246_),
    .A2(_1249_),
    .B1(_1250_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1251_));
 sky130_fd_sc_hd__mux4_2 _3899_ (.A0(clknet_1_0__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1252_));
 sky130_fd_sc_hd__o21ai_2 _3900_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0197_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1253_));
 sky130_fd_sc_hd__a21o_2 _3901_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(net36),
    .B1(_1253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_1 _3902_ (.A0(_1254_),
    .A1(_1252_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(_1255_),
    .A1(_1251_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1256_));
 sky130_fd_sc_hd__mux4_2 _3904_ (.A0(clknet_1_0__leaf__0901_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1257_));
 sky130_fd_sc_hd__mux4_2 _3905_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_0__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1258_));
 sky130_fd_sc_hd__or2_2 _3906_ (.A(_0070_),
    .B(_1258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1259_));
 sky130_fd_sc_hd__o211a_2 _3907_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .A2(_1257_),
    .B1(_1259_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1261_));
 sky130_fd_sc_hd__or3_2 _3909_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .B(_0070_),
    .C(_1261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1262_));
 sky130_fd_sc_hd__mux4_2 _3910_ (.A0(clknet_1_0__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1263_));
 sky130_fd_sc_hd__inv_2 _3925__126 (.A(_1277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net361));
 sky130_fd_sc_hd__a21oi_2 _3912_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .A2(net360),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1265_));
 sky130_fd_sc_hd__a21oi_2 _3913_ (.A1(_1262_),
    .A2(_1265_),
    .B1(_1260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1266_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_1__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1267_));
 sky130_fd_sc_hd__nor2_2 _3915_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1268_));
 sky130_fd_sc_hd__a211o_2 _3916_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1268_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1270_));
 sky130_fd_sc_hd__inv_2 _3684__82 (.A(clknet_1_0__leaf__1049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net317));
 sky130_fd_sc_hd__a21oi_2 _3919_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .A2(net316),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1272_));
 sky130_fd_sc_hd__mux4_2 _3920_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_0__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1273_));
 sky130_fd_sc_hd__a22o_2 _3921_ (.A1(_1269_),
    .A2(_1272_),
    .B1(_1273_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1274_));
 sky130_fd_sc_hd__o21ai_2 _3922_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0197_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1275_));
 sky130_fd_sc_hd__a211o_2 _3923_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(net36),
    .B1(_1275_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1276_));
 sky130_fd_sc_hd__mux4_2 _3924_ (.A0(clknet_1_0__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1277_));
 sky130_fd_sc_hd__inv_2 _3995__127 (.A(_1343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net362));
 sky130_fd_sc_hd__a21oi_2 _3926_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .A2(net361),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1279_));
 sky130_fd_sc_hd__a22o_2 _3927_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .A2(_1274_),
    .B1(_1276_),
    .B2(_1279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1280_));
 sky130_fd_sc_hd__mux2_1 _3928_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_1__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(_1267_),
    .A1(_1281_),
    .S(clknet_1_1__leaf__1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1282_));
 sky130_fd_sc_hd__nor2_2 _3930_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1283_));
 sky130_fd_sc_hd__a211o_2 _3931_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1283_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1285_));
 sky130_fd_sc_hd__o21ba_2 _3933_ (.A1(_0071_),
    .A2(_1285_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1286_));
 sky130_fd_sc_hd__mux4_2 _3934_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_0__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1287_));
 sky130_fd_sc_hd__a22o_2 _3935_ (.A1(_1284_),
    .A2(_1286_),
    .B1(_1287_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1288_));
 sky130_fd_sc_hd__mux4_2 _3936_ (.A0(clknet_1_0__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1290_));
 sky130_fd_sc_hd__or3b_2 _3938_ (.A(_1290_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1291_));
 sky130_fd_sc_hd__o21a_2 _3939_ (.A1(_0071_),
    .A2(_1289_),
    .B1(_1291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _3940_ (.A0(_1292_),
    .A1(_1288_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _3941_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_1__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _3942_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _3943_ (.A0(_1294_),
    .A1(_1295_),
    .S(clknet_1_1__leaf__1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1296_));
 sky130_fd_sc_hd__mux2_1 _3944_ (.A0(_1282_),
    .A1(_1296_),
    .S(clknet_1_1__leaf__1280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_1 _3945_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_0__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1298_));
 sky130_fd_sc_hd__mux2_1 _3946_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1299_));
 sky130_fd_sc_hd__mux2_1 _3947_ (.A0(_1298_),
    .A1(_1299_),
    .S(clknet_1_0__leaf__1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _3948_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_0__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1301_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_0__leaf__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_1 _3950_ (.A0(_1301_),
    .A1(_1302_),
    .S(clknet_1_0__leaf__1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _3951_ (.A0(_1303_),
    .A1(_1300_),
    .S(clknet_1_0__leaf__1280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(_1297_),
    .A1(_1304_),
    .S(_1293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _3953_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1305_));
 sky130_fd_sc_hd__nand2_1 _3954_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .B(_1305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(clknet_1_0__leaf__0221_),
    .A1(clknet_1_0__leaf__0624_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1306_));
 sky130_fd_sc_hd__and3b_2 _3956_ (.A_N(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ),
    .B(clknet_1_0__leaf__0561_),
    .C(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1307_));
 sky130_fd_sc_hd__a21o_2 _3957_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ),
    .A2(_1306_),
    .B1(_1307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _3959_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .A1(_1309_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1310_));
 sky130_fd_sc_hd__nand2b_2 _3960_ (.A_N(_1310_),
    .B(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1311_));
 sky130_fd_sc_hd__or3b_2 _3961_ (.A(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ),
    .B(net364),
    .C_N(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1312_));
 sky130_fd_sc_hd__o311a_2 _3962_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ),
    .A2(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ),
    .A3(_0686_),
    .B1(_1311_),
    .C1(_1312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _3963_ (.A0(_1308_),
    .A1(_1313_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1314_));
 sky130_fd_sc_hd__nand2b_1 _3964_ (.A_N(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1315_));
 sky130_fd_sc_hd__o211a_1 _3965_ (.A1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__1314_),
    .B1(_1315_),
    .C1(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1316_));
 sky130_fd_sc_hd__nand2_1 _3966_ (.A(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.Q ),
    .B(clknet_1_1__leaf__1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1317_));
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(net301),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_4 _3968_ (.A0(_1317_),
    .A1(_1318_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__mux2_1 _3969_ (.A0(clknet_1_1__leaf__0704_),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1319_));
 sky130_fd_sc_hd__mux4_1 _3970_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .A2(net343),
    .A3(_1319_),
    .S0(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_1 _3971_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1321_));
 sky130_fd_sc_hd__and3b_1 _3972_ (.A_N(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_2_.Q ),
    .B(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_1_.Q ),
    .C(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1322_));
 sky130_fd_sc_hd__a21oi_2 _3973_ (.A1(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_2_.Q ),
    .A2(_1321_),
    .B1(_1322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1323_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(_1323_),
    .A1(_1320_),
    .S(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__nor2_2 _3975_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1324_));
 sky130_fd_sc_hd__a211o_2 _3976_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1324_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1326_));
 sky130_fd_sc_hd__inv_2 _4002__75 (.A(_1350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net310));
 sky130_fd_sc_hd__a21oi_2 _3979_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .A2(net309),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1328_));
 sky130_fd_sc_hd__mux4_1 _3980_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_1__leaf_net33),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1329_));
 sky130_fd_sc_hd__a22o_1 _3981_ (.A1(_1325_),
    .A2(_1328_),
    .B1(_1329_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1330_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net37),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1331_));
 sky130_fd_sc_hd__or3b_2 _3983_ (.A(_1331_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1332_));
 sky130_fd_sc_hd__mux4_2 _3984_ (.A0(clknet_1_1__leaf_net29),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1333_));
 sky130_fd_sc_hd__inv_2 _4023__120 (.A(_1371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net355));
 sky130_fd_sc_hd__a21oi_2 _3986_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .A2(net354),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1335_));
 sky130_fd_sc_hd__a22o_1 _3987_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .A2(_1330_),
    .B1(_1332_),
    .B2(_1335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1336_));
 sky130_fd_sc_hd__mux4_2 _3988_ (.A0(clknet_1_1__leaf__0901_),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1337_));
 sky130_fd_sc_hd__mux4_2 _3989_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(clknet_1_1__leaf_net33),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1338_));
 sky130_fd_sc_hd__or2_2 _3990_ (.A(_0073_),
    .B(_1338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1339_));
 sky130_fd_sc_hd__o211a_2 _3991_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .A2(_1337_),
    .B1(_1339_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1340_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net36),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1341_));
 sky130_fd_sc_hd__or3_2 _3993_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .B(_0073_),
    .C(_1341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1342_));
 sky130_fd_sc_hd__mux4_2 _3994_ (.A0(clknet_1_1__leaf_net29),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net31),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1343_));
 sky130_fd_sc_hd__inv_2 _2803__128 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net363));
 sky130_fd_sc_hd__a21oi_2 _3996_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .A2(net362),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1345_));
 sky130_fd_sc_hd__a21oi_2 _3997_ (.A1(_1342_),
    .A2(_1345_),
    .B1(_1340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1346_));
 sky130_fd_sc_hd__mux2_1 _3998_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_0__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1347_));
 sky130_fd_sc_hd__nor2_2 _3999_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1348_));
 sky130_fd_sc_hd__a211o_2 _4000_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1348_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_1 _4001_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1350_));
 sky130_fd_sc_hd__inv_2 _4016__76 (.A(_1364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net311));
 sky130_fd_sc_hd__a21oi_2 _4003_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .A2(net310),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1352_));
 sky130_fd_sc_hd__mux4_2 _4004_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(net34),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1353_));
 sky130_fd_sc_hd__a22o_2 _4005_ (.A1(_1349_),
    .A2(_1352_),
    .B1(_1353_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1354_));
 sky130_fd_sc_hd__mux4_2 _4006_ (.A0(net30),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1355_));
 sky130_fd_sc_hd__o21ai_2 _4007_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0197_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1356_));
 sky130_fd_sc_hd__a21o_2 _4008_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .A2(net36),
    .B1(_1356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1357_));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(_1357_),
    .A1(_1355_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_1 _4010_ (.A0(_1358_),
    .A1(_1354_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _4012_ (.A0(_1347_),
    .A1(_1360_),
    .S(clknet_1_0__leaf__1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1361_));
 sky130_fd_sc_hd__nor2_2 _4013_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1362_));
 sky130_fd_sc_hd__a211o_2 _4014_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1362_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1364_));
 sky130_fd_sc_hd__inv_2 _3531__77 (.A(_0904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net312));
 sky130_fd_sc_hd__a21oi_2 _4017_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .A2(net311),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1366_));
 sky130_fd_sc_hd__mux4_2 _4018_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(net34),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1367_));
 sky130_fd_sc_hd__a22o_2 _4019_ (.A1(_1363_),
    .A2(_1366_),
    .B1(_1367_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_1 _4020_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net37),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1369_));
 sky130_fd_sc_hd__or3b_2 _4021_ (.A(_1369_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1370_));
 sky130_fd_sc_hd__mux4_2 _4022_ (.A0(net30),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1371_));
 sky130_fd_sc_hd__inv_2 _4136__121 (.A(_1479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net356));
 sky130_fd_sc_hd__a21oi_2 _4024_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .A2(net355),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1373_));
 sky130_fd_sc_hd__a22o_2 _4025_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .A2(_1368_),
    .B1(_1370_),
    .B2(_1373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1375_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(_1376_),
    .A1(_1375_),
    .S(clknet_1_0__leaf__1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(_1377_),
    .A1(_1361_),
    .S(clknet_1_0__leaf__1359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_1__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(_1379_),
    .A1(_1380_),
    .S(clknet_1_1__leaf__1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _4034_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(_1382_),
    .A1(_1383_),
    .S(clknet_1_1__leaf__1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(_1384_),
    .A1(_1381_),
    .S(clknet_1_1__leaf__1359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(_1378_),
    .A1(_1385_),
    .S(_1374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _4039_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .B(_1386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__a21o_1 _4040_ (.A1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.Q ),
    .A2(net280),
    .B1(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1387_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(net302),
    .A1(net410),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1388_));
 sky130_fd_sc_hd__mux4_2 _4042_ (.A0(net256),
    .A1(clknet_1_0__leaf__0889_),
    .A2(clknet_1_0__leaf_net35),
    .A3(_1388_),
    .S0(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1389_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1390_));
 sky130_fd_sc_hd__and3b_1 _4044_ (.A_N(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_1_.Q ),
    .B(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_2_.Q ),
    .C(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1391_));
 sky130_fd_sc_hd__a21o_1 _4045_ (.A1(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_1_.Q ),
    .A2(_1390_),
    .B1(_1391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _4046_ (.A0(_1392_),
    .A1(_1389_),
    .S(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1393_));
 sky130_fd_sc_hd__or2_2 _4047_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .B(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1394_));
 sky130_fd_sc_hd__o211a_2 _4048_ (.A1(_0154_),
    .A2(clknet_1_1__leaf__1393_),
    .B1(_1394_),
    .C1(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_2 _4049_ (.A0(clknet_1_1__leaf__1395_),
    .A1(clknet_1_0__leaf__0525_),
    .S(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1396_));
 sky130_fd_sc_hd__o21ai_4 _4050_ (.A1(_1396_),
    .A2(_0155_),
    .B1(_1387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_1 _4052_ (.A0(net15),
    .A1(clknet_1_1__leaf_net16),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1398_));
 sky130_fd_sc_hd__o21a_1 _4053_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .A2(_1398_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1399_));
 sky130_fd_sc_hd__o21ai_2 _4054_ (.A1(_0129_),
    .A2(_1397_),
    .B1(_1399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1400_));
 sky130_fd_sc_hd__mux2_1 _4055_ (.A0(clknet_1_0__leaf_net23),
    .A1(net26),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1401_));
 sky130_fd_sc_hd__nor2_1 _4056_ (.A(_0129_),
    .B(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1402_));
 sky130_fd_sc_hd__o21ba_1 _4057_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .A2(_1402_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1403_));
 sky130_fd_sc_hd__mux4_2 _4058_ (.A0(clknet_1_1__leaf_net28),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1404_));
 sky130_fd_sc_hd__nand2_2 _4059_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .B(_1404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1405_));
 sky130_fd_sc_hd__mux4_2 _4060_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_2 _4061_ (.A(_0129_),
    .B(_1406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1407_));
 sky130_fd_sc_hd__a32o_2 _4062_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .A2(_1405_),
    .A3(_1407_),
    .B1(_1400_),
    .B2(_1403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1408_));
 sky130_fd_sc_hd__mux4_2 _4063_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf_net27),
    .A2(clknet_1_1__leaf_net19),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_2 _4064_ (.A(_0127_),
    .B(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1410_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1411_));
 sky130_fd_sc_hd__nor2_2 _4066_ (.A(_0128_),
    .B(_1411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1413_));
 sky130_fd_sc_hd__nor2_2 _4068_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .B(_1413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1414_));
 sky130_fd_sc_hd__o311a_2 _4069_ (.A1(_0127_),
    .A2(_1412_),
    .A3(_1414_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .C1(_1410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1415_));
 sky130_fd_sc_hd__mux4_2 _4070_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net16),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1416_));
 sky130_fd_sc_hd__and2b_1 _4071_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf_net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1417_));
 sky130_fd_sc_hd__a211o_1 _4072_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .A2(net26),
    .B1(_0128_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1418_));
 sky130_fd_sc_hd__o22a_2 _4073_ (.A1(_0127_),
    .A2(_1416_),
    .B1(_1417_),
    .B2(_1418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1419_));
 sky130_fd_sc_hd__o21ba_2 _4074_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .A2(_1419_),
    .B1_N(_1415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1420_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .S(clknet_1_0__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1421_));
 sky130_fd_sc_hd__mux4_2 _4076_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf_net27),
    .A2(clknet_1_0__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1422_));
 sky130_fd_sc_hd__nand2_2 _4077_ (.A(_0130_),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1423_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1424_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1425_));
 sky130_fd_sc_hd__o21a_2 _4080_ (.A1(_0131_),
    .A2(_1425_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1426_));
 sky130_fd_sc_hd__o21ai_2 _4081_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .A2(_1424_),
    .B1(_1426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1427_));
 sky130_fd_sc_hd__mux2_1 _4082_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1428_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(clknet_1_0__leaf_net23),
    .A1(net25),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1429_));
 sky130_fd_sc_hd__o21a_1 _4084_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .A2(_1429_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1430_));
 sky130_fd_sc_hd__o21ai_1 _4085_ (.A1(_0130_),
    .A2(_1428_),
    .B1(_1430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1431_));
 sky130_fd_sc_hd__nand2_1 _4086_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1432_));
 sky130_fd_sc_hd__o211a_1 _4087_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0192_),
    .B1(_1432_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1433_));
 sky130_fd_sc_hd__o21ba_1 _4088_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .A2(_1433_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1434_));
 sky130_fd_sc_hd__a32o_1 _4089_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .A2(_1423_),
    .A3(_1427_),
    .B1(_1431_),
    .B2(_1434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .S(clknet_1_0__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(_1421_),
    .A1(_1436_),
    .S(clknet_1_1__leaf__1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1437_));
 sky130_fd_sc_hd__mux4_2 _4092_ (.A0(clknet_1_0__leaf_net23),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net25),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_1 _4093_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf_net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1439_));
 sky130_fd_sc_hd__o211a_1 _4094_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0192_),
    .B1(_1439_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1440_));
 sky130_fd_sc_hd__nor2_1 _4095_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .B(_1440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1441_));
 sky130_fd_sc_hd__a211oi_2 _4096_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .A2(_1438_),
    .B1(_1441_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1442_));
 sky130_fd_sc_hd__mux4_2 _4097_ (.A0(clknet_1_0__leaf_net27),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1443_));
 sky130_fd_sc_hd__nand2_2 _4098_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .B(_1443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1444_));
 sky130_fd_sc_hd__mux4_2 _4099_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net18),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1445_));
 sky130_fd_sc_hd__nand2b_2 _4100_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .B(_1445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1446_));
 sky130_fd_sc_hd__a31o_2 _4101_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .A2(_1444_),
    .A3(_1446_),
    .B1(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1447_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .S(clknet_1_0__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _4103_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .S(clknet_1_0__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _4104_ (.A0(_1449_),
    .A1(_1448_),
    .S(clknet_1_0__leaf__1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1450_));
 sky130_fd_sc_hd__mux2_1 _4105_ (.A0(_1450_),
    .A1(_1437_),
    .S(clknet_1_0__leaf__1435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .S(clknet_1_1__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .S(clknet_1_1__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(_1452_),
    .A1(_1453_),
    .S(clknet_1_0__leaf__1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .S(clknet_1_1__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1455_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .S(clknet_1_1__leaf__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(_1455_),
    .A1(_1456_),
    .S(clknet_1_1__leaf__1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_1 _4112_ (.A0(_1457_),
    .A1(_1454_),
    .S(clknet_1_1__leaf__1435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(_1451_),
    .A1(_1458_),
    .S(_1447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1459_));
 sky130_fd_sc_hd__nand2_4 _4115_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .B(_1459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__nor2_2 _4116_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1460_));
 sky130_fd_sc_hd__a211o_2 _4117_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1460_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _4118_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1462_));
 sky130_fd_sc_hd__o21ba_2 _4119_ (.A1(_0075_),
    .A2(_1462_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1463_));
 sky130_fd_sc_hd__mux4_2 _4120_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(net34),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1464_));
 sky130_fd_sc_hd__a22o_2 _4121_ (.A1(_1461_),
    .A2(_1463_),
    .B1(_1464_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1465_));
 sky130_fd_sc_hd__mux4_2 _4122_ (.A0(net30),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net37),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1467_));
 sky130_fd_sc_hd__or3b_2 _4124_ (.A(_1467_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1468_));
 sky130_fd_sc_hd__o21a_2 _4125_ (.A1(_0075_),
    .A2(_1466_),
    .B1(_1468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(_1469_),
    .A1(_1465_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1470_));
 sky130_fd_sc_hd__or2_2 _4127_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1471_));
 sky130_fd_sc_hd__a21oi_2 _4128_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .A2(net421),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _4129_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1473_));
 sky130_fd_sc_hd__a221o_2 _4130_ (.A1(_1471_),
    .A2(_1472_),
    .B1(_1473_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1474_));
 sky130_fd_sc_hd__mux4_2 _4131_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(net34),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1475_));
 sky130_fd_sc_hd__or2_2 _4132_ (.A(_0074_),
    .B(_1475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1476_));
 sky130_fd_sc_hd__o21ai_2 _4133_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0197_),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1477_));
 sky130_fd_sc_hd__a211o_2 _4134_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .A2(net37),
    .B1(_1477_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1478_));
 sky130_fd_sc_hd__mux4_2 _4135_ (.A0(net30),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1479_));
 sky130_fd_sc_hd__inv_2 _3538__122 (.A(_0911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net357));
 sky130_fd_sc_hd__a21oi_2 _4137_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .A2(net356),
    .B1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1481_));
 sky130_fd_sc_hd__a32o_2 _4138_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .A2(_1474_),
    .A3(_1476_),
    .B1(_1478_),
    .B2(_1481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .S(clknet_1_0__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1483_));
 sky130_fd_sc_hd__nor2_2 _4140_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1484_));
 sky130_fd_sc_hd__a211o_2 _4141_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1484_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _4142_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1486_));
 sky130_fd_sc_hd__o21ba_2 _4143_ (.A1(_0076_),
    .A2(_1486_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1487_));
 sky130_fd_sc_hd__mux4_2 _4144_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(net34),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1488_));
 sky130_fd_sc_hd__a22o_2 _4145_ (.A1(_1485_),
    .A2(_1487_),
    .B1(_1488_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1489_));
 sky130_fd_sc_hd__mux4_1 _4146_ (.A0(net30),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4147_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net37),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1491_));
 sky130_fd_sc_hd__or3b_2 _4148_ (.A(_1491_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1492_));
 sky130_fd_sc_hd__o21a_1 _4149_ (.A1(_0076_),
    .A2(_1490_),
    .B1(_1492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(_1493_),
    .A1(_1489_),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _4151_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .S(clknet_1_0__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(_1483_),
    .A1(_1495_),
    .S(clknet_1_0__leaf__1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1496_));
 sky130_fd_sc_hd__nor2_2 _4153_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1497_));
 sky130_fd_sc_hd__a211o_2 _4154_ (.A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(_1497_),
    .C1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _4155_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1499_));
 sky130_fd_sc_hd__o21ba_2 _4156_ (.A1(_0077_),
    .A2(_1499_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1500_));
 sky130_fd_sc_hd__mux4_2 _4157_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(net34),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1501_));
 sky130_fd_sc_hd__a22o_2 _4158_ (.A1(_1498_),
    .A2(_1500_),
    .B1(_1501_),
    .B2(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1502_));
 sky130_fd_sc_hd__mux4_2 _4159_ (.A0(net30),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net32),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _4160_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(net37),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1504_));
 sky130_fd_sc_hd__or3b_2 _4161_ (.A(_1504_),
    .B(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1505_));
 sky130_fd_sc_hd__o21a_2 _4162_ (.A1(_0077_),
    .A2(_1503_),
    .B1(_1505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _4163_ (.A0(_1506_),
    .A1(_1502_),
    .S(\dut_0.U0_formal_verification.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .S(clknet_1_0__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_1 _4165_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .S(clknet_1_0__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(_1509_),
    .A1(_1508_),
    .S(clknet_1_0__leaf__1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(_1510_),
    .A1(_1496_),
    .S(clknet_1_0__leaf__1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _4168_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .S(clknet_1_1__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .S(clknet_1_1__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(_1512_),
    .A1(_1513_),
    .S(clknet_1_1__leaf__1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .S(clknet_1_1__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _4172_ (.A0(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .S(clknet_1_1__leaf__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _4173_ (.A0(_1515_),
    .A1(_1516_),
    .S(clknet_1_1__leaf__1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(_1517_),
    .A1(_1514_),
    .S(clknet_1_1__leaf__1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(_1511_),
    .A1(_1518_),
    .S(_1507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1519_));
 sky130_fd_sc_hd__nand2_4 _4177_ (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .B(_1519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4178_ (.A1(_0078_),
    .A2(clknet_1_0__leaf__0805_),
    .B1(\dut_0.U0_formal_verification.cby_1__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1520_));
 sky130_fd_sc_hd__a21o_2 _4179_ (.A1(_0078_),
    .A2(clknet_1_0__leaf__0704_),
    .B1(_1520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4180_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(net346),
    .B1(\dut_0.U0_formal_verification.cbx_1__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1521_));
 sky130_fd_sc_hd__a21o_2 _4181_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_2.DFF_0_.Q ),
    .A2(net300),
    .B1(_1521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4182_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(net363),
    .B1(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1522_));
 sky130_fd_sc_hd__a21o_2 _4183_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .B1(_1522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_1 _4184_ (.A1(_0079_),
    .A2(clknet_1_0__leaf_net35),
    .B1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1523_));
 sky130_fd_sc_hd__a21o_2 _4185_ (.A1(_0079_),
    .A2(clknet_1_0__leaf__0700_),
    .B1(_1523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(clknet_1_1__leaf__0829_),
    .A1(clknet_1_0__leaf__0593_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1524_));
 sky130_fd_sc_hd__nand2_2 _4187_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_1_.Q ),
    .B(_1524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _4188_ (.A(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1525_));
 sky130_fd_sc_hd__o2111a_2 _4189_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0813_),
    .B1(_1525_),
    .C1(_0081_),
    .D1(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(clknet_1_0__leaf__0525_),
    .A1(clknet_1_0__leaf__1314_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(clknet_1_0__leaf__0544_),
    .A1(clknet_1_0__leaf__0646_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(_1528_),
    .A1(_1527_),
    .S(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1529_));
 sky130_fd_sc_hd__a21oi_2 _4193_ (.A1(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_2_.Q ),
    .A2(_1529_),
    .B1(_1526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(_0686_),
    .A1(clknet_1_0__leaf__0688_),
    .S(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1530_));
 sky130_fd_sc_hd__nor2_2 _4195_ (.A(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1531_));
 sky130_fd_sc_hd__a211o_2 _4196_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0193_),
    .B1(_1531_),
    .C1(_0082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1532_));
 sky130_fd_sc_hd__o211ai_2 _4197_ (.A1(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_1_.Q ),
    .A2(_1530_),
    .B1(_1532_),
    .C1(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1533_));
 sky130_fd_sc_hd__o41a_2 _4198_ (.A1(_0082_),
    .A2(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .A3(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_2_.Q ),
    .A4(clknet_1_1__leaf__0634_),
    .B1(_1533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _4199_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .B(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1534_));
 sky130_fd_sc_hd__o2111a_2 _4200_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0655_),
    .B1(_1534_),
    .C1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_1_.Q ),
    .D1(_0083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1535_));
 sky130_fd_sc_hd__nor2_2 _4201_ (.A(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1536_));
 sky130_fd_sc_hd__a211o_2 _4202_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0603_),
    .B1(_1536_),
    .C1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1537_));
 sky130_fd_sc_hd__o21ai_2 _4203_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .B1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1538_));
 sky130_fd_sc_hd__a21o_2 _4204_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0675_),
    .B1(_1538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1539_));
 sky130_fd_sc_hd__a31oi_2 _4205_ (.A1(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_2_.Q ),
    .A2(_1537_),
    .A3(_1539_),
    .B1(_1535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _4206_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1540_));
 sky130_fd_sc_hd__o2111a_2 _4207_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0811_),
    .B1(_1540_),
    .C1(_0085_),
    .D1(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(clknet_1_0__leaf__0257_),
    .A1(clknet_1_0__leaf__1316_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(clknet_1_0__leaf__0537_),
    .A1(clknet_1_0__leaf__0648_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(_1542_),
    .A1(_1543_),
    .S(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1544_));
 sky130_fd_sc_hd__a21oi_2 _4211_ (.A1(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_2_.Q ),
    .A2(_1544_),
    .B1(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__mux4_1 _4212_ (.A0(clknet_1_0__leaf_net49),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net52),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1545_));
 sky130_fd_sc_hd__nor2_1 _4213_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1546_));
 sky130_fd_sc_hd__a211o_1 _4214_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .A2(net21),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .C1(_0106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1547_));
 sky130_fd_sc_hd__o22a_1 _4215_ (.A1(_0107_),
    .A2(_1545_),
    .B1(_1546_),
    .B2(_1547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1548_));
 sky130_fd_sc_hd__mux4_2 _4216_ (.A0(clknet_1_1__leaf_net22),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1549_));
 sky130_fd_sc_hd__mux4_2 _4217_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1550_));
 sky130_fd_sc_hd__a21bo_2 _4218_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .A2(_1550_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1551_));
 sky130_fd_sc_hd__a21o_2 _4219_ (.A1(_0107_),
    .A2(_1549_),
    .B1(_1551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1552_));
 sky130_fd_sc_hd__o21ai_2 _4220_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .A2(_1548_),
    .B1(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1553_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(clknet_1_0__leaf_net49),
    .A1(clknet_1_0__leaf_net52),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1554_));
 sky130_fd_sc_hd__or3_1 _4222_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .B(_0105_),
    .C(_1554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1555_));
 sky130_fd_sc_hd__mux4_2 _4223_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net20),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1556_));
 sky130_fd_sc_hd__inv_2 _4280__171 (.A(_1610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net406));
 sky130_fd_sc_hd__a21oi_2 _4225_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .A2(net405),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1558_));
 sky130_fd_sc_hd__mux4_2 _4226_ (.A0(clknet_1_0__leaf_net22),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1559_));
 sky130_fd_sc_hd__mux4_2 _4227_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1560_));
 sky130_fd_sc_hd__or2_2 _4228_ (.A(_0105_),
    .B(_1560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1561_));
 sky130_fd_sc_hd__o211a_2 _4229_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .A2(_1559_),
    .B1(_1561_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1562_));
 sky130_fd_sc_hd__a21oi_2 _4230_ (.A1(_1555_),
    .A2(_1558_),
    .B1(_1562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_1 _4231_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_0__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1564_));
 sky130_fd_sc_hd__mux4_2 _4232_ (.A0(clknet_1_0__leaf_net50),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net53),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1565_));
 sky130_fd_sc_hd__nor2_1 _4233_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1566_));
 sky130_fd_sc_hd__a211o_1 _4234_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .A2(net20),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .C1(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1567_));
 sky130_fd_sc_hd__o22a_2 _4235_ (.A1(_0109_),
    .A2(_1565_),
    .B1(_1566_),
    .B2(_1567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1568_));
 sky130_fd_sc_hd__nor2_2 _4236_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .B(_1568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1569_));
 sky130_fd_sc_hd__mux4_2 _4237_ (.A0(clknet_1_0__leaf_net22),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1570_));
 sky130_fd_sc_hd__nand2_2 _4238_ (.A(_0109_),
    .B(_1570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1571_));
 sky130_fd_sc_hd__mux4_2 _4239_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1572_));
 sky130_fd_sc_hd__nand2_2 _4240_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .B(_1572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1573_));
 sky130_fd_sc_hd__a31o_2 _4241_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .A2(_1571_),
    .A3(_1573_),
    .B1(_1569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_0__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1575_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(_1564_),
    .A1(_1575_),
    .S(clknet_1_0__leaf__1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1576_));
 sky130_fd_sc_hd__nand2b_1 _4244_ (.A_N(_1576_),
    .B(clknet_1_0__leaf__1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1577_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_0__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_0__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(_1578_),
    .A1(_1579_),
    .S(clknet_1_0__leaf__1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1580_));
 sky130_fd_sc_hd__mux4_2 _4248_ (.A0(clknet_1_0__leaf_net50),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net53),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1581_));
 sky130_fd_sc_hd__nor2_1 _4249_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1582_));
 sky130_fd_sc_hd__a211o_1 _4250_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .A2(net20),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .C1(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1583_));
 sky130_fd_sc_hd__o22a_2 _4251_ (.A1(_0111_),
    .A2(_1581_),
    .B1(_1582_),
    .B2(_1583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1584_));
 sky130_fd_sc_hd__mux4_2 _4252_ (.A0(clknet_1_0__leaf_net22),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1585_));
 sky130_fd_sc_hd__mux4_2 _4253_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1586_));
 sky130_fd_sc_hd__a21bo_2 _4254_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .A2(_1586_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1587_));
 sky130_fd_sc_hd__a21o_2 _4255_ (.A1(_0111_),
    .A2(_1585_),
    .B1(_1587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1588_));
 sky130_fd_sc_hd__o21ai_2 _4256_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.ccff_tail ),
    .A2(_1584_),
    .B1(_1588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1589_));
 sky130_fd_sc_hd__o21ba_2 _4257_ (.A1(clknet_1_0__leaf__1574_),
    .A2(_1580_),
    .B1_N(clknet_1_1__leaf__1589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_1__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_1__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(_1591_),
    .A1(_1592_),
    .S(clknet_1_1__leaf__1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1593_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_1__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_1__leaf__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(_1595_),
    .A1(_1594_),
    .S(clknet_1_1__leaf__1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1596_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(_1596_),
    .A1(_1593_),
    .S(clknet_1_1__leaf__1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1597_));
 sky130_fd_sc_hd__a22o_1 _4265_ (.A1(_1577_),
    .A2(_1590_),
    .B1(_1597_),
    .B2(clknet_1_0__leaf__1589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1598_));
 sky130_fd_sc_hd__nand2_4 _4267_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .B(_1598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux4_2 _4268_ (.A0(clknet_1_0__leaf_net50),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net53),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1599_));
 sky130_fd_sc_hd__nor2_1 _4269_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1600_));
 sky130_fd_sc_hd__a211o_1 _4270_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(net20),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .C1(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1601_));
 sky130_fd_sc_hd__o22a_2 _4271_ (.A1(_0088_),
    .A2(_1599_),
    .B1(_1600_),
    .B2(_1601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1602_));
 sky130_fd_sc_hd__mux4_2 _4272_ (.A0(clknet_1_0__leaf_net22),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1603_));
 sky130_fd_sc_hd__mux4_2 _4273_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1604_));
 sky130_fd_sc_hd__a21bo_2 _4274_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .A2(_1604_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1605_));
 sky130_fd_sc_hd__a21o_2 _4275_ (.A1(_0088_),
    .A2(_1603_),
    .B1(_1605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1606_));
 sky130_fd_sc_hd__o21ai_2 _4276_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .A2(_1602_),
    .B1(_1606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1607_));
 sky130_fd_sc_hd__mux2_1 _4277_ (.A0(clknet_1_0__leaf_net50),
    .A1(clknet_1_0__leaf_net53),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1608_));
 sky130_fd_sc_hd__or3_1 _4278_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .B(_0086_),
    .C(_1608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1609_));
 sky130_fd_sc_hd__mux4_2 _4279_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net20),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1610_));
 sky130_fd_sc_hd__inv_2 _2837__172 (.A(clknet_1_0__leaf__0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net407));
 sky130_fd_sc_hd__a21oi_2 _4281_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .A2(net406),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1612_));
 sky130_fd_sc_hd__mux4_2 _4282_ (.A0(clknet_1_0__leaf_net22),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1613_));
 sky130_fd_sc_hd__mux4_2 _4283_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1614_));
 sky130_fd_sc_hd__or2_2 _4284_ (.A(_0086_),
    .B(_1614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1615_));
 sky130_fd_sc_hd__o211a_2 _4285_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .A2(_1613_),
    .B1(_1615_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1616_));
 sky130_fd_sc_hd__a21oi_2 _4286_ (.A1(_1609_),
    .A2(_1612_),
    .B1(_1616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1617_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .S(clknet_1_1__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1618_));
 sky130_fd_sc_hd__mux4_2 _4288_ (.A0(clknet_1_0__leaf_net50),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net53),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1619_));
 sky130_fd_sc_hd__nor2_1 _4289_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1620_));
 sky130_fd_sc_hd__a211o_1 _4290_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(net20),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .C1(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1621_));
 sky130_fd_sc_hd__o22a_2 _4291_ (.A1(_0090_),
    .A2(_1619_),
    .B1(_1620_),
    .B2(_1621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1622_));
 sky130_fd_sc_hd__mux4_2 _4292_ (.A0(clknet_1_0__leaf_net22),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1623_));
 sky130_fd_sc_hd__mux4_2 _4293_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1624_));
 sky130_fd_sc_hd__a21bo_2 _4294_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .A2(_1624_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1625_));
 sky130_fd_sc_hd__a21o_2 _4295_ (.A1(_0090_),
    .A2(_1623_),
    .B1(_1625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1626_));
 sky130_fd_sc_hd__o21ai_2 _4296_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .A2(_1622_),
    .B1(_1626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1627_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .S(clknet_1_1__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(_1628_),
    .A1(_1618_),
    .S(clknet_1_1__leaf__1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .S(clknet_1_1__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .S(clknet_1_1__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(_1630_),
    .A1(_1631_),
    .S(clknet_1_1__leaf__1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1632_));
 sky130_fd_sc_hd__nand2b_2 _4302_ (.A_N(_1632_),
    .B(clknet_1_1__leaf__1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1633_));
 sky130_fd_sc_hd__mux4_2 _4303_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net20),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1634_));
 sky130_fd_sc_hd__or2_2 _4304_ (.A(_0091_),
    .B(_1634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(clknet_1_0__leaf_net49),
    .A1(clknet_1_0__leaf_net52),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1636_));
 sky130_fd_sc_hd__or3b_1 _4306_ (.A(_1636_),
    .B(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .C_N(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1637_));
 sky130_fd_sc_hd__a21oi_2 _4307_ (.A1(_1635_),
    .A2(_1637_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1638_));
 sky130_fd_sc_hd__or2_1 _4308_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1639_));
 sky130_fd_sc_hd__a21oi_2 _4309_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1640_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1641_));
 sky130_fd_sc_hd__inv_2 _3766__192 (.A(_1127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net427));
 sky130_fd_sc_hd__a221o_2 _4312_ (.A1(_1639_),
    .A2(_1640_),
    .B1(net426),
    .B2(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1644_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1645_));
 sky130_fd_sc_hd__o21a_2 _4315_ (.A1(_0091_),
    .A2(_1645_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1646_));
 sky130_fd_sc_hd__o21ai_2 _4316_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .A2(_1644_),
    .B1(_1646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1647_));
 sky130_fd_sc_hd__a31o_2 _4317_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .A2(_1643_),
    .A3(_1647_),
    .B1(_1638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1648_));
 sky130_fd_sc_hd__o21ba_2 _4318_ (.A1(clknet_1_0__leaf__1627_),
    .A2(_1629_),
    .B1_N(clknet_1_0__leaf__1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1649_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .S(clknet_1_0__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .S(clknet_1_0__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(_1650_),
    .A1(_1651_),
    .S(clknet_1_0__leaf__1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .S(clknet_1_0__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .S(clknet_1_0__leaf__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(_1654_),
    .A1(_1653_),
    .S(clknet_1_0__leaf__1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(_1655_),
    .A1(_1652_),
    .S(clknet_1_0__leaf__1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1656_));
 sky130_fd_sc_hd__a22o_2 _4326_ (.A1(_1633_),
    .A2(_1649_),
    .B1(_1656_),
    .B2(clknet_1_1__leaf__1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1657_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .B(_1657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4329_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0596_),
    .B1(\dut_0.U0_formal_verification.cby_2__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1658_));
 sky130_fd_sc_hd__a21o_2 _4330_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_2.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .B1(_1658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(clknet_1_1__leaf__0681_),
    .A1(clknet_1_1__leaf__0688_),
    .S(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_2 _4332_ (.A(\dut_0.U0_formal_verification.cbx_1__1__1_ccff_tail ),
    .B(_1659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4333_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(net333),
    .B1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1660_));
 sky130_fd_sc_hd__a21o_2 _4334_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .B1(_1660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4335_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0849_),
    .B1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1661_));
 sky130_fd_sc_hd__a21o_2 _4336_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_0_.Q ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .B1(_1661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(clknet_1_1__leaf__0233_),
    .A1(clknet_1_1__leaf__0846_),
    .S(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1662_));
 sky130_fd_sc_hd__nand2_2 _4338_ (.A(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_1_.Q ),
    .B(_1662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__nor2_1 _4339_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1663_));
 sky130_fd_sc_hd__a211o_2 _4340_ (.A1(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0718_),
    .B1(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_2_.Q ),
    .C1(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1664_));
 sky130_fd_sc_hd__nand2_2 _4341_ (.A(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1665_));
 sky130_fd_sc_hd__o211a_2 _4342_ (.A1(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__1091_),
    .B1(_1665_),
    .C1(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(clknet_1_0__leaf__0558_),
    .A1(clknet_1_1__leaf__0574_),
    .S(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1667_));
 sky130_fd_sc_hd__a21bo_2 _4344_ (.A1(_0113_),
    .A2(_1667_),
    .B1_N(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1668_));
 sky130_fd_sc_hd__o22a_4 _4345_ (.A1(_1663_),
    .A2(_1664_),
    .B1(_1666_),
    .B2(_1668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _4346_ (.A(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .B(clknet_1_0__leaf__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1669_));
 sky130_fd_sc_hd__o2111a_2 _4347_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0599_),
    .B1(_1669_),
    .C1(_0120_),
    .D1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1670_));
 sky130_fd_sc_hd__mux4_2 _4348_ (.A0(net273),
    .A1(net323),
    .A2(clknet_1_0__leaf__1095_),
    .A3(clknet_1_0__leaf__0868_),
    .S0(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1671_));
 sky130_fd_sc_hd__a21oi_2 _4349_ (.A1(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_2_.Q ),
    .A2(_1671_),
    .B1(_1670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(clknet_1_1__leaf__0227_),
    .A1(clknet_1_1__leaf__0615_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1672_));
 sky130_fd_sc_hd__mux2_1 _4351_ (.A0(clknet_1_1__leaf__0568_),
    .A1(clknet_1_1__leaf__0639_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1673_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(_1672_),
    .A1(_1673_),
    .S(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1674_));
 sky130_fd_sc_hd__nand2_1 _4353_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ),
    .B(clknet_1_1__leaf__0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1675_));
 sky130_fd_sc_hd__o2111a_2 _4354_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__1077_),
    .B1(_1675_),
    .C1(_0121_),
    .D1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1676_));
 sky130_fd_sc_hd__a21oi_2 _4355_ (.A1(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_2_.Q ),
    .A2(_1674_),
    .B1(_1676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__nand2_2 _4356_ (.A(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_0_.Q ),
    .B(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1677_));
 sky130_fd_sc_hd__o2111a_2 _4357_ (.A1(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0883_),
    .B1(_1677_),
    .C1(_0122_),
    .D1(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1678_));
 sky130_fd_sc_hd__mux4_2 _4358_ (.A0(clknet_1_1__leaf__0555_),
    .A1(clknet_1_1__leaf__0617_),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .S0(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1679_));
 sky130_fd_sc_hd__o21ba_2 _4359_ (.A1(_0122_),
    .A2(_1679_),
    .B1_N(_1678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__mux4_1 _4360_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net16),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1680_));
 sky130_fd_sc_hd__mux2_1 _4361_ (.A0(clknet_1_1__leaf_net23),
    .A1(net26),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1681_));
 sky130_fd_sc_hd__inv_2 _4362_ (.A(_1681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1682_));
 sky130_fd_sc_hd__a21oi_1 _4363_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .A2(_1682_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1683_));
 sky130_fd_sc_hd__a211oi_1 _4364_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .A2(_1680_),
    .B1(_1683_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1684_));
 sky130_fd_sc_hd__mux4_2 _4365_ (.A0(clknet_1_1__leaf_net27),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_2 _4366_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .B(_1685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1686_));
 sky130_fd_sc_hd__mux4_2 _4367_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1687_));
 sky130_fd_sc_hd__nand2b_2 _4368_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .B(_1687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1688_));
 sky130_fd_sc_hd__a31o_2 _4369_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .A2(_1686_),
    .A3(_1688_),
    .B1(_1684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1689_));
 sky130_fd_sc_hd__mux4_2 _4370_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net16),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1690_));
 sky130_fd_sc_hd__and2_2 _4371_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .B(_1690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1691_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(clknet_1_1__leaf_net23),
    .A1(net26),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1692_));
 sky130_fd_sc_hd__inv_2 _4373_ (.A(_1692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1693_));
 sky130_fd_sc_hd__a21oi_1 _4374_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .A2(_1693_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1694_));
 sky130_fd_sc_hd__mux4_2 _4375_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1695_));
 sky130_fd_sc_hd__mux4_2 _4376_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf_net27),
    .A2(clknet_1_1__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1696_));
 sky130_fd_sc_hd__and2b_2 _4377_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .B(_1696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1697_));
 sky130_fd_sc_hd__a21bo_2 _4378_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .A2(_1695_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1698_));
 sky130_fd_sc_hd__o32a_2 _4379_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .A2(_1691_),
    .A3(_1694_),
    .B1(_1697_),
    .B2(_1698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1699_));
 sky130_fd_sc_hd__mux2_1 _4380_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .S(clknet_1_1__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1701_));
 sky130_fd_sc_hd__mux2_1 _4382_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf_net16),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1702_));
 sky130_fd_sc_hd__o21a_1 _4383_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .A2(_1702_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1703_));
 sky130_fd_sc_hd__o21ai_2 _4384_ (.A1(_0136_),
    .A2(_1701_),
    .B1(_1703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1704_));
 sky130_fd_sc_hd__mux2_1 _4385_ (.A0(clknet_1_1__leaf_net23),
    .A1(net25),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1705_));
 sky130_fd_sc_hd__nor2_1 _4386_ (.A(_0136_),
    .B(_1705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1706_));
 sky130_fd_sc_hd__o21ba_1 _4387_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .A2(_1706_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1707_));
 sky130_fd_sc_hd__mux4_2 _4388_ (.A0(clknet_1_0__leaf_net27),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1708_));
 sky130_fd_sc_hd__nand2_2 _4389_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .B(_1708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1709_));
 sky130_fd_sc_hd__mux4_2 _4390_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1710_));
 sky130_fd_sc_hd__nand2_2 _4391_ (.A(_0136_),
    .B(_1710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1711_));
 sky130_fd_sc_hd__a32o_2 _4392_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .A2(_1709_),
    .A3(_1711_),
    .B1(_1704_),
    .B2(_1707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .S(clknet_1_1__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(_1700_),
    .A1(_1713_),
    .S(clknet_1_1__leaf__1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1714_));
 sky130_fd_sc_hd__nand2b_1 _4395_ (.A_N(_1714_),
    .B(clknet_1_0__leaf__1712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1715_));
 sky130_fd_sc_hd__mux2_1 _4396_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .S(clknet_1_0__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1716_));
 sky130_fd_sc_hd__mux2_1 _4397_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .S(clknet_1_0__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1717_));
 sky130_fd_sc_hd__mux2_1 _4398_ (.A0(_1717_),
    .A1(_1716_),
    .S(clknet_1_0__leaf__1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1718_));
 sky130_fd_sc_hd__or2_2 _4399_ (.A(clknet_1_1__leaf__1712_),
    .B(_1718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1719_));
 sky130_fd_sc_hd__mux4_2 _4400_ (.A0(clknet_1_0__leaf_net23),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net25),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _4401_ (.A0(net15),
    .A1(clknet_1_1__leaf_net16),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1721_));
 sky130_fd_sc_hd__or3b_1 _4402_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .B(_1721_),
    .C_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1722_));
 sky130_fd_sc_hd__o21a_2 _4403_ (.A1(_0137_),
    .A2(_1720_),
    .B1(_1722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1723_));
 sky130_fd_sc_hd__mux4_2 _4404_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_2 _4405_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .B(_1724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1725_));
 sky130_fd_sc_hd__mux4_2 _4406_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf_net27),
    .A2(clknet_1_0__leaf_net18),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net40 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net40));
 sky130_fd_sc_hd__o211a_2 _4408_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .A2(net428),
    .B1(_1725_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1728_));
 sky130_fd_sc_hd__o21ba_2 _4409_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.ccff_tail ),
    .A2(_1723_),
    .B1_N(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1729_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .S(clknet_1_0__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1730_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .S(clknet_1_0__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1731_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(_1730_),
    .A1(_1731_),
    .S(clknet_1_0__leaf__1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1732_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .S(clknet_1_1__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1733_));
 sky130_fd_sc_hd__mux2_1 _4414_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .S(clknet_1_1__leaf__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1734_));
 sky130_fd_sc_hd__mux2_1 _4415_ (.A0(_1733_),
    .A1(_1734_),
    .S(clknet_1_1__leaf__1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1735_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(_1735_),
    .A1(_1732_),
    .S(clknet_1_0__leaf__1712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1736_));
 sky130_fd_sc_hd__and2b_2 _4417_ (.A_N(clknet_1_0__leaf__1729_),
    .B(_1736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1737_));
 sky130_fd_sc_hd__a31o_1 _4418_ (.A1(_1715_),
    .A2(_1719_),
    .A3(clknet_1_1__leaf__1729_),
    .B1(_1737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1738_));
 sky130_fd_sc_hd__nand2_2 _4420_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .B(_1738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux4_2 _4421_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_0__leaf_net27),
    .A2(clknet_1_0__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1739_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1740_));
 sky130_fd_sc_hd__or2_2 _4423_ (.A(_0124_),
    .B(_1740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1741_));
 sky130_fd_sc_hd__mux2_1 _4424_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1742_));
 sky130_fd_sc_hd__o211a_2 _4425_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .A2(_1742_),
    .B1(_1741_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1743_));
 sky130_fd_sc_hd__a21bo_2 _4426_ (.A1(_0123_),
    .A2(_1739_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1744_));
 sky130_fd_sc_hd__mux4_2 _4427_ (.A0(net15),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net16),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1745_));
 sky130_fd_sc_hd__and2b_1 _4428_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .B(clknet_1_1__leaf_net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1746_));
 sky130_fd_sc_hd__a211o_1 _4429_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .A2(net25),
    .B1(_0124_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1747_));
 sky130_fd_sc_hd__o22a_2 _4430_ (.A1(_0123_),
    .A2(_1745_),
    .B1(_1746_),
    .B2(_1747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1748_));
 sky130_fd_sc_hd__o22ai_2 _4431_ (.A1(_1743_),
    .A2(_1744_),
    .B1(_1748_),
    .B2(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1749_));
 sky130_fd_sc_hd__mux4_2 _4432_ (.A0(net15),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net17),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(clknet_1_1__leaf_net23),
    .A1(net25),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1751_));
 sky130_fd_sc_hd__inv_2 _4434_ (.A(_1751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1752_));
 sky130_fd_sc_hd__a21oi_1 _4435_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .A2(_1752_),
    .B1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1753_));
 sky130_fd_sc_hd__and2_2 _4436_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .B(_1750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1754_));
 sky130_fd_sc_hd__mux4_2 _4437_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1755_));
 sky130_fd_sc_hd__mux4_2 _4438_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(clknet_1_1__leaf_net27),
    .A2(clknet_1_1__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1756_));
 sky130_fd_sc_hd__and2b_2 _4439_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .B(_1756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1757_));
 sky130_fd_sc_hd__a21bo_2 _4440_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .A2(_1755_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1758_));
 sky130_fd_sc_hd__o32a_2 _4441_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .A2(_1753_),
    .A3(_1754_),
    .B1(_1757_),
    .B2(_1758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1759_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .S(clknet_1_1__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1760_));
 sky130_fd_sc_hd__mux4_2 _4443_ (.A0(net24),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A2(net25),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1761_));
 sky130_fd_sc_hd__nand2_1 _4444_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .B(clknet_1_0__leaf_net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1762_));
 sky130_fd_sc_hd__o211a_1 _4445_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .A2(clknet_1_1__leaf__0192_),
    .B1(_1762_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1763_));
 sky130_fd_sc_hd__nor2_1 _4446_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .B(_1763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1764_));
 sky130_fd_sc_hd__a211oi_2 _4447_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .A2(_1761_),
    .B1(_1764_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1765_));
 sky130_fd_sc_hd__mux4_2 _4448_ (.A0(clknet_1_0__leaf_net28),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_2 _4449_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .B(_1766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1767_));
 sky130_fd_sc_hd__mux4_2 _4450_ (.A0(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_0__leaf_net19),
    .A3(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1768_));
 sky130_fd_sc_hd__nand2b_2 _4451_ (.A_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .B(_1768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1769_));
 sky130_fd_sc_hd__a31o_2 _4452_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .A2(_1767_),
    .A3(_1769_),
    .B1(_1765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_1 _4453_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .S(clknet_1_1__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1771_));
 sky130_fd_sc_hd__mux2_1 _4454_ (.A0(_1760_),
    .A1(_1771_),
    .S(clknet_1_1__leaf__1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1772_));
 sky130_fd_sc_hd__mux4_2 _4455_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .A2(clknet_1_1__leaf_net18),
    .A3(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .S0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .S1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1773_));
 sky130_fd_sc_hd__mux2_1 _4456_ (.A0(clknet_1_0__leaf_net27),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1774_));
 sky130_fd_sc_hd__or2_1 _4457_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .B(_1774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1776_));
 sky130_fd_sc_hd__o211a_1 _4459_ (.A1(_0125_),
    .A2(_1776_),
    .B1(_1775_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1777_));
 sky130_fd_sc_hd__a21bo_2 _4460_ (.A1(_0126_),
    .A2(_1773_),
    .B1_N(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1778_));
 sky130_fd_sc_hd__mux2_1 _4461_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .A1(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1779_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(net15),
    .A1(net17),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1780_));
 sky130_fd_sc_hd__or2_1 _4463_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .B(_1780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1781_));
 sky130_fd_sc_hd__o211a_2 _4464_ (.A1(_0126_),
    .A2(_1779_),
    .B1(_1781_),
    .C1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1782_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(net24),
    .A1(net25),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1783_));
 sky130_fd_sc_hd__o21a_1 _4466_ (.A1(_0126_),
    .A2(_1783_),
    .B1(_0125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1784_));
 sky130_fd_sc_hd__o32a_1 _4467_ (.A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .A2(_1782_),
    .A3(_1784_),
    .B1(_1777_),
    .B2(_1778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1785_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .S(clknet_1_1__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .S(clknet_1_1__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(_1787_),
    .A1(_1786_),
    .S(clknet_1_1__leaf__1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1788_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(_1788_),
    .A1(_1772_),
    .S(clknet_1_1__leaf__1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1789_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .S(clknet_1_0__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1790_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .S(clknet_1_0__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1791_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(_1790_),
    .A1(_1791_),
    .S(clknet_1_0__leaf__1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .S(clknet_1_0__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1793_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .S(clknet_1_0__leaf__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1794_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(_1793_),
    .A1(_1794_),
    .S(clknet_1_0__leaf__1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1795_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(_1795_),
    .A1(_1792_),
    .S(clknet_1_0__leaf__1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1796_));
 sky130_fd_sc_hd__mux2_2 _4479_ (.A0(_1796_),
    .A1(_1789_),
    .S(_1785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .A1(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .S(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1797_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .B(_1797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__o21ai_2 _4482_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_2.DFF_0_.Q ),
    .A2(clknet_1_0__leaf__0668_),
    .B1(\dut_0.U0_formal_verification.cby_2__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1798_));
 sky130_fd_sc_hd__a21o_2 _4483_ (.A1(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_2.DFF_0_.Q ),
    .A2(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .B1(_1798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(net409),
    .A1(clknet_1_1__leaf__0593_),
    .S(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1799_));
 sky130_fd_sc_hd__nand2_2 _4485_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_ccff_tail ),
    .B(_1799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(net91),
    .D(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.cby_0__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.cby_0__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.cby_1__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(net170),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4525_ (.CLK_N(net244),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net221),
    .SET_B(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2157_));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(net179),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(net179),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4544_ (.CLK_N(net251),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net220),
    .SET_B(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2158_));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4563_ (.CLK_N(net241),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net220),
    .SET_B(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2159_));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(net214),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4582_ (.CLK_N(net242),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net221),
    .SET_B(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2160_));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4587_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4591_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4592_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(net173),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4595_ (.CLK(net171),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4596_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(net179),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(net179),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4599_ (.CLK(net179),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4600_ (.CLK(net173),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4603_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4604_ (.CLK(net179),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4607_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4608_ (.CLK(net180),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4611_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4612_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(net206),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4615_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4616_ (.CLK(net205),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(net206),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(net206),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4619_ (.CLK(net206),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4620_ (.CLK(net206),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4623_ (.CLK(net208),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4624_ (.CLK(net208),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4627_ (.CLK(net213),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4628_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4631_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4632_ (.CLK(net207),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4635_ (.CLK(net204),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4636_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4639_ (.CLK(net201),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4640_ (.CLK(net204),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4643_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4644_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_0_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4647_ (.CLK(net178),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4648_ (.CLK(net181),
    .D(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.cby_1__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4656_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4657_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4658_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4660_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(net60),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4665_ (.CLK_N(net236),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net222),
    .SET_B(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2161_));
 sky130_fd_sc_hd__dfxtp_1 _4666_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(net58),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(net59),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(net58),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(net58),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(net58),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(net56),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4684_ (.CLK_N(net237),
    .D(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net222),
    .SET_B(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2162_));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4689_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4703_ (.CLK_N(net238),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net222),
    .SET_B(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2163_));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(net77),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(net85),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4720_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4721_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4722_ (.CLK_N(net239),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net222),
    .SET_B(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2164_));
 sky130_fd_sc_hd__dfxtp_1 _4723_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4724_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4725_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4726_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4728_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4729_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4730_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4731_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4732_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4733_ (.CLK(net60),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4734_ (.CLK(net60),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4735_ (.CLK(net60),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4736_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4737_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4738_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4739_ (.CLK(net60),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4740_ (.CLK(net60),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4741_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4742_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4743_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4744_ (.CLK(net58),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4745_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4746_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4747_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4748_ (.CLK(net58),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4749_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4750_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4751_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4752_ (.CLK(net57),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4753_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4754_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4755_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4756_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4757_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4758_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4759_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4760_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4761_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4762_ (.CLK(net78),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4763_ (.CLK(net78),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4764_ (.CLK(net76),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4765_ (.CLK(net78),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4766_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4767_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4768_ (.CLK(net78),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4769_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4770_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4771_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4772_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4773_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4774_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4775_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4776_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4777_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4778_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4779_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4780_ (.CLK(net82),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4781_ (.CLK(net85),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4782_ (.CLK(net85),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4783_ (.CLK(net85),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4784_ (.CLK(net81),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4785_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4786_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4787_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4788_ (.CLK(net83),
    .D(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4789_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.cby_2__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4790_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4791_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4792_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4793_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4794_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4795_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4796_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4797_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4798_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4799_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4800_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4801_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4802_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4803_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4804_ (.CLK(net187),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4805_ (.CLK_N(net245),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net219),
    .SET_B(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2165_));
 sky130_fd_sc_hd__dfxtp_1 _4806_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4807_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4808_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4809_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4810_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4811_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4812_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4813_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4814_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4815_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4816_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4817_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4818_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4819_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4820_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4821_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4822_ (.CLK(net198),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4823_ (.CLK(net199),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4824_ (.CLK_N(net240),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net219),
    .SET_B(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2166_));
 sky130_fd_sc_hd__dfxtp_1 _4825_ (.CLK(net199),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4826_ (.CLK(net199),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4827_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4828_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4829_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4830_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4831_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4832_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4833_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4834_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4835_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4836_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4837_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4838_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4839_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4840_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4841_ (.CLK(net215),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4842_ (.CLK(net216),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4843_ (.CLK_N(net250),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net220),
    .SET_B(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2167_));
 sky130_fd_sc_hd__dfxtp_1 _4844_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4845_ (.CLK(net210),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4846_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4847_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4848_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4849_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4850_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4851_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4852_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4853_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4854_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4855_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4856_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4857_ (.CLK(net196),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4858_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4859_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4860_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4861_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4862_ (.CLK_N(net246),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net220),
    .SET_B(_0022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2168_));
 sky130_fd_sc_hd__dfxtp_1 _4863_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4864_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4865_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4866_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4867_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4868_ (.CLK(net162),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4869_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4870_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4871_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4872_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4873_ (.CLK(net204),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4874_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4875_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4876_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4877_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4878_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4879_ (.CLK(net204),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4880_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4881_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4882_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4883_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4884_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4885_ (.CLK(net199),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4886_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4887_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4888_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4889_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4890_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4891_ (.CLK(net199),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4892_ (.CLK(net199),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4893_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4894_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4895_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4896_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4897_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4898_ (.CLK(net216),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4899_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4900_ (.CLK(net212),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4901_ (.CLK(net210),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4902_ (.CLK(net210),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4903_ (.CLK(net210),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4904_ (.CLK(net211),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4905_ (.CLK(net210),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4906_ (.CLK(net204),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4907_ (.CLK(net204),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4908_ (.CLK(net210),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4909_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4910_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4911_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4912_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4913_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4914_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4915_ (.CLK(net203),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4916_ (.CLK(net209),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4917_ (.CLK(net197),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4918_ (.CLK(net200),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4919_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4920_ (.CLK(net190),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4921_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4922_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4923_ (.CLK(net202),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4924_ (.CLK(net191),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4925_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4926_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _4927_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4928_ (.CLK(net176),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4929_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.cby_2__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4930_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4931_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4932_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4933_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4934_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4935_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4936_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4937_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4938_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4939_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4940_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4941_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4942_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4943_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4944_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4945_ (.CLK_N(net247),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net220),
    .SET_B(_0024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2169_));
 sky130_fd_sc_hd__dfxtp_1 _4946_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4947_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4948_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4949_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4950_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4951_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4952_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4953_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4954_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4955_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4956_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4957_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4958_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4959_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4960_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4961_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4962_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4963_ (.CLK(net192),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4964_ (.CLK_N(net248),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net219),
    .SET_B(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2170_));
 sky130_fd_sc_hd__dfxtp_1 _4965_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4966_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4967_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4968_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4969_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4970_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4971_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4972_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4973_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4974_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4975_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4976_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4977_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4978_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4979_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4980_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4981_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4982_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _4983_ (.CLK_N(net243),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net221),
    .SET_B(_0028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2171_));
 sky130_fd_sc_hd__dfxtp_1 _4984_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _4985_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4986_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4987_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4988_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4989_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4990_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4991_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4992_ (.CLK(net195),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4993_ (.CLK(net195),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4994_ (.CLK(net195),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4995_ (.CLK(net195),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4996_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4997_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4998_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _4999_ (.CLK(net194),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _5000_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _5001_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfbbn_2 _5002_ (.CLK_N(net249),
    .D(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(net219),
    .SET_B(_0030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(_2172_));
 sky130_fd_sc_hd__dfxtp_1 _5003_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5004_ (.CLK(net193),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5005_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5006_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5007_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5008_ (.CLK(net189),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5009_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5010_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5011_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5012_ (.CLK(net188),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5013_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5014_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5015_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5016_ (.CLK(net161),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5017_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5018_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5019_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5020_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5021_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5022_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5023_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5024_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5025_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5026_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5027_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5028_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5029_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5030_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5031_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5032_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5033_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5034_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5035_ (.CLK(net155),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5036_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5037_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5038_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5039_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5040_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5041_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5042_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5043_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5044_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5045_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5046_ (.CLK(net154),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5047_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5048_ (.CLK(net146),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5049_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5050_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5051_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5052_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5053_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5054_ (.CLK(net185),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5055_ (.CLK(net186),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5056_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5057_ (.CLK(net184),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5058_ (.CLK(net186),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5059_ (.CLK(net186),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5060_ (.CLK(net186),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5061_ (.CLK(net184),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5062_ (.CLK(net184),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5063_ (.CLK(net183),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5064_ (.CLK(net184),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5065_ (.CLK(net156),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5066_ (.CLK(net157),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5067_ (.CLK(net157),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5068_ (.CLK(net184),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5069_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5070_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5071_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5072_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_14.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5073_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5074_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_12.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5075_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5076_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5077_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5078_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_10.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5079_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5080_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5081_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5082_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5083_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5084_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5085_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5086_ (.CLK(net95),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5087_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5088_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_right_track_0.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5089_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5090_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_14.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5091_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5092_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_12.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5093_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5094_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5095_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5096_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_10.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5097_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5098_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5099_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5100_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5101_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5102_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5103_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5104_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__0_.mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5105_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_14.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5106_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5107_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5108_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5109_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5110_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_12.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5111_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5112_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_10.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5113_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5114_ (.CLK(net88),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5115_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5116_ (.CLK(net88),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5117_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5118_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5119_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5120_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5121_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5122_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5123_ (.CLK(net97),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5124_ (.CLK(net88),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5125_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5126_ (.CLK(net89),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5127_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5128_ (.CLK(net90),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5129_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5130_ (.CLK(net97),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_bottom_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5131_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5132_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5133_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5134_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_right_track_2.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5135_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5136_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5137_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5138_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5139_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5140_ (.CLK(net75),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5141_ (.CLK(net75),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5142_ (.CLK(net75),
    .D(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.mem_top_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5143_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5144_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__1_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5145_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5146_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_15.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5147_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5148_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_13.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5149_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5150_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5151_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5152_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_11.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5153_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5154_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5155_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5156_ (.CLK(net71),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5157_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5158_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5159_ (.CLK(net73),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5160_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5161_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5162_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_bottom_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5163_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5164_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_14.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5165_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5166_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_12.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5167_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5168_ (.CLK(net74),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5169_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5170_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_10.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5171_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5172_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5173_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5174_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5175_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5176_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5177_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.grid_io_top_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5178_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_0__2_.mem_right_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5179_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5180_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5181_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5182_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5183_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5184_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5185_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5186_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5187_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5188_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5189_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5190_ (.CLK(net130),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5191_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5192_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5193_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5194_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_left_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5195_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5196_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5197_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5198_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5199_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5200_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5201_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5202_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5203_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5204_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5205_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_right_track_0.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5206_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5207_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5208_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5209_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_14.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5210_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5211_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5212_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.grid_io_left_0__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5213_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5214_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__0_.mem_top_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5215_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5216_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5217_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5218_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5219_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5220_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5221_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5222_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5223_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5224_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5225_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5226_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5227_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5228_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5229_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5230_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5231_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5232_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5233_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5234_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5235_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5236_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5237_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5238_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_left_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5239_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5240_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5241_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5242_ (.CLK(net123),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5243_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5244_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5245_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5246_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_bottom_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5247_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5248_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5249_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5250_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5251_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5252_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5253_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5254_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_right_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5255_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5256_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5257_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5258_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5259_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5260_ (.CLK(net108),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5261_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5262_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__1_.mem_top_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5263_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5264_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5265_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5266_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_15.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5267_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5268_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_13.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5269_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5270_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5271_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5272_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_11.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5273_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5274_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5275_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5276_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5277_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5278_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5279_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5280_ (.CLK(net104),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5281_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5282_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5283_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5284_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5285_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5286_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5287_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5288_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5289_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5290_ (.CLK(net104),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5291_ (.CLK(net103),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5292_ (.CLK(net100),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_left_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5293_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5294_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5295_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5296_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_bottom_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5297_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5298_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5299_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5300_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5301_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.grid_io_top_1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5302_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5303_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5304_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_1__2_.mem_right_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5305_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5306_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5307_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5308_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_15.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5309_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5310_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_13.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5311_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5312_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5313_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5314_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_11.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5315_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5316_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5317_ (.CLK(net138),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5318_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5319_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5320_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5321_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5322_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5323_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5324_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5325_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5326_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_14.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5327_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5328_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_12.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5329_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5330_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5331_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5332_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_10.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5333_ (.CLK(net135),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5334_ (.CLK(net135),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5335_ (.CLK(net164),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5336_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5337_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5338_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5339_ (.CLK(net177),
    .D(\dut_0.U0_formal_verification.grid_clb_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5340_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__0_.mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5341_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5342_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5343_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5344_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_15.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5345_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5346_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_13.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5347_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5348_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5349_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5350_ (.CLK(net119),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_11.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5351_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5352_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5353_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5354_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5355_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5356_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5357_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5358_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5359_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5360_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5361_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5362_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5363_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5364_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5365_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5366_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_9.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5367_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5368_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5369_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5370_ (.CLK(net165),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5371_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5372_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5373_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5374_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_bottom_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5375_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_3_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5376_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5377_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5378_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_8.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5379_ (.CLK(net160),
    .D(\dut_0.U0_formal_verification.grid_clb_2__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5380_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5381_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5382_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__1_.mem_top_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5383_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5384_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 _5385_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5386_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_15.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5387_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5388_ (.CLK(net111),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_13.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5389_ (.CLK(net114),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5390_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5391_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5392_ (.CLK(net114),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_11.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5393_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5394_ (.CLK(net112),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5395_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5396_ (.CLK(net114),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5397_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5398_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5399_ (.CLK(net145),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5400_ (.CLK(net145),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5401_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5402_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5403_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5404_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_15.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5405_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5406_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5407_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5408_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5409_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5410_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_11.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _5411_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5412_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5413_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5414_ (.CLK(net119),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5415_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5416_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5417_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.grid_io_right_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5418_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5419_ (.CLK(net127),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5420_ (.CLK(net129),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5421_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5422_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5423_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5424_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5425_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5426_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5427_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5428_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5429_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5430_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5431_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5432_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5433_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5434_ (.CLK(net128),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5435_ (.CLK(net129),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5436_ (.CLK(net96),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5437_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5438_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5439_ (.CLK(net96),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5440_ (.CLK(net96),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5441_ (.CLK(net96),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5442_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5443_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5444_ (.CLK(net92),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_top_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5445_ (.CLK(net129),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5446_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5447_ (.CLK(net92),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5448_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5449_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5450_ (.CLK(net125),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5451_ (.CLK(net170),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5452_ (.CLK(net170),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5453_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5454_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5455_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__0__1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5456_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5457_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5458_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5459_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5460_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5461_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5462_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5463_ (.CLK(net137),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5464_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5465_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5466_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5467_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5468_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5469_ (.CLK(net140),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5470_ (.CLK(net140),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5471_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5472_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5473_ (.CLK(net139),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5474_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5475_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5476_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_top_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5477_ (.CLK(net170),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5478_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5479_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5480_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5481_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5482_ (.CLK(net169),
    .D(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5483_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5484_ (.CLK(net134),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5485_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5486_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5487_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5488_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5489_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5490_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5491_ (.CLK(net131),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_top_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5492_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5493_ (.CLK(net121),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5494_ (.CLK(net122),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5495_ (.CLK(net109),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5496_ (.CLK(net109),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5497_ (.CLK(net109),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5498_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5499_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__1__1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5500_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5501_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5502_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5503_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5504_ (.CLK(net119),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5505_ (.CLK(net119),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5506_ (.CLK(net149),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_top_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5507_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5508_ (.CLK(net117),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5509_ (.CLK(net118),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5510_ (.CLK(net120),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5511_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5512_ (.CLK(net115),
    .D(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5513_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5514_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5515_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5516_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5517_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5518_ (.CLK(net70),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5519_ (.CLK(net70),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_top_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5520_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5521_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5522_ (.CLK(net101),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_7.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5523_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5524_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5525_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5526_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5527_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5528_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5529_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5530_ (.CLK(net66),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5531_ (.CLK(net67),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5532_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5533_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5534_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5535_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5536_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5537_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5538_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5539_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5540_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5541_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5542_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5543_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5544_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5545_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_1__2__1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5546_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5547_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5548_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5549_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5550_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_top_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5551_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5552_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5553_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_7.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5554_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5555_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5556_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5557_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5558_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5559_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5560_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5561_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5562_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5563_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5564_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5565_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5566_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5567_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5568_ (.CLK(net110),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5569_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5570_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5571_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5572_ (.CLK(net144),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5573_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5574_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5575_ (.CLK(net92),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5576_ (.CLK(net94),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5577_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5578_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5579_ (.CLK(net91),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5580_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5581_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5582_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5583_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5584_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5585_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5586_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5587_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5588_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5589_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5590_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5591_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5592_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5593_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5594_ (.CLK(net87),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5595_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5596_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5597_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5598_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5599_ (.CLK(net80),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5600_ (.CLK(net84),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_right_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5601_ (.CLK(net93),
    .D(\dut_0.U0_formal_verification.cby_0__1_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5602_ (.CLK(net92),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5603_ (.CLK(net92),
    .D(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1_.mem_left_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5604_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5605_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5606_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5607_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5608_ (.CLK(net62),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__1__1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5609_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5610_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5611_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5612_ (.CLK(net72),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5613_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5614_ (.CLK(net86),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5615_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5616_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5617_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5618_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5619_ (.CLK(net61),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5620_ (.CLK(net63),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5621_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5622_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5623_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5624_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5625_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5626_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5627_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5628_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5629_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_right_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5630_ (.CLK(net79),
    .D(\dut_0.U0_formal_verification.cby_0__2_.ccff_head ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5631_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5632_ (.CLK(net64),
    .D(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_0__2_.mem_left_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5633_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5634_ (.CLK(net170),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5635_ (.CLK(net135),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5636_ (.CLK(net168),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5637_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5638_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5639_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5640_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5641_ (.CLK(net133),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_right_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5642_ (.CLK(net129),
    .D(\dut_0.U0_formal_verification.cbx_1__0_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5643_ (.CLK(net124),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5644_ (.CLK(net132),
    .D(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1_.mem_left_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5645_ (.CLK(net105),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5646_ (.CLK(net101),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__1__1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5647_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5648_ (.CLK(net106),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5649_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5650_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _5651_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5652_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5653_ (.CLK(net107),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_right_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5654_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cbx_1__1_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5655_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5656_ (.CLK(net116),
    .D(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_1__2_.mem_left_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5657_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5658_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5659_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5660_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5661_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5662_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5663_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_right_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5664_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5665_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5666_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_7.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5667_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5668_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5669_ (.CLK(net166),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5670_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5671_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5672_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5673_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5674_ (.CLK(net174),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5675_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5676_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5677_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5678_ (.CLK(net175),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5679_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5680_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5681_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5682_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5683_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5684_ (.CLK(net150),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5685_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.cbx_1__0__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5686_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5687_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1_.mem_left_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5688_ (.CLK(net157),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5689_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__1__1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5690_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5691_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5692_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5693_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5694_ (.CLK(net153),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_right_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5695_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5696_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5697_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_7.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5698_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5699_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5700_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_6.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5701_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5702_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5703_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_5.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5704_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5705_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5706_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_4.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5707_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5708_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5709_ (.CLK(net147),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5710_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5711_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5712_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5713_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5714_ (.CLK(net159),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5715_ (.CLK(net162),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5716_ (.CLK(net152),
    .D(\dut_0.U0_formal_verification.cbx_1__1__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5717_ (.CLK(net152),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5718_ (.CLK(net162),
    .D(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.cby_2__2_.mem_left_ipin_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _5719_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_0_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5720_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5721_ (.CLK(net69),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5722_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5723_ (.CLK(net101),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5724_ (.CLK(net99),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5725_ (.CLK(net70),
    .D(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5726_ (.CLK(net68),
    .D(\dut_0.U0_formal_verification.cbx_1__2_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5727_ (.CLK(net102),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5728_ (.CLK(net104),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5729_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5730_ (.CLK(net113),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5731_ (.CLK(net114),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5732_ (.CLK(net143),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5733_ (.CLK(net145),
    .D(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5734_ (.CLK(net145),
    .D(\dut_0.U0_formal_verification.cbx_1__2__1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5735_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_0_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5736_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5737_ (.CLK(net148),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5738_ (.CLK(net145),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5739_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5740_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5741_ (.CLK(net158),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5742_ (.CLK(net151),
    .D(\dut_0.U0_formal_verification.grid_io_right_1_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5743_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_1_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5744_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5745_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5746_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5747_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5748_ (.CLK(net167),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5749_ (.CLK(net172),
    .D(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5750_ (.CLK(net170),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_0_ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5751_ (.CLK(net140),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_0_ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5752_ (.CLK(net140),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5753_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5754_ (.CLK(net141),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5755_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5756_ (.CLK(net136),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5757_ (.CLK(net129),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5758_ (.CLK(net129),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _5759_ (.CLK(net126),
    .D(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.ccff_tail ));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net234));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net235));
 sky130_fd_sc_hd__inv_2 _2556__1 (.A(clknet_1_0__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net236));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net224));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net225));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net226));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net227));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net228));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net229));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net230));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net231));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net232));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net233));
 sky130_fd_sc_hd__buf_2 _5773_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__buf_2 _5774_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__buf_2 _5775_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__buf_2 _5776_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _5777_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _5778_ (.A(\dut_0.U0_formal_verification.ccff_tail ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _5779_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__clkbuf_4 _5780_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _5781_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _5782_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _5783_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__ebufn_1 _5784_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ ),
    .TE_B(_2029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5785_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_ ),
    .TE_B(_2030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5786_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ ),
    .TE_B(_2031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.RST ));
 sky130_fd_sc_hd__ebufn_2 _5787_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .TE_B(_2032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5788_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ ),
    .TE_B(_2033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net5));
 sky130_fd_sc_hd__ebufn_1 _5789_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ ),
    .TE_B(_2034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net3));
 sky130_fd_sc_hd__ebufn_1 _5790_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ ),
    .TE_B(_2035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net9));
 sky130_fd_sc_hd__ebufn_2 _5791_ (.A(net10),
    .TE_B(_2036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_1 _5792_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_4 _5793_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5794_ (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.RST ),
    .TE_B(_2039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5795_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5796_ (.A(net5),
    .TE_B(_2041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5797_ (.A(net3),
    .TE_B(_2042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_1 _5798_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_ ),
    .TE_B(_2043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net7));
 sky130_fd_sc_hd__ebufn_1 _5799_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_ ),
    .TE_B(_2044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5800_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_ ),
    .TE_B(_2045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(clk));
 sky130_fd_sc_hd__ebufn_2 _5801_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_ ),
    .TE_B(_2046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5802_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .TE_B(_2047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5803_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ ),
    .TE_B(_2048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5804_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ ),
    .TE_B(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5805_ (.A(\dut_0.U0_formal_verification.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ ),
    .TE_B(_2050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5806_ (.A(net7),
    .TE_B(_2051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5807_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5808_ (.A(clknet_1_1__leaf_net40),
    .TE_B(_2053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5809_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .TE_B(_2054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5810_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5811_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .TE_B(_2056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5812_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ),
    .TE_B(_2057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5813_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_ ),
    .TE_B(_2058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5814_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_ ),
    .TE_B(_2059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5815_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_ ),
    .TE_B(_2060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5816_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_ ),
    .TE_B(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5817_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .TE_B(_2062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5818_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ ),
    .TE_B(_2063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5819_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ ),
    .TE_B(_2064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5820_ (.A(\dut_0.U0_formal_verification.cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ ),
    .TE_B(_2065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5821_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .TE_B(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5822_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5823_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5824_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .TE_B(_2069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5825_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5826_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .TE_B(_2071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5827_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ),
    .TE_B(_2072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5828_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5829_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5830_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5831_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5832_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5833_ (.A(net9),
    .TE_B(_2078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5834_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_2 _5835_ (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .TE_B(_2080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__ebufn_1 _5836_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_7.out ),
    .TE_B(_2081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5837_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_6.out ),
    .TE_B(_2082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5838_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_5.out ),
    .TE_B(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5839_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_4.out ),
    .TE_B(_2084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5840_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_3.out ),
    .TE_B(_2085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5841_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.out ),
    .TE_B(_2086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5842_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.out ),
    .TE_B(_2087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5843_ (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_0.out ),
    .TE_B(_2088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5844_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .TE_B(_2089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5845_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5846_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_1 _5847_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .TE_B(_2092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5848_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5849_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .TE_B(_2094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5850_ (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ),
    .TE_B(_2095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5851_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_ ),
    .TE_B(_2096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5852_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_ ),
    .TE_B(_2097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5853_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_ ),
    .TE_B(_2098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5854_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_ ),
    .TE_B(_2099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5855_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .TE_B(_2100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5856_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_ ),
    .TE_B(_2101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5857_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_ ),
    .TE_B(_2102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5858_ (.A(\dut_0.U0_formal_verification.cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_ ),
    .TE_B(_2103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5859_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .TE_B(_2104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5860_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5861_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_1 _5862_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .TE_B(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5863_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5864_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .TE_B(_2109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5865_ (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ),
    .TE_B(_2110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5866_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_ ),
    .TE_B(_2111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_4 _5867_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_ ),
    .TE_B(_2112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5868_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_ ),
    .TE_B(_2113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5869_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_ ),
    .TE_B(_2114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5870_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .TE_B(_2115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5871_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_ ),
    .TE_B(_2116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5872_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_ ),
    .TE_B(_2117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5873_ (.A(\dut_0.U0_formal_verification.cby_2__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_ ),
    .TE_B(_2118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5874_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .TE_B(_2119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5875_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5876_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5877_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .TE_B(_2122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5878_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5879_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .TE_B(_2124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5880_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ),
    .TE_B(_2125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_4 _5881_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_7.out ),
    .TE_B(_2126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net11));
 sky130_fd_sc_hd__ebufn_4 _5882_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_6.out ),
    .TE_B(_2127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5883_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_5.out ),
    .TE_B(_2128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_4 _5884_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_4.out ),
    .TE_B(_2129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net6));
 sky130_fd_sc_hd__ebufn_2 _5885_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_3.out ),
    .TE_B(_2130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5886_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_2.out ),
    .TE_B(_2131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5887_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.out ),
    .TE_B(_2132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5888_ (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.out ),
    .TE_B(_2133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5889_ (.A(net11),
    .TE_B(_2134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5890_ (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_1 _5891_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_1 _5892_ (.A(net6),
    .TE_B(_2137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5893_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .TE_B(_2138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5894_ (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .TE_B(_2139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5895_ (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__1.gfpga_pad_GPIO_PAD ),
    .TE_B(_2140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5896_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_ ),
    .TE_B(_2141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5897_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ ),
    .TE_B(_2142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5898_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_ ),
    .TE_B(_2143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5899_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ ),
    .TE_B(_2144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_1 _5900_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .TE_B(_2145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net2));
 sky130_fd_sc_hd__ebufn_4 _5901_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ ),
    .TE_B(_2146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net4));
 sky130_fd_sc_hd__ebufn_2 _5902_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ ),
    .TE_B(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net8));
 sky130_fd_sc_hd__ebufn_2 _5903_ (.A(\dut_0.U0_formal_verification.cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ ),
    .TE_B(_2148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__ebufn_2 _5904_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .TE_B(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5905_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .TE_B(_2150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5906_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.gfpga_pad_GPIO_PAD ),
    .TE_B(_2151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5907_ (.A(\dut_0.U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.gfpga_pad_GPIO_PAD ),
    .TE_B(_2152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_2 _5908_ (.A(net2),
    .TE_B(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_4 _5909_ (.A(net4),
    .TE_B(_2154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_4 _5910_ (.A(net8),
    .TE_B(_2155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__ebufn_1 _5911_ (.A(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_ ),
    .TE_B(_2156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(net10));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(uio_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(uio_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(uio_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(uio_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_4 fanout15 (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_6 fanout17 (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(clknet_1_1__leaf_net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(\dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_6 fanout26 (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(clknet_1_1__leaf_net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(\dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_4 fanout37 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_6 fanout39 (.A(clknet_1_1__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_12 fanout43 (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(clknet_1_1__leaf_net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(clknet_1_1__leaf_net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout60 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout62 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout64 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 fanout66 (.A(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 fanout68 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 fanout70 (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout72 (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 fanout73 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 fanout76 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 fanout77 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout78 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 fanout80 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__buf_2 fanout82 (.A(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout85 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__buf_1 fanout88 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__buf_1 fanout92 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout96 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout101 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__buf_1 fanout104 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout109 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 fanout113 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 fanout115 (.A(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 fanout117 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 fanout119 (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 fanout122 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 fanout135 (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 fanout138 (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 fanout139 (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 fanout140 (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 fanout141 (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 fanout144 (.A(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 fanout147 (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 fanout148 (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 fanout150 (.A(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout152 (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 fanout154 (.A(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 fanout155 (.A(net156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout157 (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 fanout159 (.A(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 fanout161 (.A(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 fanout162 (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 fanout164 (.A(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 fanout165 (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 fanout166 (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 fanout167 (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 fanout168 (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 fanout171 (.A(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 fanout172 (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 fanout175 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 fanout176 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout177 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__buf_1 fanout179 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__buf_2 fanout181 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 fanout182 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__buf_1 fanout184 (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 fanout185 (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 fanout186 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 fanout187 (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 fanout188 (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 fanout189 (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 fanout190 (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout191 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 fanout192 (.A(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 fanout193 (.A(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__buf_1 fanout195 (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 fanout196 (.A(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 fanout197 (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout199 (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 fanout204 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout206 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 fanout207 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 fanout208 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__buf_1 fanout210 (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 fanout212 (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 fanout213 (.A(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 fanout216 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__conb_1 tt_um_openfpga22_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net223));
 sky130_fd_sc_hd__inv_2 _2798__20 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _2802__22 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _2802__23 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _2802__24 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _2802__25 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _2819__27 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _2819__28 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _2819__29 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _2819__30 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _2801__32 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _2801__33 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _2801__34 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _2801__35 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _2801__36 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _2796__38 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _2793__40 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _3257__42 (.A(clknet_1_0__leaf__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _3257__43 (.A(clknet_1_0__leaf__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _3257__44 (.A(clknet_1_1__leaf__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _2790__46 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _2816__52 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _2816__53 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _2816__54 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _2817__56 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _3360__58 (.A(clknet_1_0__leaf__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _3360__59 (.A(clknet_1_1__leaf__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _3360__60 (.A(clknet_1_1__leaf__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _3186__62 (.A(clknet_1_0__leaf__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _3186__63 (.A(clknet_1_0__leaf__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _3280__66 (.A(clknet_1_0__leaf__0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _2808__68 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _2808__69 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _2808__70 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _2808__71 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _2808__72 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _2808__73 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _3684__83 (.A(clknet_1_1__leaf__1049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _2815__85 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _2815__86 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _2815__87 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _2806__89 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _2806__90 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _2806__91 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _2806__92 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _2806__93 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _2806__94 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _2797__96 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _2811__99 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _2811__100 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _2811__101 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _2811__102 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _3741__104 (.A(clknet_1_1__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _3741__105 (.A(clknet_1_1__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _3741__106 (.A(clknet_1_1__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _3741__107 (.A(clknet_1_1__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _2818__110 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _2812__112 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _2812__113 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _2812__114 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _2812__115 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _2812__116 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _2812__117 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _2812__118 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _2803__129 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _2803__130 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _2810__132 (.A(clknet_1_0__leaf_net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _2820__134 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _2820__135 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _2820__136 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _2820__137 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _2820__138 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _2820__139 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _2805__142 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _2809__146 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _2809__147 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _2809__148 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _2809__149 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _2809__150 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _2809__151 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _2809__152 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _2809__153 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _2809__154 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _2809__155 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _2809__156 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _2814__159 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _2814__160 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _2814__161 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _2814__162 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _2814__163 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _2814__164 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _3296__167 (.A(clknet_1_0__leaf__0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _2837__173 (.A(clknet_1_0__leaf__0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _2813__175 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _2813__176 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _2813__177 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _2813__178 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _2813__179 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _2813__180 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _2813__181 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _3270__183 (.A(clknet_1_0__leaf__0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _3151__189 (.A(clknet_1_0__leaf__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _3151__190 (.A(clknet_1_0__leaf__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net425));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net40 (.A(clknet_0_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net40));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net40 (.A(clknet_0_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net40));
 sky130_fd_sc_hd__bufinv_8 clkload0 (.A(clknet_1_1__leaf_net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net39 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net39));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net39 (.A(clknet_0_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net39));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net39 (.A(clknet_0_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net39));
 sky130_fd_sc_hd__inv_4 clkload1 (.A(clknet_1_1__leaf_net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0698_ (.A(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0698_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0698_ (.A(clknet_0__0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0698_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0698_ (.A(clknet_0__0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0698_));
 sky130_fd_sc_hd__bufinv_16 clkload3 (.A(clknet_1_0__leaf__0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0757_ (.A(_0757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0757_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0757_ (.A(clknet_0__0757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0757_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0757_ (.A(clknet_0__0757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0757_));
 sky130_fd_sc_hd__bufinv_8 clkload6 (.A(clknet_1_0__leaf__0757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0820_ (.A(_0820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0820_ (.A(clknet_0__0820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0820_ (.A(clknet_0__0820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0820_));
 sky130_fd_sc_hd__clkbuf_4 clkload7 (.A(clknet_1_1__leaf__0820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload9 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1134_ (.A(_1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1134_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1134_ (.A(clknet_0__1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1134_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1134_ (.A(clknet_0__1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1134_));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_1_1__leaf__1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload11 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1214_ (.A(_1214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1214_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1214_ (.A(clknet_0__1214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1214_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1214_ (.A(clknet_0__1214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1214_));
 sky130_fd_sc_hd__clkbuf_4 clkload12 (.A(clknet_1_1__leaf__1214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload13 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__bufinv_8 clkload14 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net50 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net50));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net50 (.A(clknet_0_net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net50));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net50 (.A(clknet_0_net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net50));
 sky130_fd_sc_hd__clkinv_2 clkload15 (.A(clknet_1_1__leaf_net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net49 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net49 (.A(clknet_0_net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net49 (.A(clknet_0_net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net49));
 sky130_fd_sc_hd__inv_2 clkload16 (.A(clknet_1_0__leaf_net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1199_ (.A(_1199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1199_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1199_ (.A(clknet_0__1199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1199_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1199_ (.A(clknet_0__1199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1199_));
 sky130_fd_sc_hd__clkinv_2 clkload17 (.A(clknet_1_1__leaf__1199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1178_ (.A(_1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1178_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1178_ (.A(clknet_0__1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1178_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1178_ (.A(clknet_0__1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1178_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1149_ (.A(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1149_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1149_ (.A(clknet_0__1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1149_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1149_ (.A(clknet_0__1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1149_));
 sky130_fd_sc_hd__clkbuf_4 clkload18 (.A(clknet_1_0__leaf__1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1118_ (.A(_1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1118_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1118_ (.A(clknet_0__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1118_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1118_ (.A(clknet_0__1118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1118_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1108_ (.A(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1108_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1108_ (.A(clknet_0__1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1108_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1108_ (.A(clknet_0__1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1108_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1563_ (.A(_1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1563_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1563_ (.A(clknet_0__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1563_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1563_ (.A(clknet_0__1563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1563_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload19 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload20 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1553_ (.A(_1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1553_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1553_ (.A(clknet_0__1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1553_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1553_ (.A(clknet_0__1553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1553_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1574_ (.A(_1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1574_ (.A(clknet_0__1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1574_ (.A(clknet_0__1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1574_));
 sky130_fd_sc_hd__clkbuf_4 clkload21 (.A(clknet_1_1__leaf__1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1589_ (.A(_1589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1589_ (.A(clknet_0__1589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1589_ (.A(clknet_0__1589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1589_));
 sky130_fd_sc_hd__clkbuf_4 clkload22 (.A(clknet_1_1__leaf__1589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1607_ (.A(_1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1607_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1607_ (.A(clknet_0__1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1607_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1607_ (.A(clknet_0__1607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1607_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload23 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net53 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net53));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net53 (.A(clknet_0_net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net53));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net53 (.A(clknet_0_net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net53));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_1_1__leaf_net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkinv_4 clkload25 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload26 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload27 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload28 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0527_ (.A(_0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0527_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0527_ (.A(clknet_0__0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0527_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0527_ (.A(clknet_0__0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0527_));
 sky130_fd_sc_hd__clkbuf_4 clkload29 (.A(clknet_1_1__leaf__0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0529_ (.A(_0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0529_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0529_ (.A(clknet_0__0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0529_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0529_ (.A(clknet_0__0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0529_));
 sky130_fd_sc_hd__clkinv_1 clkload30 (.A(clknet_1_0__leaf__0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0532_ (.A(_0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0532_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0532_ (.A(clknet_0__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0532_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0532_ (.A(clknet_0__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0532_));
 sky130_fd_sc_hd__clkinvlp_2 clkload31 (.A(clknet_1_1__leaf__0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1168_ (.A(_1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1168_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1168_ (.A(clknet_0__1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1168_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1168_ (.A(clknet_0__1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1168_));
 sky130_fd_sc_hd__clkbuf_4 clkload32 (.A(clknet_1_0__leaf__1168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out  (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkinv_4 clkload33 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload34 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1435_ (.A(_1435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1435_ (.A(clknet_0__1435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1435_ (.A(clknet_0__1435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1435_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload35 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload36 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1408_ (.A(_1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1408_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1408_ (.A(clknet_0__1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1408_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1408_ (.A(clknet_0__1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1408_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1699_ (.A(_1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1699_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1699_ (.A(clknet_0__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1699_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1699_ (.A(clknet_0__1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1699_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload37 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1759_ (.A(_1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1759_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1759_ (.A(clknet_0__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1759_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1759_ (.A(clknet_0__1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1759_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1749_ (.A(_1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1749_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1749_ (.A(clknet_0__1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1749_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1749_ (.A(clknet_0__1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1749_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0192_ (.A(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0192_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0192_ (.A(clknet_0__0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0192_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0192_ (.A(clknet_0__0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0192_));
 sky130_fd_sc_hd__clkinv_1 clkload38 (.A(clknet_1_1__leaf__0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1770_ (.A(_1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1770_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1770_ (.A(clknet_0__1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1770_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1770_ (.A(clknet_0__1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1770_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1238_ (.A(_1238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1238_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1238_ (.A(clknet_0__1238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1238_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1238_ (.A(clknet_0__1238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1238_));
 sky130_fd_sc_hd__clkbuf_4 clkload39 (.A(clknet_1_0__leaf__1238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out  (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_4 clkload40 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload41 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1393_ (.A(_1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1393_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1393_ (.A(clknet_0__1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1393_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1393_ (.A(clknet_0__1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1393_));
 sky130_fd_sc_hd__clkbuf_4 clkload42 (.A(clknet_1_0__leaf__1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1395_ (.A(_1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1395_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1395_ (.A(clknet_0__1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1395_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1395_ (.A(clknet_0__1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1395_));
 sky130_fd_sc_hd__clkbuf_4 clkload43 (.A(clknet_1_1__leaf__1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 clkload44 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload45 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1482_ (.A(_1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1482_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1482_ (.A(clknet_0__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1482_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1482_ (.A(clknet_0__1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1482_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload46 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1494_ (.A(_1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1494_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1494_ (.A(clknet_0__1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1494_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1494_ (.A(clknet_0__1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1494_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1470_ (.A(_1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1470_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1470_ (.A(clknet_0__1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1470_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1470_ (.A(clknet_0__1470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1470_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload47 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1336_ (.A(_1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1336_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1336_ (.A(clknet_0__1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1336_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1336_ (.A(clknet_0__1336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1336_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1359_ (.A(_1359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1359_ (.A(clknet_0__1359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1359_ (.A(clknet_0__1359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1256_ (.A(_1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1256_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1256_ (.A(clknet_0__1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1256_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1256_ (.A(clknet_0__1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1256_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload48 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net19 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net19 (.A(clknet_0_net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net19 (.A(clknet_0_net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net19));
 sky130_fd_sc_hd__clkinvlp_2 clkload49 (.A(clknet_1_1__leaf_net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1420_ (.A(_1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1420_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1420_ (.A(clknet_0__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1420_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1420_ (.A(clknet_0__1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1420_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net18 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net18));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net18 (.A(clknet_0_net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net18));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net18 (.A(clknet_0_net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net18));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1689_ (.A(_1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1689_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1689_ (.A(clknet_0__1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1689_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1689_ (.A(clknet_0__1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1689_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1712_ (.A(_1712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1712_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1712_ (.A(clknet_0__1712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1712_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1712_ (.A(clknet_0__1712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1712_));
 sky130_fd_sc_hd__inv_2 clkload50 (.A(clknet_1_1__leaf__1712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1729_ (.A(_1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1729_ (.A(clknet_0__1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1729_ (.A(clknet_0__1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1729_));
 sky130_fd_sc_hd__clkbuf_4 clkload51 (.A(clknet_1_0__leaf__1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0987_ (.A(_0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0987_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0987_ (.A(clknet_0__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0987_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0987_ (.A(clknet_0__0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0987_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload52 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net16 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net16 (.A(clknet_0_net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net16 (.A(clknet_0_net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net16));
 sky130_fd_sc_hd__clkbuf_4 clkload53 (.A(clknet_1_0__leaf_net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0534_ (.A(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0534_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0534_ (.A(clknet_0__0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0534_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0534_ (.A(clknet_0__0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0534_));
 sky130_fd_sc_hd__clkbuf_4 clkload54 (.A(clknet_1_1__leaf__0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0539_ (.A(_0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0539_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0539_ (.A(clknet_0__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0539_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0539_ (.A(clknet_0__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0539_));
 sky130_fd_sc_hd__bufinv_8 clkload55 (.A(clknet_1_1__leaf__0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0558_ (.A(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0558_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0558_ (.A(clknet_0__0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0558_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0558_ (.A(clknet_0__0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0558_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload56 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1188_ (.A(_1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1188_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1188_ (.A(clknet_0__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1188_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1188_ (.A(clknet_0__1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1188_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1648_ (.A(_1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1648_ (.A(clknet_0__1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1648_ (.A(clknet_0__1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1648_));
 sky130_fd_sc_hd__clkbuf_4 clkload57 (.A(clknet_1_0__leaf__1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1617_ (.A(_1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1617_ (.A(clknet_0__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1617_ (.A(clknet_0__1617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1627_ (.A(_1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1627_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1627_ (.A(clknet_0__1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1627_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1627_ (.A(clknet_0__1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1627_));
 sky130_fd_sc_hd__clkbuf_4 clkload58 (.A(clknet_1_1__leaf__1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1231_ (.A(_1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1231_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1231_ (.A(clknet_0__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1231_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1231_ (.A(clknet_0__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1231_));
 sky130_fd_sc_hd__bufinv_16 clkload59 (.A(clknet_1_0__leaf__1231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload60 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out  (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_4 clkload61 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload62 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload63 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0849_ (.A(_0849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0849_ (.A(clknet_0__0849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0849_ (.A(clknet_0__0849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0849_));
 sky130_fd_sc_hd__clkbuf_4 clkload64 (.A(clknet_1_0__leaf__0849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload65 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__bufinv_8 clkload66 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload67 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1054_ (.A(_1054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1054_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1054_ (.A(clknet_0__1054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1054_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1054_ (.A(clknet_0__1054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1054_));
 sky130_fd_sc_hd__clkbuf_4 clkload68 (.A(clknet_1_1__leaf__1054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload69 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload70 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload71 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0639_ (.A(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0639_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0639_ (.A(clknet_0__0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0639_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0639_ (.A(clknet_0__0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0639_));
 sky130_fd_sc_hd__bufinv_16 clkload72 (.A(clknet_1_1__leaf__0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload73 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0642_ (.A(_0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0642_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0642_ (.A(clknet_0__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0642_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0642_ (.A(clknet_0__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0642_));
 sky130_fd_sc_hd__bufinv_8 clkload74 (.A(clknet_1_0__leaf__0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0646_ (.A(_0646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0646_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0646_ (.A(clknet_0__0646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0646_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0646_ (.A(clknet_0__0646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0646_));
 sky130_fd_sc_hd__clkinv_2 clkload75 (.A(clknet_1_1__leaf__0646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload76 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0914_ (.A(_0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0914_ (.A(clknet_0__0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0914_ (.A(clknet_0__0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0914_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload77 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__inv_4 clkload78 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0524_ (.A(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0524_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0524_ (.A(clknet_0__0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0524_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0524_ (.A(clknet_0__0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0524_));
 sky130_fd_sc_hd__clkbuf_4 clkload79 (.A(clknet_1_0__leaf__0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0526_ (.A(_0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0526_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0526_ (.A(clknet_0__0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0526_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0526_ (.A(clknet_0__0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0526_));
 sky130_fd_sc_hd__clkbuf_4 clkload80 (.A(clknet_1_1__leaf__0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0528_ (.A(_0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0528_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0528_ (.A(clknet_0__0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0528_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0528_ (.A(clknet_0__0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0528_));
 sky130_fd_sc_hd__clkbuf_4 clkload81 (.A(clknet_1_0__leaf__0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0611_ (.A(_0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0611_ (.A(clknet_0__0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0611_ (.A(clknet_0__0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0611_));
 sky130_fd_sc_hd__clkbuf_4 clkload82 (.A(clknet_1_1__leaf__0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1072_ (.A(_1072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1072_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1072_ (.A(clknet_0__1072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1072_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1072_ (.A(clknet_0__1072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1072_));
 sky130_fd_sc_hd__clkbuf_4 clkload83 (.A(clknet_1_1__leaf__1072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1077_ (.A(_1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1077_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1077_ (.A(clknet_0__1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1077_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1077_ (.A(clknet_0__1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1077_));
 sky130_fd_sc_hd__bufinv_8 clkload84 (.A(clknet_1_0__leaf__1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__bufinv_8 clkload85 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload86 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload87 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0598_ (.A(_0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0598_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0598_ (.A(clknet_0__0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0598_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0598_ (.A(clknet_0__0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0598_));
 sky130_fd_sc_hd__clkbuf_4 clkload88 (.A(clknet_1_1__leaf__0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0600_ (.A(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0600_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0600_ (.A(clknet_0__0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0600_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0600_ (.A(clknet_0__0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0600_));
 sky130_fd_sc_hd__clkbuf_4 clkload89 (.A(clknet_1_1__leaf__0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0771_ (.A(_0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0771_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0771_ (.A(clknet_0__0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0771_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0771_ (.A(clknet_0__0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0771_));
 sky130_fd_sc_hd__clkbuf_4 clkload90 (.A(clknet_1_0__leaf__0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0791_ (.A(_0791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0791_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0791_ (.A(clknet_0__0791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0791_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0791_ (.A(clknet_0__0791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0791_));
 sky130_fd_sc_hd__clkbuf_4 clkload91 (.A(clknet_1_0__leaf__0791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0794_ (.A(_0794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0794_ (.A(clknet_0__0794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0794_ (.A(clknet_0__0794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0794_));
 sky130_fd_sc_hd__clkbuf_4 clkload92 (.A(clknet_1_1__leaf__0794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0805_ (.A(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0805_ (.A(clknet_0__0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0805_ (.A(clknet_0__0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0805_));
 sky130_fd_sc_hd__clkbuf_4 clkload93 (.A(clknet_1_0__leaf__0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload94 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1346_ (.A(_1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1346_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1346_ (.A(clknet_0__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1346_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1346_ (.A(clknet_0__1346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1346_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1280_ (.A(_1280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1280_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1280_ (.A(clknet_0__1280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1280_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1280_ (.A(clknet_0__1280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1280_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1266_ (.A(_1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1266_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1266_ (.A(clknet_0__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1266_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1266_ (.A(clknet_0__1266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1266_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0938_ (.A(_0938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0938_ (.A(clknet_0__0938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0938_ (.A(clknet_0__0938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0924_ (.A(_0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0924_ (.A(clknet_0__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0924_ (.A(clknet_0__0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0879_ (.A(_0879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0879_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0879_ (.A(clknet_0__0879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0879_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0879_ (.A(clknet_0__0879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0879_));
 sky130_fd_sc_hd__clkbuf_4 clkload95 (.A(clknet_1_1__leaf__0879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0881_ (.A(_0881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0881_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0881_ (.A(clknet_0__0881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0881_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0881_ (.A(clknet_0__0881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0881_));
 sky130_fd_sc_hd__clkbuf_4 clkload96 (.A(clknet_1_0__leaf__0881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0883_ (.A(_0883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0883_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0883_ (.A(clknet_0__0883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0883_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0883_ (.A(clknet_0__0883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0883_));
 sky130_fd_sc_hd__clkinv_1 clkload97 (.A(clknet_1_1__leaf__0883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1091_ (.A(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1091_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1091_ (.A(clknet_0__1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1091_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1091_ (.A(clknet_0__1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1091_));
 sky130_fd_sc_hd__clkbuf_4 clkload98 (.A(clknet_1_0__leaf__1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload99 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0744_ (.A(_0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0744_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0744_ (.A(clknet_0__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0744_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0744_ (.A(clknet_0__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0744_));
 sky130_fd_sc_hd__inv_2 clkload100 (.A(clknet_1_0__leaf__0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload101 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0742_ (.A(_0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0742_ (.A(clknet_0__0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0742_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0742_ (.A(clknet_0__0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0742_));
 sky130_fd_sc_hd__clkinvlp_2 clkload102 (.A(clknet_1_1__leaf__0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload103 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0553_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0553_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0553_ (.A(clknet_0__0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0553_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0553_ (.A(clknet_0__0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0553_));
 sky130_fd_sc_hd__clkbuf_4 clkload104 (.A(clknet_1_0__leaf__0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0554_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0554_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0554_ (.A(clknet_0__0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0554_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0554_ (.A(clknet_0__0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0554_));
 sky130_fd_sc_hd__clkbuf_4 clkload105 (.A(clknet_1_0__leaf__0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0785_ (.A(_0785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0785_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0785_ (.A(clknet_0__0785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0785_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0785_ (.A(clknet_0__0785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0785_));
 sky130_fd_sc_hd__clkbuf_4 clkload106 (.A(clknet_1_1__leaf__0785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0829_ (.A(_0829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0829_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0829_ (.A(clknet_0__0829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0829_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0829_ (.A(clknet_0__0829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0829_));
 sky130_fd_sc_hd__clkbuf_4 clkload107 (.A(clknet_1_1__leaf__0829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload108 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0831_ (.A(_0831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0831_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0831_ (.A(clknet_0__0831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0831_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0831_ (.A(clknet_0__0831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0831_));
 sky130_fd_sc_hd__clkbuf_4 clkload109 (.A(clknet_1_1__leaf__0831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload110 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1049_ (.A(_1049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1049_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1049_ (.A(clknet_0__1049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1049_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1049_ (.A(clknet_0__1049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1049_));
 sky130_fd_sc_hd__clkbuf_4 clkload111 (.A(clknet_1_1__leaf__1049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1061_ (.A(_1061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1061_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1061_ (.A(clknet_0__1061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1061_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1061_ (.A(clknet_0__1061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1061_));
 sky130_fd_sc_hd__bufinv_8 clkload112 (.A(clknet_1_1__leaf__1061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out  (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_8 clkload113 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload114 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0223_ (.A(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0223_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0223_ (.A(clknet_0__0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0223_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0223_ (.A(clknet_0__0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0223_));
 sky130_fd_sc_hd__clkbuf_4 clkload115 (.A(clknet_1_1__leaf__0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0789_ (.A(_0789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0789_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0789_ (.A(clknet_0__0789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0789_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0789_ (.A(clknet_0__0789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0789_));
 sky130_fd_sc_hd__clkbuf_2 clkload116 (.A(clknet_1_0__leaf__0789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0790_ (.A(_0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0790_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0790_ (.A(clknet_0__0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0790_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0790_ (.A(clknet_0__0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0790_));
 sky130_fd_sc_hd__inv_2 clkload117 (.A(clknet_1_1__leaf__0790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkinv_1 clkload118 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0895_ (.A(_0895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0895_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0895_ (.A(clknet_0__0895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0895_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0895_ (.A(clknet_0__0895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0895_));
 sky130_fd_sc_hd__clkbuf_4 clkload119 (.A(clknet_1_0__leaf__0895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0897_ (.A(_0897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0897_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0897_ (.A(clknet_0__0897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0897_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0897_ (.A(clknet_0__0897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0897_));
 sky130_fd_sc_hd__clkbuf_4 clkload120 (.A(clknet_1_1__leaf__0897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkinvlp_4 clkload121 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload122 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0977_ (.A(_0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0977_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0977_ (.A(clknet_0__0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0977_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0977_ (.A(clknet_0__0977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0977_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1000_ (.A(_1000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1000_ (.A(clknet_0__1000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1000_ (.A(clknet_0__1000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1314_ (.A(_1314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1314_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1314_ (.A(clknet_0__1314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1314_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1314_ (.A(clknet_0__1314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1314_));
 sky130_fd_sc_hd__clkbuf_4 clkload123 (.A(clknet_1_0__leaf__1314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1316_ (.A(_1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1316_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1316_ (.A(clknet_0__1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1316_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1316_ (.A(clknet_0__1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1316_));
 sky130_fd_sc_hd__clkbuf_4 clkload124 (.A(clknet_1_0__leaf__1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload125 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out  (.A(\dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkbuf_4 clkload126 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_left_ipin_1.INVTX1_1_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0846_ (.A(_0846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0846_ (.A(clknet_0__0846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0846_ (.A(clknet_0__0846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0846_));
 sky130_fd_sc_hd__clkbuf_4 clkload127 (.A(clknet_1_0__leaf__0846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload128 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0723_ (.A(_0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0723_ (.A(clknet_0__0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0723_ (.A(clknet_0__0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0723_));
 sky130_fd_sc_hd__clkbuf_4 clkload129 (.A(clknet_1_0__leaf__0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net33 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net33));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net33 (.A(clknet_0_net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net33));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net33 (.A(clknet_0_net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net33));
 sky130_fd_sc_hd__clkbuf_8 clkload130 (.A(clknet_1_1__leaf_net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1033_ (.A(_1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1033_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1033_ (.A(clknet_0__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1033_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1033_ (.A(clknet_0__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1033_));
 sky130_fd_sc_hd__bufinv_16 clkload131 (.A(clknet_1_1__leaf__1033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1035_ (.A(_1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1035_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1035_ (.A(clknet_0__1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1035_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1035_ (.A(clknet_0__1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1035_));
 sky130_fd_sc_hd__clkbuf_4 clkload132 (.A(clknet_1_1__leaf__1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out  (.A(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload133 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload134 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0445_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0445_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0445_ (.A(clknet_0__0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0445_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0445_ (.A(clknet_0__0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0445_));
 sky130_fd_sc_hd__clkbuf_4 clkload135 (.A(clknet_1_0__leaf__0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0426_ (.A(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0426_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0426_ (.A(clknet_0__0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0426_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0426_ (.A(clknet_0__0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0426_));
 sky130_fd_sc_hd__clkinv_1 clkload136 (.A(clknet_1_1__leaf__0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0378_ (.A(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0378_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0378_ (.A(clknet_0__0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0378_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0378_ (.A(clknet_0__0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0378_));
 sky130_fd_sc_hd__clkbuf_4 clkload137 (.A(clknet_1_0__leaf__0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload138 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0359_ (.A(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0359_ (.A(clknet_0__0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0359_ (.A(clknet_0__0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0359_));
 sky130_fd_sc_hd__clkbuf_4 clkload139 (.A(clknet_1_1__leaf__0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0345_ (.A(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0345_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0345_ (.A(clknet_0__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0345_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0345_ (.A(clknet_0__0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0345_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0333_ (.A(_0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0333_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0333_ (.A(clknet_0__0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0333_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0333_ (.A(clknet_0__0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0333_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0292_ (.A(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0292_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0292_ (.A(clknet_0__0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0292_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0292_ (.A(clknet_0__0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0292_));
 sky130_fd_sc_hd__clkbuf_4 clkload140 (.A(clknet_1_1__leaf__0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0266_ (.A(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0266_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0266_ (.A(clknet_0__0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0266_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0266_ (.A(clknet_0__0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0266_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0412_ (.A(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0412_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0412_ (.A(clknet_0__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0412_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0412_ (.A(clknet_0__0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0412_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0511_ (.A(_0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0511_ (.A(clknet_0__0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0511_ (.A(clknet_0__0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0511_));
 sky130_fd_sc_hd__clkbuf_4 clkload141 (.A(clknet_1_1__leaf__0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload142 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload143 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0311_ (.A(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0311_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0311_ (.A(clknet_0__0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0311_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0311_ (.A(clknet_0__0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0311_));
 sky130_fd_sc_hd__clkbuf_4 clkload144 (.A(clknet_1_1__leaf__0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0479_ (.A(_0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0479_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0479_ (.A(clknet_0__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0479_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0479_ (.A(clknet_0__0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0479_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0493_ (.A(_0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0493_ (.A(clknet_0__0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0493_ (.A(clknet_0__0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0493_));
 sky130_fd_sc_hd__clkinv_2 clkload145 (.A(clknet_1_1__leaf__0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0467_ (.A(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0467_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0467_ (.A(clknet_0__0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0467_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0467_ (.A(clknet_0__0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0467_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload146 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0868_ (.A(_0868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0868_ (.A(clknet_0__0868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0868_ (.A(clknet_0__0868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0868_));
 sky130_fd_sc_hd__bufinv_8 clkload147 (.A(clknet_1_1__leaf__0868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__bufinv_16 clkload148 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_0.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload149 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0530_ (.A(_0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0530_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0530_ (.A(clknet_0__0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0530_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0530_ (.A(clknet_0__0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0530_));
 sky130_fd_sc_hd__clkinv_1 clkload150 (.A(clknet_1_0__leaf__0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0531_ (.A(_0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0531_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0531_ (.A(clknet_0__0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0531_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0531_ (.A(clknet_0__0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0531_));
 sky130_fd_sc_hd__clkbuf_4 clkload151 (.A(clknet_1_0__leaf__0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0623_ (.A(_0623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0623_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0623_ (.A(clknet_0__0623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0623_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0623_ (.A(clknet_0__0623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0623_));
 sky130_fd_sc_hd__clkbuf_4 clkload152 (.A(clknet_1_0__leaf__0623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0624_ (.A(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0624_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0624_ (.A(clknet_0__0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0624_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0624_ (.A(clknet_0__0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0624_));
 sky130_fd_sc_hd__clkbuf_8 clkload153 (.A(clknet_1_1__leaf__0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0860_ (.A(_0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0860_ (.A(clknet_0__0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0860_ (.A(clknet_0__0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0860_));
 sky130_fd_sc_hd__clkinv_2 clkload154 (.A(clknet_1_1__leaf__0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload155 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0633_ (.A(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0633_ (.A(clknet_0__0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0633_ (.A(clknet_0__0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0633_));
 sky130_fd_sc_hd__clkbuf_4 clkload156 (.A(clknet_1_1__leaf__0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0634_ (.A(_0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0634_ (.A(clknet_0__0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0634_ (.A(clknet_0__0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0634_));
 sky130_fd_sc_hd__clkbuf_4 clkload157 (.A(clknet_1_1__leaf__0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload158 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload159 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0226_ (.A(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0226_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0226_ (.A(clknet_0__0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0226_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0226_ (.A(clknet_0__0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0226_));
 sky130_fd_sc_hd__clkinv_2 clkload160 (.A(clknet_1_1__leaf__0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0245_ (.A(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0245_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0245_ (.A(clknet_0__0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0245_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0245_ (.A(clknet_0__0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0245_));
 sky130_fd_sc_hd__clkinv_2 clkload161 (.A(clknet_1_1__leaf__0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0249_ (.A(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0249_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0249_ (.A(clknet_0__0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0249_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0249_ (.A(clknet_0__0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0249_));
 sky130_fd_sc_hd__clkbuf_4 clkload162 (.A(clknet_1_1__leaf__0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0252_ (.A(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0252_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0252_ (.A(clknet_0__0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0252_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0252_ (.A(clknet_0__0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0252_));
 sky130_fd_sc_hd__clkbuf_4 clkload163 (.A(clknet_1_1__leaf__0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0619_ (.A(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0619_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0619_ (.A(clknet_0__0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0619_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0619_ (.A(clknet_0__0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0619_));
 sky130_fd_sc_hd__clkbuf_4 clkload164 (.A(clknet_1_0__leaf__0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0622_ (.A(_0622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0622_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0622_ (.A(clknet_0__0622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0622_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0622_ (.A(clknet_0__0622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0622_));
 sky130_fd_sc_hd__clkbuf_4 clkload165 (.A(clknet_1_1__leaf__0622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0621_ (.A(_0621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0621_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0621_ (.A(clknet_0__0621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0621_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0621_ (.A(clknet_0__0621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0621_));
 sky130_fd_sc_hd__clkbuf_4 clkload166 (.A(clknet_1_0__leaf__0621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkinv_2 clkload167 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_top_ipin_2.INVTX1_5_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net35 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net35 (.A(clknet_0_net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net35));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net35 (.A(clknet_0_net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net35));
 sky130_fd_sc_hd__clkinvlp_2 clkload168 (.A(clknet_1_0__leaf_net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload169 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0246_ (.A(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0246_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0246_ (.A(clknet_0__0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0246_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0246_ (.A(clknet_0__0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0246_));
 sky130_fd_sc_hd__clkinv_2 clkload170 (.A(clknet_1_1__leaf__0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0248_ (.A(_0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0248_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0248_ (.A(clknet_0__0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0248_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0248_ (.A(clknet_0__0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0248_));
 sky130_fd_sc_hd__clkbuf_4 clkload171 (.A(clknet_1_1__leaf__0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0602_ (.A(_0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0602_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0602_ (.A(clknet_0__0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0602_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0602_ (.A(clknet_0__0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0602_));
 sky130_fd_sc_hd__clkbuf_4 clkload172 (.A(clknet_1_1__leaf__0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0613_ (.A(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0613_ (.A(clknet_0__0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0613_ (.A(clknet_0__0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0613_));
 sky130_fd_sc_hd__clkbuf_4 clkload173 (.A(clknet_1_1__leaf__0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0603_ (.A(_0603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0603_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0603_ (.A(clknet_0__0603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0603_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0603_ (.A(clknet_0__0603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0603_));
 sky130_fd_sc_hd__clkbuf_4 clkload174 (.A(clknet_1_1__leaf__0603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1102_ (.A(_1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1102_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1102_ (.A(clknet_0__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1102_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1102_ (.A(clknet_0__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1102_));
 sky130_fd_sc_hd__clkinv_4 clkload175 (.A(clknet_1_0__leaf__1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net22 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net22 (.A(clknet_0_net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net22));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net22 (.A(clknet_0_net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net22));
 sky130_fd_sc_hd__clkbuf_8 clkload176 (.A(clknet_1_1__leaf_net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload177 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0247_ (.A(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0247_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0247_ (.A(clknet_0__0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0247_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0247_ (.A(clknet_0__0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0247_));
 sky130_fd_sc_hd__clkinvlp_2 clkload178 (.A(clknet_1_1__leaf__0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload179 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1095_ (.A(_1095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__1095_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1095_ (.A(clknet_0__1095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__1095_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1095_ (.A(clknet_0__1095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__1095_));
 sky130_fd_sc_hd__clkbuf_4 clkload180 (.A(clknet_1_0__leaf__1095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out  (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__clkinvlp_4 clkload181 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload182 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0792_ (.A(_0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0792_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0792_ (.A(clknet_0__0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0792_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0792_ (.A(clknet_0__0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0792_));
 sky130_fd_sc_hd__clkbuf_4 clkload183 (.A(clknet_1_0__leaf__0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0793_ (.A(_0793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0793_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0793_ (.A(clknet_0__0793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0793_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0793_ (.A(clknet_0__0793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0793_));
 sky130_fd_sc_hd__bufinv_8 clkload184 (.A(clknet_1_1__leaf__0793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload185 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload186 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0681_ (.A(_0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0681_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0681_ (.A(clknet_0__0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0681_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0681_ (.A(clknet_0__0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0681_));
 sky130_fd_sc_hd__clkinv_1 clkload187 (.A(clknet_1_1__leaf__0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0730_ (.A(_0730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0730_ (.A(clknet_0__0730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0730_ (.A(clknet_0__0730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0730_));
 sky130_fd_sc_hd__clkinv_2 clkload188 (.A(clknet_1_1__leaf__0730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload189 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload190 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload191 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0250_ (.A(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0250_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0250_ (.A(clknet_0__0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0250_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0250_ (.A(clknet_0__0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0250_));
 sky130_fd_sc_hd__clkbuf_4 clkload192 (.A(clknet_1_1__leaf__0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0251_ (.A(_0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0251_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0251_ (.A(clknet_0__0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0251_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0251_ (.A(clknet_0__0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0251_));
 sky130_fd_sc_hd__clkbuf_4 clkload193 (.A(clknet_1_1__leaf__0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\dut_0.U0_formal_verification.cbx_1__2_.mem_bottom_ipin_3.DFF_2_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\dut_0.U0_formal_verification.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinvlp_2 clkload194 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__1_.mux_top_ipin_2.INVTX1_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0236_ (.A(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0236_ (.A(clknet_0__0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0236_ (.A(clknet_0__0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0236_));
 sky130_fd_sc_hd__bufinv_8 clkload195 (.A(clknet_1_0__leaf__0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload196 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0738_ (.A(_0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0738_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0738_ (.A(clknet_0__0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0738_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0738_ (.A(clknet_0__0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0738_));
 sky130_fd_sc_hd__clkbuf_4 clkload197 (.A(clknet_1_0__leaf__0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\dut_0.U0_formal_verification.cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_6 clkload198 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.INVTX1_2_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0811_ (.A(_0811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0811_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0811_ (.A(clknet_0__0811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0811_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0811_ (.A(clknet_0__0811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0811_));
 sky130_fd_sc_hd__clkinvlp_2 clkload199 (.A(clknet_1_1__leaf__0811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0816_ (.A(_0816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0816_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0816_ (.A(clknet_0__0816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0816_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0816_ (.A(clknet_0__0816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0816_));
 sky130_fd_sc_hd__inv_2 clkload200 (.A(clknet_1_1__leaf__0816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0889_ (.A(_0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0889_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0889_ (.A(clknet_0__0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0889_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0889_ (.A(clknet_0__0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0889_));
 sky130_fd_sc_hd__bufinv_8 clkload201 (.A(clknet_1_1__leaf__0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net28 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net28));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net28 (.A(clknet_0_net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net28));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net28 (.A(clknet_0_net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net28));
 sky130_fd_sc_hd__clkinvlp_2 clkload202 (.A(clknet_1_1__leaf_net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net27 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net27 (.A(clknet_0_net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net27 (.A(clknet_0_net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net27));
 sky130_fd_sc_hd__clkinv_1 clkload203 (.A(clknet_1_1__leaf_net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0813_ (.A(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0813_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0813_ (.A(clknet_0__0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0813_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0813_ (.A(clknet_0__0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0813_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload204 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload205 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload206 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0812_ (.A(_0812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0812_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0812_ (.A(clknet_0__0812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0812_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0812_ (.A(clknet_0__0812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0812_));
 sky130_fd_sc_hd__clkbuf_4 clkload207 (.A(clknet_1_0__leaf__0812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload208 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload209 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0592_ (.A(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0592_ (.A(clknet_0__0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0592_ (.A(clknet_0__0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0592_));
 sky130_fd_sc_hd__clkbuf_4 clkload210 (.A(clknet_1_0__leaf__0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0594_ (.A(_0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0594_ (.A(clknet_0__0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0594_ (.A(clknet_0__0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0594_));
 sky130_fd_sc_hd__clkbuf_4 clkload211 (.A(clknet_1_1__leaf__0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0597_ (.A(_0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0597_ (.A(clknet_0__0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0597_ (.A(clknet_0__0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0597_));
 sky130_fd_sc_hd__clkbuf_4 clkload212 (.A(clknet_1_1__leaf__0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0599_ (.A(_0599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0599_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0599_ (.A(clknet_0__0599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0599_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0599_ (.A(clknet_0__0599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0599_));
 sky130_fd_sc_hd__clkbuf_4 clkload213 (.A(clknet_1_0__leaf__0599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload214 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0570_ (.A(_0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0570_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0570_ (.A(clknet_0__0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0570_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0570_ (.A(clknet_0__0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0570_));
 sky130_fd_sc_hd__clkbuf_4 clkload215 (.A(clknet_1_0__leaf__0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0588_ (.A(_0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0588_ (.A(clknet_0__0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0588_ (.A(clknet_0__0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0588_));
 sky130_fd_sc_hd__clkbuf_4 clkload216 (.A(clknet_1_0__leaf__0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0591_ (.A(_0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0591_ (.A(clknet_0__0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0591_ (.A(clknet_0__0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0591_));
 sky130_fd_sc_hd__clkbuf_4 clkload217 (.A(clknet_1_0__leaf__0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0593_ (.A(_0593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0593_ (.A(clknet_0__0593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0593_ (.A(clknet_0__0593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0593_));
 sky130_fd_sc_hd__bufinv_8 clkload218 (.A(clknet_1_1__leaf__0593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload219 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0650_ (.A(_0650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0650_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0650_ (.A(clknet_0__0650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0650_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0650_ (.A(clknet_0__0650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0650_));
 sky130_fd_sc_hd__clkbuf_4 clkload220 (.A(clknet_1_1__leaf__0650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload221 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload222 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0775_ (.A(_0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0775_ (.A(clknet_0__0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0775_ (.A(clknet_0__0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0775_));
 sky130_fd_sc_hd__clkbuf_4 clkload223 (.A(clknet_1_0__leaf__0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0535_ (.A(_0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0535_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0535_ (.A(clknet_0__0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0535_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0535_ (.A(clknet_0__0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0535_));
 sky130_fd_sc_hd__clkbuf_4 clkload224 (.A(clknet_1_0__leaf__0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0542_ (.A(_0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0542_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0542_ (.A(clknet_0__0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0542_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0542_ (.A(clknet_0__0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0542_));
 sky130_fd_sc_hd__clkbuf_4 clkload225 (.A(clknet_1_0__leaf__0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0545_ (.A(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0545_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0545_ (.A(clknet_0__0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0545_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0545_ (.A(clknet_0__0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0545_));
 sky130_fd_sc_hd__clkbuf_4 clkload226 (.A(clknet_1_1__leaf__0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0548_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0548_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0548_ (.A(clknet_0__0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0548_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0548_ (.A(clknet_0__0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0548_));
 sky130_fd_sc_hd__clkbuf_4 clkload227 (.A(clknet_1_0__leaf__0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0551_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0551_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0551_ (.A(clknet_0__0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0551_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0551_ (.A(clknet_0__0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0551_));
 sky130_fd_sc_hd__clkbuf_4 clkload228 (.A(clknet_1_0__leaf__0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0555_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0555_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0555_ (.A(clknet_0__0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0555_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0555_ (.A(clknet_0__0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0555_));
 sky130_fd_sc_hd__clkbuf_4 clkload229 (.A(clknet_1_0__leaf__0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0550_ (.A(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0550_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0550_ (.A(clknet_0__0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0550_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0550_ (.A(clknet_0__0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0550_));
 sky130_fd_sc_hd__clkbuf_4 clkload230 (.A(clknet_1_0__leaf__0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0702_ (.A(_0702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0702_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0702_ (.A(clknet_0__0702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0702_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0702_ (.A(clknet_0__0702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0702_));
 sky130_fd_sc_hd__bufinv_8 clkload231 (.A(clknet_1_0__leaf__0702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0704_ (.A(_0704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0704_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0704_ (.A(clknet_0__0704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0704_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0704_ (.A(clknet_0__0704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0704_));
 sky130_fd_sc_hd__clkbuf_4 clkload232 (.A(clknet_1_0__leaf__0704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload233 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload234 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0665_ (.A(_0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0665_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0665_ (.A(clknet_0__0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0665_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0665_ (.A(clknet_0__0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0665_));
 sky130_fd_sc_hd__clkinv_1 clkload235 (.A(clknet_1_1__leaf__0665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload236 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__2_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0667_ (.A(_0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0667_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0667_ (.A(clknet_0__0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0667_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0667_ (.A(clknet_0__0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0667_));
 sky130_fd_sc_hd__clkinv_1 clkload237 (.A(clknet_1_0__leaf__0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0669_ (.A(_0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0669_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0669_ (.A(clknet_0__0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0669_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0669_ (.A(clknet_0__0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0669_));
 sky130_fd_sc_hd__bufinv_8 clkload238 (.A(clknet_1_1__leaf__0669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0795_ (.A(_0795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0795_ (.A(clknet_0__0795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0795_ (.A(clknet_0__0795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0795_));
 sky130_fd_sc_hd__clkbuf_4 clkload239 (.A(clknet_1_1__leaf__0795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0796_ (.A(_0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0796_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0796_ (.A(clknet_0__0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0796_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0796_ (.A(clknet_0__0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0796_));
 sky130_fd_sc_hd__clkinv_1 clkload240 (.A(clknet_1_1__leaf__0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0671_ (.A(_0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0671_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0671_ (.A(clknet_0__0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0671_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0671_ (.A(clknet_0__0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0671_));
 sky130_fd_sc_hd__bufinv_8 clkload241 (.A(clknet_1_1__leaf__0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0675_ (.A(_0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0675_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0675_ (.A(clknet_0__0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0675_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0675_ (.A(clknet_0__0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0675_));
 sky130_fd_sc_hd__clkbuf_4 clkload242 (.A(clknet_1_1__leaf__0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload243 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0668_ (.A(_0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0668_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0668_ (.A(clknet_0__0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0668_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0668_ (.A(clknet_0__0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0668_));
 sky130_fd_sc_hd__inv_2 clkload244 (.A(clknet_1_1__leaf__0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_2 clkload245 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload246 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0567_ (.A(_0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0567_ (.A(clknet_0__0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0567_ (.A(clknet_0__0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0567_));
 sky130_fd_sc_hd__clkbuf_4 clkload247 (.A(clknet_1_0__leaf__0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0569_ (.A(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0569_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0569_ (.A(clknet_0__0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0569_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0569_ (.A(clknet_0__0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0569_));
 sky130_fd_sc_hd__clkbuf_4 clkload248 (.A(clknet_1_0__leaf__0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0572_ (.A(_0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0572_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0572_ (.A(clknet_0__0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0572_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0572_ (.A(clknet_0__0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0572_));
 sky130_fd_sc_hd__inv_1 clkload249 (.A(clknet_1_1__leaf__0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0574_ (.A(_0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0574_ (.A(clknet_0__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0574_ (.A(clknet_0__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0574_));
 sky130_fd_sc_hd__inv_6 clkload250 (.A(clknet_1_1__leaf__0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__inv_4 clkload251 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload252 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0571_ (.A(_0571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0571_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0571_ (.A(clknet_0__0571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0571_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0571_ (.A(clknet_0__0571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0571_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload253 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0546_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0546_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0546_ (.A(clknet_0__0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0546_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0546_ (.A(clknet_0__0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0546_));
 sky130_fd_sc_hd__clkbuf_4 clkload254 (.A(clknet_1_1__leaf__0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0547_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0547_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0547_ (.A(clknet_0__0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0547_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0547_ (.A(clknet_0__0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0547_));
 sky130_fd_sc_hd__clkinv_1 clkload255 (.A(clknet_1_0__leaf__0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0568_ (.A(_0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0568_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0568_ (.A(clknet_0__0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0568_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0568_ (.A(clknet_0__0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0568_));
 sky130_fd_sc_hd__clkbuf_4 clkload256 (.A(clknet_1_1__leaf__0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload257 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0230_ (.A(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0230_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0230_ (.A(clknet_0__0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0230_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0230_ (.A(clknet_0__0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0230_));
 sky130_fd_sc_hd__clkbuf_4 clkload258 (.A(clknet_1_0__leaf__0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0255_ (.A(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0255_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0255_ (.A(clknet_0__0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0255_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0255_ (.A(clknet_0__0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0255_));
 sky130_fd_sc_hd__clkbuf_4 clkload259 (.A(clknet_1_0__leaf__0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0523_ (.A(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0523_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0523_ (.A(clknet_0__0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0523_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0523_ (.A(clknet_0__0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0523_));
 sky130_fd_sc_hd__clkbuf_4 clkload260 (.A(clknet_1_0__leaf__0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0525_ (.A(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0525_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0525_ (.A(clknet_0__0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0525_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0525_ (.A(clknet_0__0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0525_));
 sky130_fd_sc_hd__clkbuf_4 clkload261 (.A(clknet_1_1__leaf__0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload262 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload263 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0543_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0543_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0543_ (.A(clknet_0__0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0543_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0543_ (.A(clknet_0__0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0543_));
 sky130_fd_sc_hd__clkbuf_4 clkload264 (.A(clknet_1_0__leaf__0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0544_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0544_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0544_ (.A(clknet_0__0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0544_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0544_ (.A(clknet_0__0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0544_));
 sky130_fd_sc_hd__clkbuf_4 clkload265 (.A(clknet_1_0__leaf__0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0688_ (.A(_0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0688_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0688_ (.A(clknet_0__0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0688_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0688_ (.A(clknet_0__0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0688_));
 sky130_fd_sc_hd__clkbuf_4 clkload266 (.A(clknet_1_1__leaf__0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload267 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload268 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0764_ (.A(_0764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0764_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0764_ (.A(clknet_0__0764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0764_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0764_ (.A(clknet_0__0764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0764_));
 sky130_fd_sc_hd__clkbuf_4 clkload269 (.A(clknet_1_1__leaf__0764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0766_ (.A(_0766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0766_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0766_ (.A(clknet_0__0766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0766_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0766_ (.A(clknet_0__0766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0766_));
 sky130_fd_sc_hd__clkbuf_4 clkload270 (.A(clknet_1_1__leaf__0766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload271 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0578_ (.A(_0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0578_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0578_ (.A(clknet_0__0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0578_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0578_ (.A(clknet_0__0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0578_));
 sky130_fd_sc_hd__clkinv_1 clkload272 (.A(clknet_1_1__leaf__0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0677_ (.A(_0677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0677_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0677_ (.A(clknet_0__0677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0677_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0677_ (.A(clknet_0__0677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0677_));
 sky130_fd_sc_hd__clkinv_2 clkload273 (.A(clknet_1_0__leaf__0677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0700_ (.A(_0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0700_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0700_ (.A(clknet_0__0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0700_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0700_ (.A(clknet_0__0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0700_));
 sky130_fd_sc_hd__bufinv_8 clkload274 (.A(clknet_1_1__leaf__0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload275 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_1__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0679_ (.A(_0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0679_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0679_ (.A(clknet_0__0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0679_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0679_ (.A(clknet_0__0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0679_));
 sky130_fd_sc_hd__clkinv_1 clkload276 (.A(clknet_1_0__leaf__0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0714_ (.A(_0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0714_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0714_ (.A(clknet_0__0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0714_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0714_ (.A(clknet_0__0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0714_));
 sky130_fd_sc_hd__clkbuf_4 clkload277 (.A(clknet_1_1__leaf__0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0718_ (.A(_0718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0718_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0718_ (.A(clknet_0__0718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0718_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0718_ (.A(clknet_0__0718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0718_));
 sky130_fd_sc_hd__clkbuf_4 clkload278 (.A(clknet_1_1__leaf__0718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload279 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload280 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__2.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload281 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload282 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0256_ (.A(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0256_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0256_ (.A(clknet_0__0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0256_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0256_ (.A(clknet_0__0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0256_));
 sky130_fd_sc_hd__clkbuf_4 clkload283 (.A(clknet_1_0__leaf__0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0257_ (.A(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0257_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0257_ (.A(clknet_0__0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0257_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0257_ (.A(clknet_0__0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0257_));
 sky130_fd_sc_hd__clkinv_1 clkload284 (.A(clknet_1_0__leaf__0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0259_ (.A(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0259_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0259_ (.A(clknet_0__0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0259_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0259_ (.A(clknet_0__0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0259_));
 sky130_fd_sc_hd__inv_2 clkload285 (.A(clknet_1_1__leaf__0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0261_ (.A(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0261_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0261_ (.A(clknet_0__0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0261_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0261_ (.A(clknet_0__0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0261_));
 sky130_fd_sc_hd__clkbuf_8 clkload286 (.A(clknet_1_0__leaf__0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload287 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0653_ (.A(_0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0653_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0653_ (.A(clknet_0__0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0653_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0653_ (.A(clknet_0__0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0653_));
 sky130_fd_sc_hd__clkbuf_4 clkload288 (.A(clknet_1_0__leaf__0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0655_ (.A(_0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0655_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0655_ (.A(clknet_0__0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0655_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0655_ (.A(clknet_0__0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0655_));
 sky130_fd_sc_hd__clkbuf_4 clkload289 (.A(clknet_1_1__leaf__0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload290 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload291 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0626_ (.A(_0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0626_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0626_ (.A(clknet_0__0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0626_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0626_ (.A(clknet_0__0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0626_));
 sky130_fd_sc_hd__clkinv_1 clkload292 (.A(clknet_1_1__leaf__0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0628_ (.A(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0628_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0628_ (.A(clknet_0__0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0628_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0628_ (.A(clknet_0__0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0628_));
 sky130_fd_sc_hd__clkbuf_4 clkload293 (.A(clknet_1_1__leaf__0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_8 clkload294 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__2_.mux_top_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload295 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0648_ (.A(_0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0648_ (.A(clknet_0__0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0648_ (.A(clknet_0__0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0648_));
 sky130_fd_sc_hd__clkbuf_4 clkload296 (.A(clknet_1_0__leaf__0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload297 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0253_ (.A(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0253_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0253_ (.A(clknet_0__0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0253_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0253_ (.A(clknet_0__0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0253_));
 sky130_fd_sc_hd__clkbuf_4 clkload298 (.A(clknet_1_1__leaf__0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0254_ (.A(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0254_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0254_ (.A(clknet_0__0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0254_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0254_ (.A(clknet_0__0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0254_));
 sky130_fd_sc_hd__clkbuf_4 clkload299 (.A(clknet_1_0__leaf__0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload300 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload301 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0661_ (.A(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0661_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0661_ (.A(clknet_0__0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0661_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0661_ (.A(clknet_0__0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0661_));
 sky130_fd_sc_hd__clkbuf_4 clkload302 (.A(clknet_1_0__leaf__0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0899_ (.A(_0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0899_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0899_ (.A(clknet_0__0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0899_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0899_ (.A(clknet_0__0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0899_));
 sky130_fd_sc_hd__clkinv_1 clkload303 (.A(clknet_1_0__leaf__0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0901_ (.A(_0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0901_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0901_ (.A(clknet_0__0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0901_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0901_ (.A(clknet_0__0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0901_));
 sky130_fd_sc_hd__clkbuf_4 clkload304 (.A(clknet_1_1__leaf__0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0900_ (.A(_0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0900_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0900_ (.A(clknet_0__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0900_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0900_ (.A(clknet_0__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0900_));
 sky130_fd_sc_hd__inv_4 clkload305 (.A(clknet_1_1__leaf__0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0663_ (.A(_0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0663_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0663_ (.A(clknet_0__0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0663_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0663_ (.A(clknet_0__0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0663_));
 sky130_fd_sc_hd__clkbuf_4 clkload306 (.A(clknet_1_0__leaf__0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload307 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0709_ (.A(_0709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0709_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0709_ (.A(clknet_0__0709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0709_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0709_ (.A(clknet_0__0709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0709_));
 sky130_fd_sc_hd__clkbuf_4 clkload308 (.A(clknet_1_1__leaf__0709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0710_ (.A(_0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0710_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0710_ (.A(clknet_0__0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0710_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0710_ (.A(clknet_0__0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0710_));
 sky130_fd_sc_hd__clkbuf_4 clkload309 (.A(clknet_1_0__leaf__0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0711_ (.A(_0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0711_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0711_ (.A(clknet_0__0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0711_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0711_ (.A(clknet_0__0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0711_));
 sky130_fd_sc_hd__clkbuf_4 clkload310 (.A(clknet_1_1__leaf__0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ));
 sky130_fd_sc_hd__clkbuf_4 clkload311 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload312 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0219_ (.A(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0219_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0219_ (.A(clknet_0__0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0219_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0219_ (.A(clknet_0__0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0219_));
 sky130_fd_sc_hd__clkbuf_4 clkload313 (.A(clknet_1_0__leaf__0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0222_ (.A(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0222_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0222_ (.A(clknet_0__0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0222_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0222_ (.A(clknet_0__0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0222_));
 sky130_fd_sc_hd__clkbuf_4 clkload314 (.A(clknet_1_1__leaf__0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0225_ (.A(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0225_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0225_ (.A(clknet_0__0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0225_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0225_ (.A(clknet_0__0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0225_));
 sky130_fd_sc_hd__clkinv_2 clkload315 (.A(clknet_1_1__leaf__0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0228_ (.A(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0228_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0228_ (.A(clknet_0__0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0228_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0228_ (.A(clknet_0__0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0228_));
 sky130_fd_sc_hd__inv_2 clkload316 (.A(clknet_1_1__leaf__0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0233_ (.A(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0233_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0233_ (.A(clknet_0__0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0233_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0233_ (.A(clknet_0__0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0233_));
 sky130_fd_sc_hd__clkinv_1 clkload317 (.A(clknet_1_1__leaf__0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0227_ (.A(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0227_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0227_ (.A(clknet_0__0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0227_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0227_ (.A(clknet_0__0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0227_));
 sky130_fd_sc_hd__clkbuf_4 clkload318 (.A(clknet_1_0__leaf__0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0224_ (.A(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0224_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0224_ (.A(clknet_0__0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0224_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0224_ (.A(clknet_0__0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0224_));
 sky130_fd_sc_hd__clkbuf_4 clkload319 (.A(clknet_1_0__leaf__0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload320 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0563_ (.A(_0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0563_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0563_ (.A(clknet_0__0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0563_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0563_ (.A(clknet_0__0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0563_));
 sky130_fd_sc_hd__clkbuf_8 clkload321 (.A(clknet_1_1__leaf__0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0566_ (.A(_0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0566_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0566_ (.A(clknet_0__0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0566_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0566_ (.A(clknet_0__0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0566_));
 sky130_fd_sc_hd__clkbuf_4 clkload322 (.A(clknet_1_1__leaf__0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0565_ (.A(_0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0565_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0565_ (.A(clknet_0__0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0565_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0565_ (.A(clknet_0__0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0565_));
 sky130_fd_sc_hd__bufinv_8 clkload323 (.A(clknet_1_0__leaf__0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0564_ (.A(_0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0564_ (.A(clknet_0__0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0564_ (.A(clknet_0__0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0564_));
 sky130_fd_sc_hd__clkbuf_4 clkload324 (.A(clknet_1_0__leaf__0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0221_ (.A(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0221_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0221_ (.A(clknet_0__0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0221_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0221_ (.A(clknet_0__0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0221_));
 sky130_fd_sc_hd__clkbuf_4 clkload325 (.A(clknet_1_1__leaf__0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkinv_1 clkload326 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0559_ (.A(_0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0559_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0559_ (.A(clknet_0__0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0559_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0559_ (.A(clknet_0__0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0559_));
 sky130_fd_sc_hd__clkbuf_4 clkload327 (.A(clknet_1_1__leaf__0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0562_ (.A(_0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0562_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0562_ (.A(clknet_0__0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0562_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0562_ (.A(clknet_0__0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0562_));
 sky130_fd_sc_hd__clkinv_1 clkload328 (.A(clknet_1_1__leaf__0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0561_ (.A(_0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0561_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0561_ (.A(clknet_0__0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0561_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0561_ (.A(clknet_0__0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0561_));
 sky130_fd_sc_hd__clkbuf_4 clkload329 (.A(clknet_1_0__leaf__0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload330 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0607_ (.A(_0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0607_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0607_ (.A(clknet_0__0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0607_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0607_ (.A(clknet_0__0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0607_));
 sky130_fd_sc_hd__clkbuf_4 clkload331 (.A(clknet_1_0__leaf__0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0609_ (.A(_0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0609_ (.A(clknet_0__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0609_ (.A(clknet_0__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0609_));
 sky130_fd_sc_hd__bufinv_8 clkload332 (.A(clknet_1_0__leaf__0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload333 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload334 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_4 clkload335 (.A(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0589_ (.A(_0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0589_ (.A(clknet_0__0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0589_ (.A(clknet_0__0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0589_));
 sky130_fd_sc_hd__clkbuf_4 clkload336 (.A(clknet_1_0__leaf__0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0590_ (.A(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0590_ (.A(clknet_0__0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0590_ (.A(clknet_0__0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0590_));
 sky130_fd_sc_hd__clkbuf_4 clkload337 (.A(clknet_1_1__leaf__0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0232_ (.A(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0232_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0232_ (.A(clknet_0__0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0232_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0232_ (.A(clknet_0__0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0232_));
 sky130_fd_sc_hd__clkbuf_4 clkload338 (.A(clknet_1_1__leaf__0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload339 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload340 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0620_ (.A(_0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0620_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0620_ (.A(clknet_0__0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0620_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0620_ (.A(clknet_0__0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0620_));
 sky130_fd_sc_hd__clkbuf_4 clkload341 (.A(clknet_1_0__leaf__0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0537_ (.A(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0537_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0537_ (.A(clknet_0__0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0537_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0537_ (.A(clknet_0__0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0537_));
 sky130_fd_sc_hd__clkbuf_4 clkload342 (.A(clknet_1_1__leaf__0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload343 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0596_ (.A(_0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0596_ (.A(clknet_0__0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0596_ (.A(clknet_0__0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0596_));
 sky130_fd_sc_hd__bufinv_16 clkload344 (.A(clknet_1_0__leaf__0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload345 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload346 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0595_ (.A(_0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0595_ (.A(clknet_0__0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0595_ (.A(clknet_0__0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0595_));
 sky130_fd_sc_hd__clkbuf_4 clkload347 (.A(clknet_1_1__leaf__0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload348 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cby_2__2_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ));
 sky130_fd_sc_hd__clkbuf_4 clkload349 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0231_ (.A(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0231_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0231_ (.A(clknet_0__0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0231_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0231_ (.A(clknet_0__0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0231_));
 sky130_fd_sc_hd__clkbuf_4 clkload350 (.A(clknet_1_1__leaf__0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in  (.A(\clknet_0_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ));
 sky130_fd_sc_hd__clkinv_1 clkload351 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.direct_interc_0_.in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0560_ (.A(_0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0560_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0560_ (.A(clknet_0__0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0560_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0560_ (.A(clknet_0__0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0560_));
 sky130_fd_sc_hd__clkbuf_4 clkload352 (.A(clknet_1_1__leaf__0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0536_ (.A(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0536_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0536_ (.A(clknet_0__0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0536_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0536_ (.A(clknet_0__0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0536_));
 sky130_fd_sc_hd__clkbuf_4 clkload353 (.A(clknet_1_0__leaf__0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0202_ (.A(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0202_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0202_ (.A(clknet_0__0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0202_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0202_ (.A(clknet_0__0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0202_));
 sky130_fd_sc_hd__clkbuf_4 clkload354 (.A(clknet_1_1__leaf__0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload355 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_2__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0197_ (.A(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0197_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0197_ (.A(clknet_0__0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0197_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0197_ (.A(clknet_0__0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0197_));
 sky130_fd_sc_hd__clkbuf_4 clkload356 (.A(clknet_1_1__leaf__0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0586_ (.A(_0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0586_ (.A(clknet_0__0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0586_ (.A(clknet_0__0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0586_));
 sky130_fd_sc_hd__clkbuf_4 clkload357 (.A(clknet_1_0__leaf__0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0549_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0549_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0549_ (.A(clknet_0__0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0549_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0549_ (.A(clknet_0__0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0549_));
 sky130_fd_sc_hd__clkbuf_4 clkload358 (.A(clknet_1_0__leaf__0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0615_ (.A(_0615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0615_ (.A(clknet_0__0615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0615_ (.A(clknet_0__0615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0615_));
 sky130_fd_sc_hd__bufinv_8 clkload359 (.A(clknet_1_1__leaf__0615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0617_ (.A(_0617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0617_ (.A(clknet_0__0617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0617_ (.A(clknet_0__0617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0617_));
 sky130_fd_sc_hd__bufinv_16 clkload360 (.A(clknet_1_1__leaf__0617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0193_ (.A(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0193_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0193_ (.A(clknet_0__0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0193_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0193_ (.A(clknet_0__0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0193_));
 sky130_fd_sc_hd__clkinv_1 clkload361 (.A(clknet_1_1__leaf__0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net31 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net31));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net31 (.A(clknet_0_net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net31));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net31 (.A(clknet_0_net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net31));
 sky130_fd_sc_hd__bufinv_8 clkload362 (.A(clknet_1_1__leaf_net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net29 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net29 (.A(clknet_0_net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net29 (.A(clknet_0_net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net29));
 sky130_fd_sc_hd__clkbuf_8 clkload363 (.A(clknet_1_1__leaf_net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net23 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net23 (.A(clknet_0_net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net23));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net23 (.A(clknet_0_net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net23));
 sky130_fd_sc_hd__clkbuf_4 clkload364 (.A(clknet_1_1__leaf_net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out  (.A(\clknet_0_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clknet_1_1__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__clkinv_1 clkload365 (.A(\clknet_1_0__leaf_dut_0.U0_formal_verification.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0220_ (.A(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0__0220_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0220_ (.A(clknet_0__0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf__0220_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0220_ (.A(clknet_0__0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf__0220_));
 sky130_fd_sc_hd__clkbuf_4 clkload366 (.A(clknet_1_0__leaf__0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net52 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_net52));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net52 (.A(clknet_0_net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_net52));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net52 (.A(clknet_0_net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_net52));
 sky130_fd_sc_hd__clkinv_1 clkload367 (.A(clknet_1_0__leaf_net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\dut_0.U0_formal_verification.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\dut_0.U0_formal_verification.cby_1__2_.mux_left_ipin_0.mux_l3_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\dut_0.U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\dut_0.U0_formal_verification.sb_2__0_.mem_left_track_5.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_9.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(clknet_1_0__leaf__0820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__6.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(clknet_1_1__leaf__0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\clknet_1_0__leaf_dut_0.U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__3.gfpga_pad_GPIO_PAD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\dut_0.U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.DFF_0_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\dut_0.U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\clknet_1_1__leaf_dut_0.U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\dut_0.U0_formal_verification.sb_2__2_.mem_bottom_track_13.DFF_1_.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_408 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_511 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_523 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_707 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_797 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_825 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_849 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_869 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_881 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_909 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_997 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_86 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_98 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_1_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_185 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_1_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_262 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_604 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_1_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_635 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_749 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_772 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_1_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_835 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_847 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_934 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_942 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_999 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_1_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_2_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_2_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_2_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_509 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_603 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_2_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_728 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_754 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_774 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_801 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_846 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_2_858 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_866 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_873 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_2_885 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_941 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_974 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_999 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1011 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1023 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_82 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_185 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_3_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_603 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_3_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_797 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_809 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_821 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_841 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_853 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_888 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_909 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_929 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_971 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_991 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_3_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_612 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_707 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_748 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_766 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_770 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_796 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_808 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_832 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_844 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_856 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_866 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_880 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_901 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_4_913 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_963 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_976 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_1007 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1019 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_40 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_185 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_5_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_256 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_5_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_577 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_5_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_648 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_660 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_769 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_801 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_841 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_853 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_857 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_872 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_884 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_888 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_918 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_1002 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_1025 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_5_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_5_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_217 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_229 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_6_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_668 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_680 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_738 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_849 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_878 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_898 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_966 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_1006 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1018 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_7_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_655 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_705 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_732 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_766 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_868 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_876 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_911 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_962 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_974 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_7_986 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_1004 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_7_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_605 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_763 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_866 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_869 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_8_881 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_908 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_912 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_916 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_937 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_998 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1010 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1022 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_9_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_516 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_9_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_550 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_598 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_633 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_9_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_815 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_834 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_875 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_9_887 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_903 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_927 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_935 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_9_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_10_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_540 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_606 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_628 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_659 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_777 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_10_789 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_825 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_847 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_885 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_937 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_941 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_958 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_968 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1001 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1013 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_11_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_760 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_877 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_11_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_957 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_969 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_993 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_11_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_1034 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1046 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_11_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_11_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_767 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_771 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_810 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_907 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_942 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_985 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_13_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_13_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_702 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_834 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_884 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_901 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_940 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_1018 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_1036 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1048 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_1060 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_13_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_72 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_14_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_14_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_650 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_662 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_674 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_686 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_14_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_817 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_911 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_975 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_990 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_996 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_15_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_15_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_15_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_720 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_758 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_835 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_884 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_913 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_15_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_942 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_976 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_1035 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1047 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_1059 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_15_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_16_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_16_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_908 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_1021 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_703 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_771 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_17_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_830 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_904 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_947 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_1000 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_1046 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_17_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_17_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_18_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_108 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_728 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_734 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_877 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_997 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_1028 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_19_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_478 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_538 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_707 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_735 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_754 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_775 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_803 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_19_815 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_838 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_875 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_887 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_907 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_916 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_928 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_936 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_1025 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_19_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_19_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_40 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_20_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_751 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_795 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_824 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_865 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_891 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_903 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_20_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_957 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_978 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_997 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_20_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_82 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_21_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_745 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_21_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_823 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_831 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_927 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_953 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_989 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_21_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_740 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_776 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_22_788 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_831 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_843 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_855 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_22_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_899 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_949 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_965 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_993 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_23_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_95 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_23_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_748 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_772 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_789 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_832 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_859 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_23_871 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_904 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_23_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_1002 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_23_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_810 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_839 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_851 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_24_863 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_869 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_24_881 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_898 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_914 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_941 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_961 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_24_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_990 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_1007 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_1019 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_24_1031 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_25_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_762 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_770 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_791 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_802 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_808 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_832 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_845 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_864 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_876 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_888 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_912 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_935 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_980 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_738 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_761 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_800 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_26_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_885 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_902 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_931 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_957 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_963 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_1013 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_73 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_27_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_716 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_744 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_770 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_27_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_827 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_838 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_962 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_1004 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_1028 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_1040 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_1052 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_27_1065 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_1082 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_28_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_799 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_862 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_914 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_1022 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_1032 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_28_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_882 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_29_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_999 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_1022 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_1040 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_1060 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_30_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_575 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_748 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_761 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_779 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_826 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_866 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_869 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_881 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_902 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_978 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_997 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_30_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_1071 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_662 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_738 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_756 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_768 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_31_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_797 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_809 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_31_821 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_829 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_888 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_913 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_938 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_962 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_966 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_983 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_995 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_1017 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_1065 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_1087 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_749 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_769 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_781 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_793 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_32_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_817 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_843 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_847 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_885 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_957 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_32_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_985 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_1027 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_20 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_606 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_716 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_749 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_766 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_850 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_948 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_994 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_1013 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_1020 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_751 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_773 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_795 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_808 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_850 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_854 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_898 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_989 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_1008 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_37 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_732 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_744 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_756 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_776 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_822 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_913 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_959 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_980 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_986 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_1013 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_36_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_537 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_564 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_674 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_744 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_780 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_36_792 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_862 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_968 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_36_993 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_1053 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_37_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_751 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_37_797 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_931 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_978 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_997 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_1032 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_1036 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_1054 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_1069 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_38_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_47 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_38_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_622 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_749 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_761 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_786 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_806 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_829 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_860 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_886 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_916 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_38_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_38_993 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_1015 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_1019 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_38_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_1069 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_1087 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_39_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_737 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_791 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_39_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_822 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_863 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_871 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_891 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_39_909 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_39_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_927 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_957 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_976 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_984 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_39_1021 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_1044 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_1071 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_1088 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_40_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_40_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_728 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_40_740 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_40_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_789 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_793 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_40_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_40_825 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_40_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_843 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_874 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_898 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_939 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_40_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_955 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_974 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_40_993 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_1028 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_1088 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_520 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_41_532 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_714 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_41_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_41_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_749 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_41_761 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_41_797 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_41_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_820 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_41_832 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_41_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_918 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_928 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_939 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_41_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_958 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_988 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_41_1021 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_1070 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_636 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_748 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_774 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_793 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_801 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_829 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_42_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_941 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_960 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_42_1057 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_42_1069 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_42_1081 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_43_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_483 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_43_495 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_723 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_749 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_43_761 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_43_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_43_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_793 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_913 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_971 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_1043 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_43_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_1072 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_43_1084 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_44_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_721 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_733 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_44_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_775 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_787 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_44_799 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_824 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_900 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_1022 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_1067 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_45_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_486 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_729 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_45_741 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_45_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_774 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_778 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_790 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_800 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_1003 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_1047 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_45_1062 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_1068 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_750 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_46_769 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_828 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_952 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_1024 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_46_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_1045 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_1060 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_46_1072 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_47_758 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_47_790 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_798 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_1032 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_47_1044 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_47_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_745 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_778 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_48_806 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_48_825 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_845 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_972 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_985 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_48_1030 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_1043 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_48_1055 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_1072 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_48_1084 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_508 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_735 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_49_747 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_772 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_49_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_49_797 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_820 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_828 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_835 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_857 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_904 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_1048 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_49_1060 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_49_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_596 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_715 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_736 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_50_748 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_769 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_781 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_793 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_50_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_825 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_50_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_845 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_904 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_935 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_959 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_50_1004 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_1012 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_1054 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_1071 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_751 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_51_763 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_51_775 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_804 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_51_816 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_820 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_841 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_51_853 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_883 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_943 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_973 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_992 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_51_1004 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_1017 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_1056 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_1065 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_463 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_810 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_842 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_862 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_869 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_52_881 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_988 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_1010 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_52_1022 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_52_1049 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_1053 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_1070 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_761 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_53_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_810 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_836 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_847 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_880 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_53_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_903 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_913 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_986 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_1018 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_53_1030 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_53_1042 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_53_1054 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_571 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_731 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_54_743 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_885 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_54_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_54_909 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_976 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_989 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_1024 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_54_1053 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_1070 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_478 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_729 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_55_741 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_749 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_760 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_55_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_837 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_868 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_55_880 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_55_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_55_909 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_929 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_985 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_993 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_1049 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_55_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_706 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_754 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_784 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_806 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_836 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_56_848 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_56_860 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_877 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_911 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_56_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_936 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_966 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_976 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_989 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_1024 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_1081 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_57_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_523 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_692 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_738 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_57_750 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_57_762 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_821 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_57_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_847 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_908 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_57_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_942 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_975 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_57_987 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_1013 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_1053 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_57_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_58_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_720 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_724 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_58_736 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_58_748 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_773 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_58_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_822 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_861 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_905 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_58_937 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_945 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_952 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_999 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_1021 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_550 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_59_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_59_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_703 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_59_715 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_59_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_747 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_802 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_59_814 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_822 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_860 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_59_872 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_878 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_59_909 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_59_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_929 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_996 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_1000 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_1017 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_1081 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_60_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_60_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_60_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_60_713 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_719 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_747 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_757 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_791 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_60_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_813 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_60_825 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_850 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_60_862 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_890 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_60_902 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_60_914 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_60_918 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_937 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_60_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_981 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_987 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_60_999 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_1062 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_1066 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_60_1083 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_61_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_61_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_478 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_705 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_750 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_778 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_789 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_797 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_801 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_819 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_827 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_858 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_866 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_885 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_937 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_943 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_1009 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_1017 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_1059 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_1065 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_62_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_48 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_62_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_616 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_740 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_62_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_764 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_62_776 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_784 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_809 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_62_818 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_863 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_878 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_62_890 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_939 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_62_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_955 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_965 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_979 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_62_1064 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_1086 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_1090 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_63_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_678 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_63_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_754 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_774 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_800 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_817 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_855 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_867 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_879 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_63_891 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_63_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_967 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_993 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_63_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_63_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_1051 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_1065 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_63_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_64_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_64_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_752 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_762 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_810 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_827 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_858 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_864 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_880 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_892 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_904 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_64_916 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_64_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_957 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_997 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_64_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_65_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_703 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_830 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_888 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_909 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_65_921 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_65_930 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_953 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_65_965 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_1000 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_1025 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_65_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_65_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_66_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_46 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_66_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_677 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_66_760 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_816 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_66_916 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_943 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_955 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_66_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_87 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_67_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_637 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_649 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_67_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_67_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_762 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_827 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_67_916 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_1041 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_67_1053 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_67_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_68_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_68_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_68_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_682 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_718 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_766 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_787 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_791 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_68_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_821 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_863 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_880 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_903 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_919 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_68_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_69_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_69_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_590 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_69_602 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_637 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_649 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_69_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_69_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_69_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_706 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_714 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_723 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_735 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_756 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_779 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_783 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_69_797 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_835 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_846 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_886 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_905 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_910 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_922 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_934 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_946 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_953 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_69_965 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_69_978 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_1034 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_1046 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_1058 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_69_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_148 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_70_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_70_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_674 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_686 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_70_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_764 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_817 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_823 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_835 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_847 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_886 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_894 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_941 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_70_1010 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_71_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_71_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_71_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_71_595 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_626 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_71_638 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_71_646 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_71_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_734 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_71_746 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_756 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_71_768 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_776 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_785 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_817 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_828 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_71_859 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_878 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_890 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_927 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_944 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_1000 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_1025 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_71_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_71_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_52 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_72_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_72_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_450 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_656 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_676 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_743 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_755 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_779 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_824 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_72_836 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_857 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_867 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_888 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_72_900 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_918 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_954 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_72_966 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_970 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_990 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_72_1025 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_20 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_32 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_73_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_73_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_524 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_73_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_579 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_599 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_73_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_628 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_729 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_73_741 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_770 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_780 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_73_792 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_817 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_834 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_841 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_73_853 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_870 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_73_909 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_73_942 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_950 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_73_1000 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_73_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_74_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_74_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_74_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_74_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_592 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_74_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_74_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_722 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_74_734 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_738 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_74_764 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_784 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_802 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_74_822 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_889 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_914 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_943 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_955 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_961 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_978 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_1010 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_1022 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_37 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_75_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_75_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_510 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_75_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_544 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_75_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_587 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_599 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_75_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_741 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_753 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_765 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_797 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_809 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_75_821 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_832 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_841 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_75_853 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_892 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_897 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_909 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_921 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_75_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_946 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_953 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_973 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_985 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_75_997 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_75_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_75_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_76_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_160 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_172 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_76_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_517 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_547 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_76_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_566 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_574 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_76_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_76_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_76_622 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_733 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_779 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_791 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_76_803 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_822 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_828 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_861 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_869 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_933 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_968 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_993 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_77_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_40 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_77_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_77_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_77_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_77_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_491 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_77_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_77_516 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_77_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_77_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_579 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_77_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_77_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_716 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_749 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_770 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_77_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_77_794 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_838 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_77_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_897 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_77_915 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_939 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_77_951 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_961 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_77_973 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_77_985 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_77_997 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_77_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_77_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_78_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_78_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_78_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_494 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_78_506 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_78_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_78_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_658 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_675 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_773 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_807 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_811 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_78_833 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_839 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_78_860 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_923 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_925 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_935 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_945 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_957 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_78_969 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_993 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_1061 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_1073 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_79_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_79_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_79_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_142 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_79_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_79_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_79_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_79_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_79_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_79_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_79_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_700 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_737 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_79_751 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_759 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_770 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_79_782 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_794 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_79_841 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_79_893 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_79_913 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_946 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_953 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_965 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_977 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_989 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_79_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_80_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_80_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_80_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_80_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_484 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_80_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_80_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_660 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_80_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_80_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_729 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_741 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_753 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_757 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_769 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_781 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_785 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_80_797 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_805 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_813 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_80_830 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_838 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_841 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_853 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_865 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_80_878 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_886 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_80_891 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_895 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_917 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_922 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_925 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_937 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_949 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_953 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_965 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_977 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_981 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_993 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_1005 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_1009 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_1021 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_1033 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_80_1061 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_1065 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_1077 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_80_1089 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net223;
 assign uio_oe[1] = net224;
 assign uio_oe[2] = net225;
 assign uio_oe[3] = net226;
 assign uio_oe[4] = net227;
 assign uio_oe[5] = net233;
 assign uio_oe[6] = net234;
 assign uio_oe[7] = net235;
 assign uio_out[0] = net228;
 assign uio_out[1] = net229;
 assign uio_out[2] = net230;
 assign uio_out[3] = net231;
 assign uio_out[4] = net232;
endmodule
