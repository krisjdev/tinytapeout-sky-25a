module tt_um_swangust3 (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire net114;
 wire clknet_leaf_0_clk;
 wire net97;
 wire \p8div.B_decode.F[0] ;
 wire \p8div.B_decode.F[1] ;
 wire \p8div.B_decode.F[2] ;
 wire \p8div.B_decode.F[3] ;
 wire \p8div.B_decode.F[4] ;
 wire \p8div.a_piped[0] ;
 wire \p8div.a_piped[1] ;
 wire \p8div.a_piped[2] ;
 wire \p8div.a_piped[3] ;
 wire \p8div.a_piped[4] ;
 wire \p8div.a_piped[5] ;
 wire \p8div.a_piped[6] ;
 wire \p8div.a_piped[7] ;
 wire \p8div.b_piped[0] ;
 wire \p8div.b_piped[1] ;
 wire \p8div.b_piped[2] ;
 wire \p8div.b_piped[3] ;
 wire \p8div.b_piped[4] ;
 wire \p8div.b_piped[5] ;
 wire \p8div.b_piped[6] ;
 wire \p8div.c_decoded[10] ;
 wire \p8div.c_decoded[11] ;
 wire \p8div.c_decoded[1] ;
 wire \p8div.c_decoded[2] ;
 wire \p8div.c_decoded[3] ;
 wire \p8div.c_decoded[4] ;
 wire \p8div.c_decoded[5] ;
 wire \p8div.c_decoded[6] ;
 wire \p8div.c_decoded[7] ;
 wire \p8div.c_decoded[8] ;
 wire \p8div.c_decoded[9] ;
 wire \p8div.c_scale[0] ;
 wire \p8div.c_scale[1] ;
 wire \p8div.c_scale[2] ;
 wire \p8div.c_scale[3] ;
 wire \p8div.c_scale[4] ;
 wire \p8div.d_sign ;
 wire \p8div.pipe_A.a_q[0][0] ;
 wire \p8div.pipe_A.a_q[0][1] ;
 wire \p8div.pipe_A.a_q[0][2] ;
 wire \p8div.pipe_A.a_q[0][3] ;
 wire \p8div.pipe_A.a_q[0][4] ;
 wire \p8div.pipe_A.a_q[0][5] ;
 wire \p8div.pipe_A.a_q[0][6] ;
 wire \p8div.pipe_A.a_q[0][7] ;
 wire \p8div.pipe_A.a_q[1][0] ;
 wire \p8div.pipe_A.a_q[1][1] ;
 wire \p8div.pipe_A.a_q[1][2] ;
 wire \p8div.pipe_A.a_q[1][3] ;
 wire \p8div.pipe_A.a_q[1][4] ;
 wire \p8div.pipe_A.a_q[1][5] ;
 wire \p8div.pipe_A.a_q[1][6] ;
 wire \p8div.pipe_A.a_q[1][7] ;
 wire \p8div.pipe_A.a_q[2][0] ;
 wire \p8div.pipe_A.a_q[2][1] ;
 wire \p8div.pipe_A.a_q[2][2] ;
 wire \p8div.pipe_A.a_q[2][3] ;
 wire \p8div.pipe_A.a_q[2][4] ;
 wire \p8div.pipe_A.a_q[2][5] ;
 wire \p8div.pipe_A.a_q[2][6] ;
 wire \p8div.pipe_A.a_q[2][7] ;
 wire \p8div.pipe_A.a_q[3][0] ;
 wire \p8div.pipe_A.a_q[3][1] ;
 wire \p8div.pipe_A.a_q[3][2] ;
 wire \p8div.pipe_A.a_q[3][3] ;
 wire \p8div.pipe_A.a_q[3][4] ;
 wire \p8div.pipe_A.a_q[3][5] ;
 wire \p8div.pipe_A.a_q[3][6] ;
 wire \p8div.pipe_A.a_q[3][7] ;
 wire \p8div.pipe_A.a_q[4][0] ;
 wire \p8div.pipe_A.a_q[4][1] ;
 wire \p8div.pipe_A.a_q[4][2] ;
 wire \p8div.pipe_A.a_q[4][3] ;
 wire \p8div.pipe_A.a_q[4][4] ;
 wire \p8div.pipe_A.a_q[4][5] ;
 wire \p8div.pipe_A.a_q[4][6] ;
 wire \p8div.pipe_A.a_q[4][7] ;
 wire \p8div.pipe_A.a_q[5][0] ;
 wire \p8div.pipe_A.a_q[5][1] ;
 wire \p8div.pipe_A.a_q[5][2] ;
 wire \p8div.pipe_A.a_q[5][3] ;
 wire \p8div.pipe_A.a_q[5][4] ;
 wire \p8div.pipe_A.a_q[5][5] ;
 wire \p8div.pipe_A.a_q[5][6] ;
 wire \p8div.pipe_A.a_q[5][7] ;
 wire \p8div.pipe_A.a_q[6][0] ;
 wire \p8div.pipe_A.a_q[6][1] ;
 wire \p8div.pipe_A.a_q[6][2] ;
 wire \p8div.pipe_A.a_q[6][3] ;
 wire \p8div.pipe_A.a_q[6][4] ;
 wire \p8div.pipe_A.a_q[6][5] ;
 wire \p8div.pipe_A.a_q[6][6] ;
 wire \p8div.pipe_A.a_q[6][7] ;
 wire \p8div.pipe_A.a_q[7][0] ;
 wire \p8div.pipe_A.a_q[7][1] ;
 wire \p8div.pipe_A.a_q[7][2] ;
 wire \p8div.pipe_A.a_q[7][3] ;
 wire \p8div.pipe_A.a_q[7][4] ;
 wire \p8div.pipe_A.a_q[7][5] ;
 wire \p8div.pipe_A.a_q[7][6] ;
 wire \p8div.pipe_A.a_q[7][7] ;
 wire \p8div.pipe_A.a_q[8][0] ;
 wire \p8div.pipe_A.a_q[8][1] ;
 wire \p8div.pipe_A.a_q[8][2] ;
 wire \p8div.pipe_A.a_q[8][3] ;
 wire \p8div.pipe_A.a_q[8][4] ;
 wire \p8div.pipe_A.a_q[8][5] ;
 wire \p8div.pipe_A.a_q[8][6] ;
 wire \p8div.pipe_A.a_q[8][7] ;
 wire \p8div.pipe_A.a_q[9][0] ;
 wire \p8div.pipe_A.a_q[9][1] ;
 wire \p8div.pipe_A.a_q[9][2] ;
 wire \p8div.pipe_A.a_q[9][3] ;
 wire \p8div.pipe_A.a_q[9][4] ;
 wire \p8div.pipe_A.a_q[9][5] ;
 wire \p8div.pipe_A.a_q[9][6] ;
 wire \p8div.pipe_A.a_q[9][7] ;
 wire \p8div.pipe_B.a_q[0][0] ;
 wire \p8div.pipe_B.a_q[0][1] ;
 wire \p8div.pipe_B.a_q[0][2] ;
 wire \p8div.pipe_B.a_q[0][3] ;
 wire \p8div.pipe_B.a_q[0][4] ;
 wire \p8div.pipe_B.a_q[0][5] ;
 wire \p8div.pipe_B.a_q[0][6] ;
 wire \p8div.pipe_B.a_q[1][0] ;
 wire \p8div.pipe_B.a_q[1][1] ;
 wire \p8div.pipe_B.a_q[1][2] ;
 wire \p8div.pipe_B.a_q[1][3] ;
 wire \p8div.pipe_B.a_q[1][4] ;
 wire \p8div.pipe_B.a_q[1][5] ;
 wire \p8div.pipe_B.a_q[1][6] ;
 wire \p8div.pipe_B.a_q[2][0] ;
 wire \p8div.pipe_B.a_q[2][1] ;
 wire \p8div.pipe_B.a_q[2][2] ;
 wire \p8div.pipe_B.a_q[2][3] ;
 wire \p8div.pipe_B.a_q[2][4] ;
 wire \p8div.pipe_B.a_q[2][5] ;
 wire \p8div.pipe_B.a_q[2][6] ;
 wire \p8div.pipe_B.a_q[3][0] ;
 wire \p8div.pipe_B.a_q[3][1] ;
 wire \p8div.pipe_B.a_q[3][2] ;
 wire \p8div.pipe_B.a_q[3][3] ;
 wire \p8div.pipe_B.a_q[3][4] ;
 wire \p8div.pipe_B.a_q[3][5] ;
 wire \p8div.pipe_B.a_q[3][6] ;
 wire \p8div.pipe_B.a_q[4][0] ;
 wire \p8div.pipe_B.a_q[4][1] ;
 wire \p8div.pipe_B.a_q[4][2] ;
 wire \p8div.pipe_B.a_q[4][3] ;
 wire \p8div.pipe_B.a_q[4][4] ;
 wire \p8div.pipe_B.a_q[4][5] ;
 wire \p8div.pipe_B.a_q[4][6] ;
 wire \p8div.pipe_B.a_q[5][0] ;
 wire \p8div.pipe_B.a_q[5][1] ;
 wire \p8div.pipe_B.a_q[5][2] ;
 wire \p8div.pipe_B.a_q[5][3] ;
 wire \p8div.pipe_B.a_q[5][4] ;
 wire \p8div.pipe_B.a_q[5][5] ;
 wire \p8div.pipe_B.a_q[5][6] ;
 wire \p8div.pipe_B.a_q[6][0] ;
 wire \p8div.pipe_B.a_q[6][1] ;
 wire \p8div.pipe_B.a_q[6][2] ;
 wire \p8div.pipe_B.a_q[6][3] ;
 wire \p8div.pipe_B.a_q[6][4] ;
 wire \p8div.pipe_B.a_q[6][5] ;
 wire \p8div.pipe_B.a_q[6][6] ;
 wire \p8div.pipe_B.a_q[7][0] ;
 wire \p8div.pipe_B.a_q[7][1] ;
 wire \p8div.pipe_B.a_q[7][2] ;
 wire \p8div.pipe_B.a_q[7][3] ;
 wire \p8div.pipe_B.a_q[7][4] ;
 wire \p8div.pipe_B.a_q[7][5] ;
 wire \p8div.pipe_B.a_q[7][6] ;
 wire \p8div.pipe_B.a_q[8][0] ;
 wire \p8div.pipe_B.a_q[8][1] ;
 wire \p8div.pipe_B.a_q[8][2] ;
 wire \p8div.pipe_B.a_q[8][3] ;
 wire \p8div.pipe_B.a_q[8][4] ;
 wire \p8div.pipe_B.a_q[8][5] ;
 wire \p8div.pipe_B.a_q[8][6] ;
 wire \p8div.pipe_B.a_q[9][0] ;
 wire \p8div.pipe_B.a_q[9][1] ;
 wire \p8div.pipe_B.a_q[9][2] ;
 wire \p8div.pipe_B.a_q[9][3] ;
 wire \p8div.pipe_B.a_q[9][4] ;
 wire \p8div.pipe_B.a_q[9][5] ;
 wire \p8div.pipe_B.a_q[9][6] ;
 wire \p8div.pipe_sign.A ;
 wire \p8div.pipe_sign.a_q[0] ;
 wire \p8div.pipe_sign.a_q[1] ;
 wire \p8div.pipe_sign.a_q[2] ;
 wire \p8div.pipe_sign.a_q[3] ;
 wire \p8div.pipe_sign.a_q[4] ;
 wire \p8div.pipe_sign.a_q[5] ;
 wire \p8div.pipe_sign.a_q[6] ;
 wire \p8div.pipe_sign.a_q[7] ;
 wire \p8div.pipe_sign.a_q[8] ;
 wire \p8div.pipe_sign.a_q[9] ;
 wire \p8div.sa.add_frac_sum_a.C ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_0_HCA.hca_stage_0.SUM ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.acc[10][0] ;
 wire \p8div.sa.div.acc[10][1] ;
 wire \p8div.sa.div.acc[10][2] ;
 wire \p8div.sa.div.acc[10][3] ;
 wire \p8div.sa.div.acc[10][4] ;
 wire \p8div.sa.div.acc[10][5] ;
 wire \p8div.sa.div.b[0][0] ;
 wire \p8div.sa.div.b[0][1] ;
 wire \p8div.sa.div.b[0][2] ;
 wire \p8div.sa.div.b[0][3] ;
 wire \p8div.sa.div.b[0][4] ;
 wire \p8div.sa.div.b[0][5] ;
 wire \p8div.sa.div.b[10][0] ;
 wire \p8div.sa.div.b[10][1] ;
 wire \p8div.sa.div.b[10][2] ;
 wire \p8div.sa.div.b[10][3] ;
 wire \p8div.sa.div.b[10][4] ;
 wire \p8div.sa.div.b[10][5] ;
 wire \p8div.sa.div.b[1][0] ;
 wire \p8div.sa.div.b[1][1] ;
 wire \p8div.sa.div.b[1][2] ;
 wire \p8div.sa.div.b[1][3] ;
 wire \p8div.sa.div.b[1][4] ;
 wire \p8div.sa.div.b[1][5] ;
 wire \p8div.sa.div.b[2][0] ;
 wire \p8div.sa.div.b[2][1] ;
 wire \p8div.sa.div.b[2][2] ;
 wire \p8div.sa.div.b[2][3] ;
 wire \p8div.sa.div.b[2][4] ;
 wire \p8div.sa.div.b[2][5] ;
 wire \p8div.sa.div.b[3][0] ;
 wire \p8div.sa.div.b[3][1] ;
 wire \p8div.sa.div.b[3][2] ;
 wire \p8div.sa.div.b[3][3] ;
 wire \p8div.sa.div.b[3][4] ;
 wire \p8div.sa.div.b[3][5] ;
 wire \p8div.sa.div.b[4][0] ;
 wire \p8div.sa.div.b[4][1] ;
 wire \p8div.sa.div.b[4][2] ;
 wire \p8div.sa.div.b[4][3] ;
 wire \p8div.sa.div.b[4][4] ;
 wire \p8div.sa.div.b[4][5] ;
 wire \p8div.sa.div.b[5][0] ;
 wire \p8div.sa.div.b[5][1] ;
 wire \p8div.sa.div.b[5][2] ;
 wire \p8div.sa.div.b[5][3] ;
 wire \p8div.sa.div.b[5][4] ;
 wire \p8div.sa.div.b[5][5] ;
 wire \p8div.sa.div.b[6][0] ;
 wire \p8div.sa.div.b[6][1] ;
 wire \p8div.sa.div.b[6][2] ;
 wire \p8div.sa.div.b[6][3] ;
 wire \p8div.sa.div.b[6][4] ;
 wire \p8div.sa.div.b[6][5] ;
 wire \p8div.sa.div.b[7][0] ;
 wire \p8div.sa.div.b[7][1] ;
 wire \p8div.sa.div.b[7][2] ;
 wire \p8div.sa.div.b[7][3] ;
 wire \p8div.sa.div.b[7][4] ;
 wire \p8div.sa.div.b[7][5] ;
 wire \p8div.sa.div.b[8][0] ;
 wire \p8div.sa.div.b[8][1] ;
 wire \p8div.sa.div.b[8][2] ;
 wire \p8div.sa.div.b[8][3] ;
 wire \p8div.sa.div.b[8][4] ;
 wire \p8div.sa.div.b[8][5] ;
 wire \p8div.sa.div.b[9][0] ;
 wire \p8div.sa.div.b[9][1] ;
 wire \p8div.sa.div.b[9][2] ;
 wire \p8div.sa.div.b[9][3] ;
 wire \p8div.sa.div.b[9][4] ;
 wire \p8div.sa.div.b[9][5] ;
 wire \p8div.sa.div.div_0.a_ge_b ;
 wire \p8div.sa.div.div_0.sub_acc.C ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[0] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[1] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[2] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[3] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[4] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[5] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[6] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[7] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[8] ;
 wire \p8div.sa.div.genblk1[10].div_n.Q_I[9] ;
 wire \p8div.sa.div.genblk1[10].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[1].div_n.Q_I ;
 wire \p8div.sa.div.genblk1[1].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[1].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[1].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[2].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[2].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[2].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[2].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[3].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[3].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[3].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[3].div_n.Q_O[3] ;
 wire \p8div.sa.div.genblk1[3].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[4].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[4].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[4].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[4].div_n.Q_O[3] ;
 wire \p8div.sa.div.genblk1[4].div_n.Q_O[4] ;
 wire \p8div.sa.div.genblk1[4].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[5].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[5].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[5].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[5].div_n.Q_O[3] ;
 wire \p8div.sa.div.genblk1[5].div_n.Q_O[4] ;
 wire \p8div.sa.div.genblk1[5].div_n.Q_O[5] ;
 wire \p8div.sa.div.genblk1[5].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[3] ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[4] ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[5] ;
 wire \p8div.sa.div.genblk1[6].div_n.Q_O[6] ;
 wire \p8div.sa.div.genblk1[6].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[3] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[4] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[5] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[6] ;
 wire \p8div.sa.div.genblk1[7].div_n.Q_O[7] ;
 wire \p8div.sa.div.genblk1[7].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[0] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[1] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[2] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[3] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[4] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[5] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[6] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[7] ;
 wire \p8div.sa.div.genblk1[8].div_n.Q_O[8] ;
 wire \p8div.sa.div.genblk1[8].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[9].div_n.a_ge_b ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ;
 wire \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ;
 wire \p8div.sa.pipe_scale_c.a_q[0][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[0][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[0][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[0][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[0][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[1][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[1][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[1][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[1][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[1][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[2][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[2][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[2][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[2][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[2][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[3][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[3][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[3][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[3][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[3][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[4][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[4][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[4][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[4][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[4][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[5][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[5][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[5][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[5][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[5][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[6][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[6][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[6][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[6][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[6][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[7][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[7][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[7][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[7][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[7][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[8][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[8][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[8][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[8][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[8][4] ;
 wire \p8div.sa.pipe_scale_c.a_q[9][0] ;
 wire \p8div.sa.pipe_scale_c.a_q[9][1] ;
 wire \p8div.sa.pipe_scale_c.a_q[9][2] ;
 wire \p8div.sa.pipe_scale_c.a_q[9][3] ;
 wire \p8div.sa.pipe_scale_c.a_q[9][4] ;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;

 sky130_fd_sc_hd__inv_2 _0487_ (.A(\p8div.sa.div.b[4][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0488_ (.A(\p8div.sa.div.b[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0489_ (.A(\p8div.sa.div.b[4][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(\p8div.sa.div.b[4][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(\p8div.sa.div.b[4][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0492_ (.A(\p8div.sa.div.b[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0493_ (.A(\p8div.sa.div.b[3][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0494_ (.A(\p8div.sa.div.b[3][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0495_ (.A(\p8div.sa.div.b[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\p8div.sa.div.b[3][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(\p8div.sa.div.b[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0498_ (.A(\p8div.sa.div.b[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0499_ (.A(\p8div.sa.div.b[2][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(\p8div.sa.div.b[2][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(\p8div.sa.div.b[2][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(\p8div.sa.div.b[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\p8div.sa.div.b[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(\p8div.sa.div.b[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(\p8div.sa.div.b[1][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(\p8div.sa.div.b[1][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0507_ (.A(\p8div.sa.div.b[1][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(\p8div.sa.div.b[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(\p8div.sa.div.b[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(\p8div.sa.div.b[0][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(\p8div.sa.div.b[0][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(\p8div.sa.div.b[0][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(\p8div.sa.div.b[0][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(\p8div.sa.div.b[0][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(\p8div.sa.div.b[0][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0516_ (.A(\p8div.sa.div.b[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(\p8div.sa.div.b[9][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0518_ (.A(\p8div.sa.div.b[9][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0519_ (.A(\p8div.sa.div.b[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(\p8div.sa.div.b[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(\p8div.sa.div.b[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(net441),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(\p8div.sa.div.b[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(\p8div.sa.div.b[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(\p8div.sa.div.b[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(\p8div.sa.div.b[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(\p8div.sa.div.b[6][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(\p8div.sa.div.b[6][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(\p8div.sa.div.b[5][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\p8div.sa.div.b[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(\p8div.sa.div.b[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(\p8div.sa.div.b[5][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(\p8div.sa.div.b[5][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0536_ (.A(\p8div.sa.div.b[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(\p8div.sa.div.b[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\p8div.sa.div.b[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(\p8div.sa.div.b[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(\p8div.sa.div.b[7][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(\p8div.sa.div.b[7][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(\p8div.sa.div.b[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0543_ (.A(\p8div.sa.div.b[8][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(\p8div.sa.div.b[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(\p8div.sa.div.b[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(\p8div.sa.div.b[8][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(\p8div.sa.div.b[8][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(\p8div.sa.div.b[4][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ));
 sky130_fd_sc_hd__inv_2 _0549_ (.A(\p8div.sa.div.b[10][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(\p8div.sa.div.acc[10][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(\p8div.sa.div.acc[10][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0070_));
 sky130_fd_sc_hd__o21a_1 _0552_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__a221o_1 _0553_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .C1(_0071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__o221a_1 _0554_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .C1(_0072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__a221o_1 _0555_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__o221a_1 _0556_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .C1(_0074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__or2_1 _0557_ (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .B(_0075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__a21o_2 _0558_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(_0076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[5].div_n.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(\p8div.sa.div.genblk1[5].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0077_));
 sky130_fd_sc_hd__o21a_1 _0560_ (.A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_1 _0561_ (.A(\p8div.sa.div.b[3][0] ),
    .B(\p8div.sa.div.b[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0079_));
 sky130_fd_sc_hd__a211o_1 _0562_ (.A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B1(_0078_),
    .C1(_0079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__o221a_1 _0563_ (.A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .C1(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__a221o_1 _0564_ (.A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__o22a_1 _0565_ (.A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__a221o_2 _0566_ (.A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(_0082_),
    .B2(_0083_),
    .C1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[4].div_n.a_ge_b ));
 sky130_fd_sc_hd__o21a_1 _0567_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__a221o_1 _0568_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .C1(_0084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__o221a_1 _0569_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .C1(_0085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__a221o_1 _0570_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__o221a_1 _0571_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .C1(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__or2_1 _0572_ (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .B(_0088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_2 _0573_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[3].div_n.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(\p8div.sa.div.genblk1[3].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0090_));
 sky130_fd_sc_hd__o21a_1 _0575_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__a221o_1 _0576_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .C1(_0091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__o221a_1 _0577_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .C1(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__a221o_1 _0578_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__o221a_1 _0579_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .C1(_0094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__or2_1 _0580_ (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .B(_0095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__a21o_2 _0581_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(_0096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[2].div_n.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(\p8div.sa.div.genblk1[2].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0097_));
 sky130_fd_sc_hd__o21a_1 _0583_ (.A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__a221o_1 _0584_ (.A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .C1(_0098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__o221a_1 _0585_ (.A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .C1(_0099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__a221o_1 _0586_ (.A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__o22a_1 _0587_ (.A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__a221o_2 _0588_ (.A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(_0101_),
    .B2(_0102_),
    .C1(net440),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[1].div_n.a_ge_b ));
 sky130_fd_sc_hd__o21a_1 _0589_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__nor2_1 _0590_ (.A(\p8div.sa.div.b[9][0] ),
    .B(\p8div.sa.div.b[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0104_));
 sky130_fd_sc_hd__a211o_1 _0591_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B1(_0103_),
    .C1(_0104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__o221a_1 _0592_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .C1(_0105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__a221o_1 _0593_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__o221a_1 _0594_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .C1(_0107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__or2_1 _0595_ (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .B(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__a21o_2 _0596_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B1(_0109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[10].div_n.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0597_ (.A(\p8div.sa.div.genblk1[10].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0110_));
 sky130_fd_sc_hd__or2_1 _0598_ (.A(_0066_),
    .B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _0599_ (.A(_0066_),
    .B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0112_));
 sky130_fd_sc_hd__nand2_1 _0600_ (.A(_0111_),
    .B(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0113_));
 sky130_fd_sc_hd__and2_1 _0601_ (.A(net39),
    .B(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.B_decode.F[0] ));
 sky130_fd_sc_hd__nand2b_1 _0602_ (.A_N(net7),
    .B(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0114_));
 sky130_fd_sc_hd__nand2b_1 _0603_ (.A_N(net8),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0115_));
 sky130_fd_sc_hd__nand2_2 _0604_ (.A(_0114_),
    .B(_0115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0116_));
 sky130_fd_sc_hd__nand3b_1 _0605_ (.A_N(net6),
    .B(net7),
    .C(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0117_));
 sky130_fd_sc_hd__nor2_1 _0606_ (.A(net8),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0118_));
 sky130_fd_sc_hd__nand2_1 _0607_ (.A(net6),
    .B(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_1 _0608_ (.A(_0117_),
    .B(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0120_));
 sky130_fd_sc_hd__a22o_1 _0609_ (.A1(net32),
    .A2(_0116_),
    .B1(_0120_),
    .B2(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__and3_1 _0610_ (.A(net33),
    .B(net29),
    .C(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0122_));
 sky130_fd_sc_hd__xor2_2 _0611_ (.A(_0121_),
    .B(_0122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__or3b_1 _0612_ (.A(_0066_),
    .B(net14),
    .C_N(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_1 _0613_ (.A(net15),
    .B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2_1 _0614_ (.A(net14),
    .B(_0124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0125_));
 sky130_fd_sc_hd__nand2_1 _0615_ (.A(_0123_),
    .B(_0125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0126_));
 sky130_fd_sc_hd__a22o_1 _0616_ (.A1(net38),
    .A2(_0113_),
    .B1(_0126_),
    .B2(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__nand2_1 _0617_ (.A(net39),
    .B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0128_));
 sky130_fd_sc_hd__and3_1 _0618_ (.A(net39),
    .B(net35),
    .C(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__xnor2_2 _0619_ (.A(_0127_),
    .B(_0129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0620_ (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.B_decode.F[1] ));
 sky130_fd_sc_hd__or4b_1 _0621_ (.A(net8),
    .B(net7),
    .C(net6),
    .D_N(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__and3_1 _0622_ (.A(net8),
    .B(net7),
    .C(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__nand3_1 _0623_ (.A(net8),
    .B(net7),
    .C(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0132_));
 sky130_fd_sc_hd__or2_1 _0624_ (.A(net31),
    .B(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__nand2_1 _0625_ (.A(_0130_),
    .B(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0134_));
 sky130_fd_sc_hd__a22o_1 _0626_ (.A1(net31),
    .A2(_0116_),
    .B1(_0120_),
    .B2(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__and3b_1 _0627_ (.A_N(net4),
    .B(net31),
    .C(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__nor2_1 _0628_ (.A(net31),
    .B(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0137_));
 sky130_fd_sc_hd__or2_1 _0629_ (.A(net31),
    .B(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__and3_1 _0630_ (.A(net4),
    .B(_0118_),
    .C(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__or2_1 _0631_ (.A(_0136_),
    .B(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _0632_ (.A1(net32),
    .A2(_0134_),
    .B1(_0140_),
    .B2(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__or2_1 _0633_ (.A(_0135_),
    .B(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__a22o_1 _0634_ (.A1(net32),
    .A2(_0120_),
    .B1(_0134_),
    .B2(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__a21oi_2 _0635_ (.A1(net4),
    .A2(_0116_),
    .B1(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0144_));
 sky130_fd_sc_hd__and2_1 _0636_ (.A(net33),
    .B(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__or3b_1 _0637_ (.A(_0121_),
    .B(_0145_),
    .C_N(_0144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__nand2_1 _0638_ (.A(net29),
    .B(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0147_));
 sky130_fd_sc_hd__xnor2_2 _0639_ (.A(_0142_),
    .B(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__or4b_1 _0640_ (.A(net15),
    .B(net16),
    .C(net14),
    .D_N(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__and3_1 _0641_ (.A(net15),
    .B(net16),
    .C(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__nand2b_1 _0642_ (.A_N(net36),
    .B(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0150_));
 sky130_fd_sc_hd__nand2_1 _0643_ (.A(_0148_),
    .B(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0151_));
 sky130_fd_sc_hd__and3b_1 _0644_ (.A_N(net37),
    .B(net36),
    .C(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__nor2_1 _0645_ (.A(net36),
    .B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0153_));
 sky130_fd_sc_hd__and3_1 _0646_ (.A(net37),
    .B(_0124_),
    .C(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__o21a_1 _0647_ (.A1(_0152_),
    .A2(_0154_),
    .B1(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__a221o_1 _0648_ (.A1(net36),
    .A2(_0113_),
    .B1(_0126_),
    .B2(net37),
    .C1(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__a21o_1 _0649_ (.A1(net38),
    .A2(_0151_),
    .B1(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_1 _0650_ (.A1(net38),
    .A2(_0126_),
    .B1(_0151_),
    .B2(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0158_));
 sky130_fd_sc_hd__a21oi_1 _0651_ (.A1(net37),
    .A2(_0113_),
    .B1(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0159_));
 sky130_fd_sc_hd__or3b_2 _0652_ (.A(\p8div.B_decode.F[0] ),
    .B(_0127_),
    .C_N(_0159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _0653_ (.A(net35),
    .B(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0161_));
 sky130_fd_sc_hd__xor2_2 _0654_ (.A(_0157_),
    .B(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.B_decode.F[3] ));
 sky130_fd_sc_hd__o21a_1 _0656_ (.A1(\p8div.B_decode.F[0] ),
    .A2(_0127_),
    .B1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__xnor2_1 _0657_ (.A(_0159_),
    .B(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.B_decode.F[2] ));
 sky130_fd_sc_hd__inv_2 _0658_ (.A(\p8div.B_decode.F[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__and4b_1 _0659_ (.A_N(net4),
    .B(_0118_),
    .C(_0137_),
    .D(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _0660_ (.A(net4),
    .B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__nand2_1 _0661_ (.A(net6),
    .B(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0165_));
 sky130_fd_sc_hd__and2_1 _0662_ (.A(_0131_),
    .B(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__and2b_1 _0663_ (.A_N(net32),
    .B(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__o21a_1 _0664_ (.A1(_0163_),
    .A2(_0167_),
    .B1(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _0665_ (.A1(net31),
    .A2(_0120_),
    .B1(_0134_),
    .B2(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__a221o_1 _0666_ (.A1(net6),
    .A2(_0116_),
    .B1(_0140_),
    .B2(net32),
    .C1(_0169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__or2_1 _0667_ (.A(_0168_),
    .B(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__o21ai_1 _0668_ (.A1(_0142_),
    .A2(_0146_),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0172_));
 sky130_fd_sc_hd__xnor2_2 _0669_ (.A(_0171_),
    .B(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__and4b_1 _0670_ (.A_N(net37),
    .B(_0124_),
    .C(_0153_),
    .D(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__and3_1 _0671_ (.A(net37),
    .B(net13),
    .C(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__nand3_1 _0672_ (.A(net12),
    .B(net13),
    .C(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0175_));
 sky130_fd_sc_hd__o21bai_1 _0673_ (.A1(net38),
    .A2(_0175_),
    .B1_N(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0176_));
 sky130_fd_sc_hd__a22o_1 _0674_ (.A1(net36),
    .A2(_0126_),
    .B1(_0151_),
    .B2(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__o21a_1 _0675_ (.A1(_0152_),
    .A2(_0154_),
    .B1(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0178_));
 sky130_fd_sc_hd__a211o_1 _0676_ (.A1(net14),
    .A2(_0113_),
    .B1(_0177_),
    .C1(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__a21o_1 _0677_ (.A1(net39),
    .A2(_0176_),
    .B1(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__o21a_1 _0678_ (.A1(_0157_),
    .A2(_0160_),
    .B1(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__xnor2_2 _0679_ (.A(_0180_),
    .B(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.B_decode.F[4] ));
 sky130_fd_sc_hd__o21a_1 _0681_ (.A1(_0121_),
    .A2(_0145_),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__xnor2_2 _0682_ (.A(_0144_),
    .B(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__nand2b_1 _0683_ (.A_N(_0145_),
    .B(\p8div.B_decode.F[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ));
 sky130_fd_sc_hd__or2_1 _0684_ (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__a21o_1 _0685_ (.A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ),
    .B1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__o211a_1 _0686_ (.A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(_0183_),
    .C1(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__a221o_1 _0687_ (.A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .C1(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__o221a_1 _0688_ (.A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .C1(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_2 _0689_ (.A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B1(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.div_0.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(\p8div.sa.div.div_0.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0188_));
 sky130_fd_sc_hd__o21a_1 _0691_ (.A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__nor2_1 _0692_ (.A(\p8div.sa.div.b[6][0] ),
    .B(\p8div.sa.div.b[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0190_));
 sky130_fd_sc_hd__a211o_1 _0693_ (.A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(_0189_),
    .C1(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__o221a_1 _0694_ (.A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0192_));
 sky130_fd_sc_hd__a221o_1 _0695_ (.A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .C1(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__o22a_1 _0696_ (.A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0194_));
 sky130_fd_sc_hd__a221o_2 _0697_ (.A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B1(_0193_),
    .B2(_0194_),
    .C1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[7].div_n.a_ge_b ));
 sky130_fd_sc_hd__o21a_1 _0698_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__a221o_1 _0699_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .C1(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__o221a_1 _0700_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__a221o_1 _0701_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .C1(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__o221a_1 _0702_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .C1(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__or2_1 _0703_ (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .B(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__a21o_2 _0704_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B1(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[6].div_n.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(\p8div.sa.div.genblk1[6].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0201_));
 sky130_fd_sc_hd__o21a_1 _0706_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__nor2_1 _0707_ (.A(\p8div.sa.div.b[7][0] ),
    .B(\p8div.sa.div.b[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0203_));
 sky130_fd_sc_hd__a211o_1 _0708_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(_0202_),
    .C1(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__o221a_1 _0709_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__a221o_1 _0710_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .C1(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__o221a_1 _0711_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .C1(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0207_));
 sky130_fd_sc_hd__or2_1 _0712_ (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .B(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__a21o_2 _0713_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B1(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[8].div_n.a_ge_b ));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(\p8div.sa.div.genblk1[8].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0209_));
 sky130_fd_sc_hd__o21a_1 _0715_ (.A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0210_));
 sky130_fd_sc_hd__a221o_1 _0716_ (.A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .A2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .B1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .C1(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__o221a_1 _0717_ (.A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .C1(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__a221o_1 _0718_ (.A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .C1(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__o22a_1 _0719_ (.A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .B2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__a221o_2 _0720_ (.A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .A2(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B1(_0213_),
    .B2(_0214_),
    .C1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.div.genblk1[9].div_n.a_ge_b ));
 sky130_fd_sc_hd__nor2_1 _0721_ (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0006_));
 sky130_fd_sc_hd__mux2_1 _0722_ (.A0(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[10].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[10].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0724_ (.A0(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[10].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0725_ (.A0(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[10].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__o22a_1 _0726_ (.A1(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(_0109_),
    .B1(_0110_),
    .B2(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(net427),
    .B(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0731_ (.A0(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__nor2_1 _0733_ (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0054_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[8].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[8].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[8].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0737_ (.A0(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[8].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__o22a_1 _0738_ (.A1(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(_0208_),
    .B1(_0209_),
    .B2(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _0739_ (.A(\p8div.sa.div.b[6][0] ),
    .B(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__nor2_1 _0745_ (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0042_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[6].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0747_ (.A0(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[6].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[6].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0749_ (.A0(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[6].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__o22a_1 _0750_ (.A1(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(_0200_),
    .B1(_0201_),
    .B2(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__nor2_1 _0751_ (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B(_0077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0036_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[5].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0753_ (.A0(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[5].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0754_ (.A0(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[5].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[5].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__o22a_1 _0756_ (.A1(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _0757_ (.A(\p8div.sa.div.b[3][0] ),
    .B(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0759_ (.A0(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _0763_ (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0024_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[3].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[3].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0766_ (.A0(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[3].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[3].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__o22a_1 _0768_ (.A1(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(_0089_),
    .B1(_0090_),
    .B2(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _0769_ (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .B(_0097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0018_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[2].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[2].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[2].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[2].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__o22a_1 _0774_ (.A1(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A2(_0096_),
    .B1(_0097_),
    .B2(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(net419),
    .B(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .A1(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .S(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0017_));
 sky130_fd_sc_hd__nand2_1 _0781_ (.A(\p8div.B_decode.F[0] ),
    .B(\p8div.sa.div.div_0.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0215_));
 sky130_fd_sc_hd__xnor2_1 _0782_ (.A(_0145_),
    .B(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0000_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .S(\p8div.sa.div.div_0.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .S(\p8div.sa.div.div_0.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .S(\p8div.sa.div.div_0.a_ge_b ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0003_));
 sky130_fd_sc_hd__o22a_1 _0786_ (.A1(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__or2_1 _0787_ (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ),
    .B(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0005_));
 sky130_fd_sc_hd__or4_1 _0788_ (.A(\p8div.a_piped[1] ),
    .B(\p8div.a_piped[0] ),
    .C(\p8div.a_piped[3] ),
    .D(\p8div.a_piped[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__nor4_1 _0789_ (.A(\p8div.a_piped[5] ),
    .B(\p8div.a_piped[4] ),
    .C(\p8div.a_piped[6] ),
    .D(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0217_));
 sky130_fd_sc_hd__or4_1 _0790_ (.A(\p8div.b_piped[1] ),
    .B(\p8div.b_piped[0] ),
    .C(\p8div.b_piped[3] ),
    .D(\p8div.b_piped[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__nor4_1 _0791_ (.A(\p8div.b_piped[5] ),
    .B(\p8div.b_piped[4] ),
    .C(\p8div.b_piped[6] ),
    .D(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0219_));
 sky130_fd_sc_hd__or2_2 _0792_ (.A(net22),
    .B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__or4_4 _0793_ (.A(net28),
    .B(\p8div.c_scale[0] ),
    .C(\p8div.c_scale[1] ),
    .D(\p8div.c_scale[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__o21ai_1 _0794_ (.A1(\p8div.c_scale[3] ),
    .A2(_0221_),
    .B1(\p8div.c_scale[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0222_));
 sky130_fd_sc_hd__or3_1 _0795_ (.A(\p8div.c_scale[3] ),
    .B(\p8div.c_scale[4] ),
    .C(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_2 _0796_ (.A(_0222_),
    .B(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0224_));
 sky130_fd_sc_hd__or3_1 _0797_ (.A(net28),
    .B(\p8div.c_scale[0] ),
    .C(\p8div.c_scale[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__a21boi_1 _0798_ (.A1(\p8div.c_scale[2] ),
    .A2(_0225_),
    .B1_N(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0226_));
 sky130_fd_sc_hd__a21bo_1 _0799_ (.A1(\p8div.c_scale[2] ),
    .A2(_0225_),
    .B1_N(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__xor2_1 _0800_ (.A(\p8div.c_scale[3] ),
    .B(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__xnor2_4 _0801_ (.A(\p8div.c_scale[3] ),
    .B(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0229_));
 sky130_fd_sc_hd__a211o_4 _0802_ (.A1(_0222_),
    .A2(_0223_),
    .B1(_0226_),
    .C1(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__xor2_4 _0803_ (.A(net28),
    .B(\p8div.c_scale[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__nand2b_2 _0804_ (.A_N(\p8div.c_scale[1] ),
    .B(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0232_));
 sky130_fd_sc_hd__o21ai_1 _0805_ (.A1(\p8div.c_decoded[11] ),
    .A2(\p8div.c_scale[0] ),
    .B1(\p8div.c_scale[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _0806_ (.A(_0225_),
    .B(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0234_));
 sky130_fd_sc_hd__a21o_2 _0807_ (.A1(_0225_),
    .A2(_0233_),
    .B1(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0236_));
 sky130_fd_sc_hd__or3_4 _0809_ (.A(\p8div.c_scale[3] ),
    .B(\p8div.c_scale[4] ),
    .C(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__o22ai_4 _0810_ (.A1(_0230_),
    .A2(_0232_),
    .B1(_0235_),
    .B2(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_1 _0811_ (.A(\p8div.c_scale[4] ),
    .B(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0239_));
 sky130_fd_sc_hd__nor2_1 _0812_ (.A(_0231_),
    .B(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0240_));
 sky130_fd_sc_hd__or2_2 _0813_ (.A(_0231_),
    .B(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _0814_ (.A(_0227_),
    .B(_0239_),
    .C(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _0815_ (.A(\p8div.c_scale[3] ),
    .B(\p8div.c_scale[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_2 _0816_ (.A(\p8div.c_scale[1] ),
    .B(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0244_));
 sky130_fd_sc_hd__nor3_1 _0817_ (.A(_0227_),
    .B(_0243_),
    .C(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0245_));
 sky130_fd_sc_hd__a31o_2 _0818_ (.A1(_0227_),
    .A2(_0239_),
    .A3(_0240_),
    .B1(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_4 _0819_ (.A0(\p8div.c_decoded[5] ),
    .A1(\p8div.c_decoded[6] ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__o22a_1 _0820_ (.A1(_0069_),
    .A2(\p8div.sa.div.b[10][4] ),
    .B1(_0070_),
    .B2(\p8div.sa.div.b[10][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0248_));
 sky130_fd_sc_hd__a21bo_1 _0821_ (.A1(\p8div.sa.div.b[10][1] ),
    .A2(\p8div.sa.div.b[10][0] ),
    .B1_N(\p8div.sa.div.acc[10][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _0822_ (.A(\p8div.sa.div.b[10][1] ),
    .B(\p8div.sa.div.b[10][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__nand2b_1 _0823_ (.A_N(\p8div.sa.div.b[10][2] ),
    .B(\p8div.sa.div.acc[10][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0251_));
 sky130_fd_sc_hd__and2b_1 _0824_ (.A_N(\p8div.sa.div.acc[10][2] ),
    .B(\p8div.sa.div.b[10][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__and2b_1 _0825_ (.A_N(\p8div.sa.div.acc[10][1] ),
    .B(\p8div.sa.div.b[10][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__a311o_1 _0826_ (.A1(_0249_),
    .A2(_0250_),
    .A3(_0251_),
    .B1(_0252_),
    .C1(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__nor2_1 _0827_ (.A(\p8div.sa.div.acc[10][4] ),
    .B(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0255_));
 sky130_fd_sc_hd__a221o_1 _0828_ (.A1(_0069_),
    .A2(\p8div.sa.div.b[10][4] ),
    .B1(_0248_),
    .B2(_0254_),
    .C1(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__or4_1 _0829_ (.A(\p8div.sa.div.acc[10][5] ),
    .B(\p8div.c_decoded[1] ),
    .C(\p8div.c_decoded[2] ),
    .D(\p8div.c_decoded[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__a221oi_1 _0830_ (.A1(net28),
    .A2(\p8div.c_decoded[4] ),
    .B1(\p8div.sa.div.acc[10][4] ),
    .B2(_0068_),
    .C1(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0258_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(\p8div.c_decoded[4] ),
    .A1(\p8div.c_decoded[5] ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(\p8div.c_decoded[6] ),
    .A1(\p8div.c_decoded[7] ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _0833_ (.A(_0259_),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0261_));
 sky130_fd_sc_hd__nand3_1 _0834_ (.A(_0256_),
    .B(_0258_),
    .C(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0262_));
 sky130_fd_sc_hd__o22ai_2 _0835_ (.A1(_0238_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0263_));
 sky130_fd_sc_hd__nand3b_1 _0836_ (.A_N(_0247_),
    .B(_0256_),
    .C(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0264_));
 sky130_fd_sc_hd__o22ai_4 _0837_ (.A1(_0230_),
    .A2(_0241_),
    .B1(_0244_),
    .B2(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0265_));
 sky130_fd_sc_hd__o21ai_2 _0838_ (.A1(_0259_),
    .A2(_0264_),
    .B1(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0266_));
 sky130_fd_sc_hd__or3_1 _0839_ (.A(_0227_),
    .B(_0235_),
    .C(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__or4_1 _0840_ (.A(\p8div.c_scale[4] ),
    .B(_0226_),
    .C(_0229_),
    .D(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_2 _0841_ (.A(_0267_),
    .B(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0269_));
 sky130_fd_sc_hd__mux2_4 _0842_ (.A0(\p8div.c_decoded[9] ),
    .A1(\p8div.c_decoded[10] ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(_0270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0271_));
 sky130_fd_sc_hd__or4_1 _0844_ (.A(\p8div.sa.div.acc[10][3] ),
    .B(\p8div.sa.div.acc[10][2] ),
    .C(\p8div.sa.div.acc[10][1] ),
    .D(\p8div.sa.div.acc[10][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__or4_1 _0845_ (.A(\p8div.sa.div.acc[10][4] ),
    .B(\p8div.sa.div.acc[10][5] ),
    .C(_0245_),
    .D(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(\p8div.c_decoded[7] ),
    .A1(\p8div.c_decoded[8] ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _0847_ (.A0(\p8div.c_decoded[8] ),
    .A1(\p8div.c_decoded[9] ),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _0848_ (.A(net25),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__o31a_1 _0849_ (.A1(_0247_),
    .A2(_0262_),
    .A3(net26),
    .B1(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__or2_2 _0850_ (.A(_0230_),
    .B(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__o22ai_4 _0851_ (.A1(_0230_),
    .A2(_0235_),
    .B1(_0237_),
    .B2(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0279_));
 sky130_fd_sc_hd__o22a_1 _0852_ (.A1(_0237_),
    .A2(_0241_),
    .B1(_0244_),
    .B2(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__o22ai_4 _0853_ (.A1(_0237_),
    .A2(_0241_),
    .B1(_0244_),
    .B2(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0281_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(_0264_),
    .A2(_0279_),
    .B1(_0281_),
    .B2(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__a221o_1 _0855_ (.A1(_0265_),
    .A2(net25),
    .B1(_0276_),
    .B2(_0242_),
    .C1(_0273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(_0269_),
    .A2(_0270_),
    .B1(net24),
    .B2(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__nor4_1 _0857_ (.A(_0277_),
    .B(_0282_),
    .C(_0283_),
    .D(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0285_));
 sky130_fd_sc_hd__a22o_1 _0858_ (.A1(_0246_),
    .A2(_0270_),
    .B1(_0279_),
    .B2(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(net27),
    .A2(_0265_),
    .B1(_0281_),
    .B2(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _0860_ (.A(_0269_),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _0861_ (.A(_0238_),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0289_));
 sky130_fd_sc_hd__and4bb_1 _0862_ (.A_N(_0286_),
    .B_N(_0287_),
    .C(_0288_),
    .D(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__a31oi_4 _0863_ (.A1(_0263_),
    .A2(_0266_),
    .A3(net19),
    .B1(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0291_));
 sky130_fd_sc_hd__a31o_2 _0864_ (.A1(_0263_),
    .A2(_0266_),
    .A3(_0285_),
    .B1(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _0865_ (.A(_0279_),
    .B(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__and2_1 _0866_ (.A(_0247_),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__and2_1 _0867_ (.A(net25),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__nand2_1 _0868_ (.A(net25),
    .B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0296_));
 sky130_fd_sc_hd__nand2_1 _0869_ (.A(_0294_),
    .B(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _0870_ (.A(_0271_),
    .B(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0298_));
 sky130_fd_sc_hd__a21o_1 _0871_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__or2_1 _0872_ (.A(_0238_),
    .B(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__a32o_1 _0873_ (.A1(_0270_),
    .A2(_0295_),
    .A3(_0300_),
    .B1(_0298_),
    .B2(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__nor2_1 _0874_ (.A(_0299_),
    .B(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0302_));
 sky130_fd_sc_hd__or2_2 _0875_ (.A(_0299_),
    .B(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__nand2_4 _0876_ (.A(_0291_),
    .B(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(_0247_),
    .B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0305_));
 sky130_fd_sc_hd__and3_1 _0878_ (.A(_0247_),
    .B(_0259_),
    .C(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _0879_ (.A(_0261_),
    .B(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__or3b_1 _0880_ (.A(_0307_),
    .B(_0306_),
    .C_N(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__nand2b_1 _0881_ (.A_N(net27),
    .B(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0309_));
 sky130_fd_sc_hd__o311a_1 _0882_ (.A1(_0280_),
    .A2(_0294_),
    .A3(_0305_),
    .B1(_0308_),
    .C1(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(_0246_),
    .B(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__o31ai_1 _0884_ (.A1(_0238_),
    .A2(_0292_),
    .A3(_0311_),
    .B1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0312_));
 sky130_fd_sc_hd__o21ai_1 _0885_ (.A1(_0292_),
    .A2(_0310_),
    .B1(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0291_),
    .B(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0314_));
 sky130_fd_sc_hd__xnor2_1 _0887_ (.A(_0247_),
    .B(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0315_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(_0313_),
    .A1(_0315_),
    .S(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__a21oi_2 _0889_ (.A1(_0291_),
    .A2(_0303_),
    .B1(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0317_));
 sky130_fd_sc_hd__and4_2 _0890_ (.A(_0241_),
    .B(_0244_),
    .C(_0291_),
    .D(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__or3b_2 _0891_ (.A(_0302_),
    .B(_0292_),
    .C_N(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _0892_ (.A1(_0291_),
    .A2(_0303_),
    .B1(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__a211oi_1 _0893_ (.A1(_0319_),
    .A2(_0320_),
    .B1(_0317_),
    .C1(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0321_));
 sky130_fd_sc_hd__a211o_1 _0894_ (.A1(_0319_),
    .A2(_0320_),
    .B1(_0317_),
    .C1(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__o31a_1 _0895_ (.A1(_0278_),
    .A2(_0292_),
    .A3(_0302_),
    .B1(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__o31ai_1 _0896_ (.A1(_0278_),
    .A2(_0292_),
    .A3(_0302_),
    .B1(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0324_));
 sky130_fd_sc_hd__a31o_2 _0897_ (.A1(_0236_),
    .A2(_0291_),
    .A3(_0303_),
    .B1(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _0898_ (.A(_0323_),
    .B(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0326_));
 sky130_fd_sc_hd__o21a_1 _0899_ (.A1(_0278_),
    .A2(_0304_),
    .B1(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__o31ai_1 _0900_ (.A1(_0278_),
    .A2(_0292_),
    .A3(_0302_),
    .B1(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0328_));
 sky130_fd_sc_hd__and3_1 _0901_ (.A(_0224_),
    .B(_0323_),
    .C(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _0902_ (.A(_0321_),
    .B(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0330_));
 sky130_fd_sc_hd__o21ai_1 _0903_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0331_));
 sky130_fd_sc_hd__o221a_1 _0904_ (.A1(_0278_),
    .A2(_0304_),
    .B1(_0325_),
    .B2(_0229_),
    .C1(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__and3_1 _0905_ (.A(_0228_),
    .B(_0325_),
    .C(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__a2bb2oi_2 _0906_ (.A1_N(_0317_),
    .A2_N(_0318_),
    .B1(_0319_),
    .B2(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0334_));
 sky130_fd_sc_hd__a22o_1 _0907_ (.A1(_0331_),
    .A2(_0332_),
    .B1(_0333_),
    .B2(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__o211a_1 _0908_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0319_),
    .C1(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_1 _0909_ (.A(_0333_),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0337_));
 sky130_fd_sc_hd__o32ai_4 _0910_ (.A1(_0224_),
    .A2(_0229_),
    .A3(_0325_),
    .B1(_0304_),
    .B2(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0338_));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(_0321_),
    .B(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _0912_ (.A1(_0333_),
    .A2(_0336_),
    .B1(_0338_),
    .B2(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _0913_ (.A(_0335_),
    .B(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__and4bb_1 _0914_ (.A_N(_0317_),
    .B_N(_0318_),
    .C(_0319_),
    .D(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(_0338_),
    .B(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0343_));
 sky130_fd_sc_hd__o21a_1 _0916_ (.A1(_0334_),
    .A2(_0342_),
    .B1(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__or4_1 _0917_ (.A(_0327_),
    .B(_0335_),
    .C(_0340_),
    .D(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__a21boi_1 _0918_ (.A1(_0330_),
    .A2(_0345_),
    .B1_N(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0346_));
 sky130_fd_sc_hd__and2_1 _0919_ (.A(_0329_),
    .B(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _0920_ (.A1(_0334_),
    .A2(_0338_),
    .B1(_0342_),
    .B2(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__xor2_1 _0921_ (.A(_0260_),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__o21a_1 _0922_ (.A1(_0292_),
    .A2(_0349_),
    .B1(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__o21a_1 _0923_ (.A1(_0238_),
    .A2(_0293_),
    .B1(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__nor3_1 _0924_ (.A(_0269_),
    .B(_0293_),
    .C(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0352_));
 sky130_fd_sc_hd__and2b_1 _0925_ (.A_N(_0246_),
    .B(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__o21ai_1 _0926_ (.A1(net25),
    .A2(_0294_),
    .B1(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0354_));
 sky130_fd_sc_hd__a21oi_1 _0927_ (.A1(net25),
    .A2(_0294_),
    .B1(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0355_));
 sky130_fd_sc_hd__o21ai_1 _0928_ (.A1(net25),
    .A2(_0306_),
    .B1(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0356_));
 sky130_fd_sc_hd__a21oi_1 _0929_ (.A1(net25),
    .A2(_0306_),
    .B1(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0357_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(_0238_),
    .A1(_0311_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__or4_1 _0931_ (.A(_0353_),
    .B(_0355_),
    .C(_0357_),
    .D(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__o32a_1 _0932_ (.A1(_0350_),
    .A2(_0351_),
    .A3(_0359_),
    .B1(_0291_),
    .B2(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(_0360_),
    .A1(_0313_),
    .S(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _0934_ (.A1(_0329_),
    .A2(_0334_),
    .B1(_0338_),
    .B2(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__a31o_1 _0935_ (.A1(_0247_),
    .A2(net27),
    .A3(net25),
    .B1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__and3_1 _0936_ (.A(_0281_),
    .B(_0297_),
    .C(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _0937_ (.A(net27),
    .B(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0365_));
 sky130_fd_sc_hd__a21o_1 _0938_ (.A1(net27),
    .A2(net25),
    .B1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__and3_1 _0939_ (.A(_0265_),
    .B(_0365_),
    .C(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__a311o_1 _0940_ (.A1(_0238_),
    .A2(_0276_),
    .A3(_0296_),
    .B1(_0364_),
    .C1(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_1 _0941_ (.A(_0246_),
    .B(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0369_));
 sky130_fd_sc_hd__o21ai_1 _0942_ (.A1(_0291_),
    .A2(_0352_),
    .B1(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0370_));
 sky130_fd_sc_hd__nand3_1 _0943_ (.A(net26),
    .B(net24),
    .C(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0371_));
 sky130_fd_sc_hd__a21o_1 _0944_ (.A1(net26),
    .A2(_0306_),
    .B1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__and3_1 _0945_ (.A(_0279_),
    .B(_0371_),
    .C(_0372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__a21oi_1 _0946_ (.A1(_0267_),
    .A2(_0268_),
    .B1(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0374_));
 sky130_fd_sc_hd__o31a_1 _0947_ (.A1(_0368_),
    .A2(_0373_),
    .A3(_0374_),
    .B1(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0375_));
 sky130_fd_sc_hd__a211o_1 _0948_ (.A1(_0275_),
    .A2(_0370_),
    .B1(_0375_),
    .C1(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(_0376_),
    .A1(_0360_),
    .S(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_1 _0950_ (.A1(_0348_),
    .A2(_0361_),
    .B1(_0362_),
    .B2(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(_0329_),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__or4_1 _0952_ (.A(net24),
    .B(_0293_),
    .C(_0300_),
    .D(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0380_));
 sky130_fd_sc_hd__o2111a_1 _0953_ (.A1(_0339_),
    .A2(_0379_),
    .B1(_0380_),
    .C1(_0376_),
    .D1(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__o211a_1 _0954_ (.A1(_0322_),
    .A2(_0324_),
    .B1(_0326_),
    .C1(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__a21oi_1 _0955_ (.A1(_0331_),
    .A2(_0332_),
    .B1(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0383_));
 sky130_fd_sc_hd__or4_1 _0956_ (.A(_0322_),
    .B(_0324_),
    .C(_0325_),
    .D(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__o21ai_1 _0957_ (.A1(_0270_),
    .A2(_0295_),
    .B1(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0385_));
 sky130_fd_sc_hd__a21oi_1 _0958_ (.A1(_0270_),
    .A2(_0295_),
    .B1(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0386_));
 sky130_fd_sc_hd__or2_1 _0959_ (.A(_0271_),
    .B(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _0960_ (.A(_0271_),
    .B(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0388_));
 sky130_fd_sc_hd__and3_1 _0961_ (.A(_0265_),
    .B(_0387_),
    .C(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__nor2_1 _0962_ (.A(_0386_),
    .B(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0390_));
 sky130_fd_sc_hd__xnor2_1 _0963_ (.A(_0270_),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _0964_ (.A(_0279_),
    .B(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0392_));
 sky130_fd_sc_hd__and2_1 _0965_ (.A(_0271_),
    .B(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__or3_1 _0966_ (.A(_0280_),
    .B(_0298_),
    .C(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__o2111a_1 _0967_ (.A1(_0270_),
    .A2(_0288_),
    .B1(_0390_),
    .C1(_0392_),
    .D1(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(_0271_),
    .A1(_0395_),
    .S(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__a21oi_1 _0969_ (.A1(_0337_),
    .A2(_0384_),
    .B1(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0397_));
 sky130_fd_sc_hd__or4b_1 _0970_ (.A(_0378_),
    .B(_0381_),
    .C(_0397_),
    .D_N(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _0971_ (.A(_0346_),
    .B(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__and2b_2 _0972_ (.A_N(_0220_),
    .B(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(_0355_),
    .B(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__or3b_1 _0974_ (.A(_0400_),
    .B(_0367_),
    .C_N(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__or3b_2 _0975_ (.A(_0335_),
    .B(_0401_),
    .C_N(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__a21oi_1 _0976_ (.A1(\p8div.d_sign ),
    .A2(_0399_),
    .B1(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0403_));
 sky130_fd_sc_hd__a31o_1 _0977_ (.A1(\p8div.d_sign ),
    .A2(_0399_),
    .A3(_0402_),
    .B1(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__nor2_4 _0978_ (.A(_0403_),
    .B(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uo_out[1]));
 sky130_fd_sc_hd__or3_1 _0979_ (.A(_0357_),
    .B(_0364_),
    .C(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__or3_2 _0980_ (.A(_0332_),
    .B(_0379_),
    .C(_0405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__or3_2 _0981_ (.A(_0346_),
    .B(_0398_),
    .C(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__a21oi_1 _0982_ (.A1(\p8div.d_sign ),
    .A2(_0407_),
    .B1(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0408_));
 sky130_fd_sc_hd__a31o_1 _0983_ (.A1(\p8div.d_sign ),
    .A2(_0406_),
    .A3(_0407_),
    .B1(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__nor2_4 _0984_ (.A(_0408_),
    .B(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uo_out[2]));
 sky130_fd_sc_hd__a21bo_1 _0985_ (.A1(_0329_),
    .A2(_0334_),
    .B1_N(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__or3_4 _0986_ (.A(_0341_),
    .B(_0373_),
    .C(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__o21a_1 _0987_ (.A1(_0406_),
    .A2(_0407_),
    .B1(\p8div.d_sign ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__o21bai_1 _0988_ (.A1(_0411_),
    .A2(_0412_),
    .B1_N(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0413_));
 sky130_fd_sc_hd__a21oi_4 _0989_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uo_out[3]));
 sky130_fd_sc_hd__or4bb_4 _0990_ (.A(_0347_),
    .B(_0341_),
    .C_N(_0343_),
    .D_N(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__o31a_1 _0991_ (.A1(_0406_),
    .A2(_0407_),
    .A3(_0411_),
    .B1(\p8div.d_sign ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__o21bai_1 _0992_ (.A1(_0414_),
    .A2(_0415_),
    .B1_N(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0416_));
 sky130_fd_sc_hd__a21oi_4 _0993_ (.A1(_0414_),
    .A2(_0415_),
    .B1(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uo_out[4]));
 sky130_fd_sc_hd__or3b_2 _0994_ (.A(_0341_),
    .B(_0344_),
    .C_N(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0418_));
 sky130_fd_sc_hd__o41ai_1 _0996_ (.A1(_0406_),
    .A2(_0407_),
    .A3(_0411_),
    .A4(_0414_),
    .B1(\p8div.d_sign ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0419_));
 sky130_fd_sc_hd__a21oi_1 _0997_ (.A1(_0418_),
    .A2(net18),
    .B1(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0420_));
 sky130_fd_sc_hd__o21a_2 _0998_ (.A1(_0418_),
    .A2(_0419_),
    .B1(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__nand2_1 _0999_ (.A(\p8div.d_sign ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0421_));
 sky130_fd_sc_hd__a21oi_1 _1000_ (.A1(net18),
    .A2(_0421_),
    .B1(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0422_));
 sky130_fd_sc_hd__a31o_1 _1001_ (.A1(_0327_),
    .A2(net18),
    .A3(_0421_),
    .B1(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__nor2_4 _1002_ (.A(_0422_),
    .B(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uo_out[6]));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(\p8div.d_sign ),
    .A1(\p8div.a_piped[7] ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__or2_4 _1004_ (.A(net20),
    .B(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__or4b_1 _1005_ (.A(net32),
    .B(net4),
    .C(net31),
    .D_N(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__nor2_1 _1006_ (.A(_0146_),
    .B(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0426_));
 sky130_fd_sc_hd__and3b_1 _1007_ (.A_N(net33),
    .B(_0166_),
    .C(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _1008_ (.A(_0117_),
    .B(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0428_));
 sky130_fd_sc_hd__o21a_1 _1009_ (.A1(_0427_),
    .A2(_0428_),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0429_));
 sky130_fd_sc_hd__o21ai_1 _1010_ (.A1(net32),
    .A2(net33),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0431_));
 sky130_fd_sc_hd__a21o_1 _1012_ (.A1(net4),
    .A2(net29),
    .B1(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__a21o_1 _1013_ (.A1(net31),
    .A2(net30),
    .B1(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__o21a_1 _1014_ (.A1(_0132_),
    .A2(_0164_),
    .B1(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_1 _1015_ (.A(_0433_),
    .B(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0435_));
 sky130_fd_sc_hd__and2_1 _1016_ (.A(_0067_),
    .B(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__a31o_1 _1017_ (.A1(net32),
    .A2(net33),
    .A3(_0166_),
    .B1(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0437_));
 sky130_fd_sc_hd__a32o_1 _1018_ (.A1(net2),
    .A2(net29),
    .A3(_0167_),
    .B1(_0431_),
    .B2(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__a21oi_1 _1019_ (.A1(net30),
    .A2(_0138_),
    .B1(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0439_));
 sky130_fd_sc_hd__or2_1 _1020_ (.A(_0114_),
    .B(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0440_));
 sky130_fd_sc_hd__o21ai_1 _1021_ (.A1(net30),
    .A2(_0115_),
    .B1(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0441_));
 sky130_fd_sc_hd__or4_1 _1022_ (.A(_0435_),
    .B(_0437_),
    .C(_0438_),
    .D(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0442_));
 sky130_fd_sc_hd__or3_1 _1023_ (.A(_0426_),
    .B(_0429_),
    .C(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__o21a_1 _1024_ (.A1(_0163_),
    .A2(_0426_),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__a41o_1 _1025_ (.A1(net8),
    .A2(net7),
    .A3(net30),
    .A4(_0165_),
    .B1(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0444_));
 sky130_fd_sc_hd__a31o_1 _1026_ (.A1(_0067_),
    .A2(_0118_),
    .A3(_0138_),
    .B1(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__o21a_1 _1027_ (.A1(_0139_),
    .A2(_0166_),
    .B1(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__or3_1 _1028_ (.A(_0443_),
    .B(_0445_),
    .C(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__o21a_1 _1029_ (.A1(_0139_),
    .A2(_0426_),
    .B1(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0447_));
 sky130_fd_sc_hd__a2111o_2 _1030_ (.A1(net30),
    .A2(_0166_),
    .B1(_0436_),
    .C1(_0445_),
    .D1(_0447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__or4b_1 _1031_ (.A(net38),
    .B(net37),
    .C(net36),
    .D_N(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__o21bai_1 _1032_ (.A1(_0152_),
    .A2(_0173_),
    .B1_N(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0449_));
 sky130_fd_sc_hd__o31a_1 _1033_ (.A1(net38),
    .A2(net12),
    .A3(net10),
    .B1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0450_));
 sky130_fd_sc_hd__a21o_1 _1034_ (.A1(net13),
    .A2(net34),
    .B1(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__o221a_1 _1035_ (.A1(_0150_),
    .A2(_0450_),
    .B1(_0451_),
    .B2(_0125_),
    .C1(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0452_));
 sky130_fd_sc_hd__o21a_1 _1036_ (.A1(net36),
    .A2(net14),
    .B1(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__o21bai_1 _1037_ (.A1(_0450_),
    .A2(_0453_),
    .B1_N(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0454_));
 sky130_fd_sc_hd__o21a_1 _1038_ (.A1(net34),
    .A2(_0111_),
    .B1(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0455_));
 sky130_fd_sc_hd__o21ai_1 _1039_ (.A1(net38),
    .A2(net10),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2b_1 _1040_ (.A_N(_0456_),
    .B(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0457_));
 sky130_fd_sc_hd__o31a_1 _1041_ (.A1(net11),
    .A2(_0128_),
    .A3(_0175_),
    .B1(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0458_));
 sky130_fd_sc_hd__a21bo_1 _1042_ (.A1(_0123_),
    .A2(_0148_),
    .B1_N(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(net11),
    .B(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0460_));
 sky130_fd_sc_hd__a2bb2o_1 _1044_ (.A1_N(net39),
    .A2_N(net35),
    .B1(_0459_),
    .B2(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0461_));
 sky130_fd_sc_hd__and4_1 _1045_ (.A(_0452_),
    .B(_0455_),
    .C(_0458_),
    .D(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0462_));
 sky130_fd_sc_hd__o21a_1 _1046_ (.A1(_0160_),
    .A2(_0448_),
    .B1(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ));
 sky130_fd_sc_hd__o21bai_1 _1047_ (.A1(_0160_),
    .A2(_0448_),
    .B1_N(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(net34),
    .B(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0464_));
 sky130_fd_sc_hd__o41a_1 _1049_ (.A1(net15),
    .A2(net16),
    .A3(net34),
    .A4(_0153_),
    .B1(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0465_));
 sky130_fd_sc_hd__nand3_1 _1050_ (.A(net15),
    .B(net16),
    .C(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0466_));
 sky130_fd_sc_hd__a31o_1 _1051_ (.A1(net37),
    .A2(net36),
    .A3(net14),
    .B1(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0467_));
 sky130_fd_sc_hd__o21ai_1 _1052_ (.A1(_0154_),
    .A2(_0174_),
    .B1(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0468_));
 sky130_fd_sc_hd__and4_1 _1053_ (.A(_0464_),
    .B(_0465_),
    .C(_0467_),
    .D(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ));
 sky130_fd_sc_hd__nor2_1 _1054_ (.A(_0154_),
    .B(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0469_));
 sky130_fd_sc_hd__o211a_1 _1055_ (.A1(net34),
    .A2(_0469_),
    .B1(_0466_),
    .C1(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ));
 sky130_fd_sc_hd__a2bb2o_1 _1056_ (.A1_N(_0163_),
    .A2_N(_0427_),
    .B1(net2),
    .B2(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0470_));
 sky130_fd_sc_hd__nand2b_1 _1057_ (.A_N(_0115_),
    .B(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0471_));
 sky130_fd_sc_hd__mux2_1 _1058_ (.A0(_0130_),
    .A1(_0133_),
    .S(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1059_ (.A0(_0117_),
    .A1(_0119_),
    .S(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0473_));
 sky130_fd_sc_hd__and3_1 _1060_ (.A(_0440_),
    .B(_0470_),
    .C(_0471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0474_));
 sky130_fd_sc_hd__and3_1 _1061_ (.A(_0472_),
    .B(_0473_),
    .C(_0474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0475_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0476_));
 sky130_fd_sc_hd__a211o_1 _1063_ (.A1(_0136_),
    .A2(_0430_),
    .B1(_0438_),
    .C1(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(_0123_),
    .A1(_0125_),
    .S(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1065_ (.A0(_0148_),
    .A1(_0150_),
    .S(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0479_));
 sky130_fd_sc_hd__a22oi_1 _1066_ (.A1(_0128_),
    .A2(_0173_),
    .B1(_0456_),
    .B2(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0480_));
 sky130_fd_sc_hd__o31a_1 _1067_ (.A1(_0111_),
    .A2(_0450_),
    .A3(_0453_),
    .B1(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0481_));
 sky130_fd_sc_hd__and4_1 _1068_ (.A(_0458_),
    .B(_0479_),
    .C(_0480_),
    .D(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0482_));
 sky130_fd_sc_hd__o211a_1 _1069_ (.A1(net39),
    .A2(_0460_),
    .B1(_0478_),
    .C1(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0483_));
 sky130_fd_sc_hd__or2_1 _1070_ (.A(_0477_),
    .B(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ));
 sky130_fd_sc_hd__xnor2_1 _1071_ (.A(_0477_),
    .B(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_0_HCA.hca_stage_0.SUM ));
 sky130_fd_sc_hd__xor2_1 _1072_ (.A(net30),
    .B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\p8div.pipe_sign.A ));
 sky130_fd_sc_hd__dfrtp_1 _1073_ (.CLK(clknet_leaf_8_clk),
    .D(net10),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1074_ (.CLK(clknet_leaf_8_clk),
    .D(net38),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1075_ (.CLK(clknet_leaf_8_clk),
    .D(net37),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1076_ (.CLK(clknet_leaf_8_clk),
    .D(net36),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1077_ (.CLK(clknet_leaf_7_clk),
    .D(net14),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1078_ (.CLK(clknet_leaf_7_clk),
    .D(net15),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1079_ (.CLK(clknet_leaf_7_clk),
    .D(net16),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_leaf_13_clk),
    .D(net239),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_leaf_14_clk),
    .D(net319),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1082_ (.CLK(clknet_leaf_14_clk),
    .D(net197),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1083_ (.CLK(clknet_leaf_14_clk),
    .D(net224),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1084_ (.CLK(clknet_leaf_13_clk),
    .D(net198),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1085_ (.CLK(clknet_leaf_13_clk),
    .D(net231),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1086_ (.CLK(clknet_leaf_13_clk),
    .D(net210),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.b_piped[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_leaf_14_clk),
    .D(net259),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_leaf_14_clk),
    .D(net196),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1089_ (.CLK(clknet_leaf_14_clk),
    .D(net262),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_leaf_14_clk),
    .D(net364),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_leaf_13_clk),
    .D(net152),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1092_ (.CLK(clknet_leaf_14_clk),
    .D(net209),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_leaf_13_clk),
    .D(net247),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_leaf_14_clk),
    .D(net344),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_leaf_14_clk),
    .D(net241),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_leaf_14_clk),
    .D(net384),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_leaf_14_clk),
    .D(net366),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_leaf_14_clk),
    .D(net336),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_leaf_14_clk),
    .D(net281),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_leaf_14_clk),
    .D(net278),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_leaf_8_clk),
    .D(net254),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_leaf_8_clk),
    .D(net299),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_leaf_8_clk),
    .D(net170),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_leaf_8_clk),
    .D(net335),
    .RESET_B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_leaf_8_clk),
    .D(net137),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_leaf_7_clk),
    .D(net148),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_leaf_7_clk),
    .D(net156),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_leaf_14_clk),
    .D(net279),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_leaf_14_clk),
    .D(net300),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_leaf_15_clk),
    .D(net348),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_leaf_10_clk),
    .D(net172),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_leaf_12_clk),
    .D(net283),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_leaf_12_clk),
    .D(net261),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1114_ (.CLK(clknet_leaf_12_clk),
    .D(net214),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1115_ (.CLK(clknet_leaf_9_clk),
    .D(net166),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1116_ (.CLK(clknet_leaf_9_clk),
    .D(net178),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1117_ (.CLK(clknet_leaf_9_clk),
    .D(net182),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_leaf_9_clk),
    .D(net174),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_leaf_9_clk),
    .D(net204),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_leaf_10_clk),
    .D(net136),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_leaf_10_clk),
    .D(net131),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_leaf_14_clk),
    .D(net353),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_leaf_14_clk),
    .D(net324),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1124_ (.CLK(clknet_leaf_15_clk),
    .D(net119),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_leaf_9_clk),
    .D(net159),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_leaf_10_clk),
    .D(net296),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_leaf_10_clk),
    .D(net269),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_leaf_12_clk),
    .D(net203),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_leaf_10_clk),
    .D(net207),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_leaf_10_clk),
    .D(net153),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_leaf_9_clk),
    .D(net158),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_leaf_9_clk),
    .D(net352),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1133_ (.CLK(clknet_leaf_10_clk),
    .D(net235),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_leaf_10_clk),
    .D(net252),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_leaf_10_clk),
    .D(net275),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_leaf_9_clk),
    .D(net177),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_leaf_9_clk),
    .D(net175),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_leaf_8_clk),
    .D(net332),
    .RESET_B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_leaf_8_clk),
    .D(net258),
    .RESET_B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1140_ (.CLK(clknet_leaf_8_clk),
    .D(net161),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1141_ (.CLK(clknet_leaf_7_clk),
    .D(net238),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1142_ (.CLK(clknet_leaf_7_clk),
    .D(net146),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(clknet_leaf_10_clk),
    .D(net167),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(clknet_leaf_9_clk),
    .D(net267),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(clknet_leaf_9_clk),
    .D(net176),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1146_ (.CLK(clknet_leaf_9_clk),
    .D(net333),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(clknet_leaf_10_clk),
    .D(net155),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1148_ (.CLK(clknet_leaf_10_clk),
    .D(net187),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1149_ (.CLK(clknet_leaf_10_clk),
    .D(net213),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_B.a_q[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1150_ (.CLK(clknet_leaf_7_clk),
    .D(net2),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1151_ (.CLK(clknet_leaf_6_clk),
    .D(net3),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1152_ (.CLK(clknet_leaf_6_clk),
    .D(net4),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1153_ (.CLK(clknet_leaf_6_clk),
    .D(net5),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1154_ (.CLK(clknet_leaf_6_clk),
    .D(net6),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1155_ (.CLK(clknet_leaf_11_clk),
    .D(net7),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1156_ (.CLK(clknet_leaf_11_clk),
    .D(net8),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1157_ (.CLK(clknet_leaf_5_clk),
    .D(net30),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(clknet_leaf_13_clk),
    .D(net232),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(clknet_leaf_13_clk),
    .D(net363),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(clknet_leaf_13_clk),
    .D(net322),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(clknet_leaf_13_clk),
    .D(net349),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(clknet_leaf_13_clk),
    .D(net287),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(clknet_leaf_13_clk),
    .D(net308),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(clknet_leaf_13_clk),
    .D(net314),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1165_ (.CLK(clknet_leaf_11_clk),
    .D(net356),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.a_piped[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(clknet_leaf_13_clk),
    .D(net266),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(clknet_leaf_12_clk),
    .D(net191),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(clknet_leaf_12_clk),
    .D(net216),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(clknet_leaf_12_clk),
    .D(net264),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1170_ (.CLK(clknet_leaf_12_clk),
    .D(net240),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(clknet_leaf_13_clk),
    .D(net295),
    .RESET_B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1172_ (.CLK(clknet_leaf_13_clk),
    .D(net226),
    .RESET_B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1173_ (.CLK(clknet_leaf_6_clk),
    .D(net334),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1174_ (.CLK(clknet_leaf_12_clk),
    .D(net215),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1175_ (.CLK(clknet_leaf_12_clk),
    .D(net180),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(clknet_leaf_12_clk),
    .D(net188),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1177_ (.CLK(clknet_leaf_12_clk),
    .D(net173),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1178_ (.CLK(clknet_leaf_12_clk),
    .D(net151),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1179_ (.CLK(clknet_leaf_12_clk),
    .D(net205),
    .RESET_B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1180_ (.CLK(clknet_leaf_13_clk),
    .D(net234),
    .RESET_B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1181_ (.CLK(clknet_leaf_6_clk),
    .D(net223),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1182_ (.CLK(clknet_leaf_7_clk),
    .D(net201),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1183_ (.CLK(clknet_leaf_6_clk),
    .D(net243),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1184_ (.CLK(clknet_leaf_7_clk),
    .D(net378),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1185_ (.CLK(clknet_leaf_6_clk),
    .D(net225),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1186_ (.CLK(clknet_leaf_6_clk),
    .D(net326),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1187_ (.CLK(clknet_leaf_11_clk),
    .D(net162),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1188_ (.CLK(clknet_leaf_11_clk),
    .D(net168),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1189_ (.CLK(clknet_leaf_5_clk),
    .D(net249),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(clknet_leaf_12_clk),
    .D(net339),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(clknet_leaf_12_clk),
    .D(net217),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1192_ (.CLK(clknet_leaf_11_clk),
    .D(net306),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1193_ (.CLK(clknet_leaf_12_clk),
    .D(net219),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1194_ (.CLK(clknet_leaf_11_clk),
    .D(net160),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1195_ (.CLK(clknet_leaf_13_clk),
    .D(net276),
    .RESET_B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(clknet_leaf_13_clk),
    .D(net256),
    .RESET_B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1197_ (.CLK(clknet_leaf_6_clk),
    .D(net272),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1198_ (.CLK(clknet_leaf_7_clk),
    .D(net369),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1199_ (.CLK(clknet_leaf_7_clk),
    .D(net367),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_leaf_7_clk),
    .D(net368),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1201_ (.CLK(clknet_leaf_11_clk),
    .D(net365),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1202_ (.CLK(clknet_leaf_6_clk),
    .D(net220),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1203_ (.CLK(clknet_leaf_11_clk),
    .D(net358),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1204_ (.CLK(clknet_leaf_11_clk),
    .D(net165),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1205_ (.CLK(clknet_leaf_5_clk),
    .D(net265),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_leaf_11_clk),
    .D(net305),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1207_ (.CLK(clknet_leaf_11_clk),
    .D(net310),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1208_ (.CLK(clknet_leaf_10_clk),
    .D(net193),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1209_ (.CLK(clknet_leaf_11_clk),
    .D(net211),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1210_ (.CLK(clknet_leaf_11_clk),
    .D(net347),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1211_ (.CLK(clknet_leaf_12_clk),
    .D(net206),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(clknet_leaf_12_clk),
    .D(net263),
    .RESET_B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1213_ (.CLK(clknet_leaf_6_clk),
    .D(net228),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1214_ (.CLK(clknet_leaf_10_clk),
    .D(net189),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1215_ (.CLK(clknet_leaf_10_clk),
    .D(net186),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1216_ (.CLK(clknet_leaf_10_clk),
    .D(net202),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1217_ (.CLK(clknet_leaf_11_clk),
    .D(net285),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1218_ (.CLK(clknet_leaf_10_clk),
    .D(net184),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1219_ (.CLK(clknet_leaf_12_clk),
    .D(net312),
    .RESET_B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1220_ (.CLK(clknet_leaf_12_clk),
    .D(net171),
    .RESET_B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1221_ (.CLK(clknet_leaf_6_clk),
    .D(net115),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1222_ (.CLK(clknet_leaf_6_clk),
    .D(net120),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1223_ (.CLK(clknet_leaf_6_clk),
    .D(net230),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1224_ (.CLK(clknet_leaf_6_clk),
    .D(net123),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1225_ (.CLK(clknet_leaf_6_clk),
    .D(net327),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1226_ (.CLK(clknet_leaf_6_clk),
    .D(net309),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1227_ (.CLK(clknet_leaf_11_clk),
    .D(net218),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1228_ (.CLK(clknet_leaf_11_clk),
    .D(net302),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1229_ (.CLK(clknet_leaf_5_clk),
    .D(net303),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1230_ (.CLK(clknet_leaf_10_clk),
    .D(net133),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1231_ (.CLK(clknet_leaf_10_clk),
    .D(net134),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1232_ (.CLK(clknet_leaf_10_clk),
    .D(net126),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1233_ (.CLK(clknet_leaf_11_clk),
    .D(net271),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1234_ (.CLK(clknet_leaf_11_clk),
    .D(net359),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1235_ (.CLK(clknet_leaf_12_clk),
    .D(net145),
    .RESET_B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1236_ (.CLK(clknet_leaf_12_clk),
    .D(net212),
    .RESET_B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1237_ (.CLK(clknet_leaf_5_clk),
    .D(net150),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_A.a_q[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1238_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.sa.div.div_0.a_ge_b ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.Q_I ));
 sky130_fd_sc_hd__dfrtp_1 _1239_ (.CLK(clknet_leaf_5_clk),
    .D(\p8div.pipe_sign.A ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1240_ (.CLK(clknet_leaf_6_clk),
    .D(net246),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.d_sign ));
 sky130_fd_sc_hd__dfrtp_1 _1241_ (.CLK(clknet_leaf_6_clk),
    .D(net257),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1242_ (.CLK(clknet_leaf_6_clk),
    .D(net222),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1243_ (.CLK(clknet_leaf_5_clk),
    .D(net144),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1244_ (.CLK(clknet_leaf_6_clk),
    .D(net311),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1245_ (.CLK(clknet_leaf_5_clk),
    .D(net208),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1246_ (.CLK(clknet_leaf_6_clk),
    .D(net116),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1247_ (.CLK(clknet_leaf_5_clk),
    .D(net169),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1248_ (.CLK(clknet_leaf_5_clk),
    .D(net200),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1249_ (.CLK(clknet_leaf_5_clk),
    .D(net141),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.pipe_sign.a_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1250_ (.CLK(clknet_leaf_17_clk),
    .D(_0006_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.acc[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1251_ (.CLK(clknet_leaf_17_clk),
    .D(_0007_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.acc[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1252_ (.CLK(clknet_leaf_17_clk),
    .D(_0008_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.acc[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1253_ (.CLK(clknet_leaf_17_clk),
    .D(_0009_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.acc[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1254_ (.CLK(clknet_leaf_16_clk),
    .D(_0010_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.acc[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1255_ (.CLK(clknet_leaf_16_clk),
    .D(_0011_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.acc[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1256_ (.CLK(clknet_leaf_17_clk),
    .D(net433),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1257_ (.CLK(clknet_leaf_17_clk),
    .D(net432),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1258_ (.CLK(clknet_leaf_17_clk),
    .D(net405),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1259_ (.CLK(clknet_leaf_17_clk),
    .D(net409),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1260_ (.CLK(clknet_leaf_16_clk),
    .D(net426),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1261_ (.CLK(clknet_leaf_19_clk),
    .D(net395),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1262_ (.CLK(clknet_leaf_16_clk),
    .D(\p8div.sa.div.genblk1[10].div_n.a_ge_b ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1263_ (.CLK(clknet_leaf_16_clk),
    .D(net375),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1264_ (.CLK(clknet_leaf_16_clk),
    .D(net374),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1265_ (.CLK(clknet_leaf_16_clk),
    .D(net253),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1266_ (.CLK(clknet_leaf_16_clk),
    .D(net376),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1267_ (.CLK(clknet_leaf_15_clk),
    .D(net143),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1268_ (.CLK(clknet_leaf_15_clk),
    .D(net195),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1269_ (.CLK(clknet_leaf_15_clk),
    .D(net154),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1270_ (.CLK(clknet_leaf_15_clk),
    .D(net360),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1271_ (.CLK(clknet_leaf_15_clk),
    .D(net289),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1272_ (.CLK(clknet_leaf_15_clk),
    .D(net297),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_decoded[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1273_ (.CLK(clknet_leaf_17_clk),
    .D(_0060_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1274_ (.CLK(clknet_leaf_17_clk),
    .D(_0061_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1275_ (.CLK(clknet_leaf_17_clk),
    .D(_0062_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1276_ (.CLK(clknet_leaf_17_clk),
    .D(_0063_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1277_ (.CLK(clknet_leaf_17_clk),
    .D(_0064_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1278_ (.CLK(clknet_leaf_17_clk),
    .D(_0065_),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1279_ (.CLK(clknet_leaf_17_clk),
    .D(net427),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1280_ (.CLK(clknet_leaf_17_clk),
    .D(net397),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1281_ (.CLK(clknet_leaf_17_clk),
    .D(net406),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1282_ (.CLK(clknet_leaf_17_clk),
    .D(net412),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1283_ (.CLK(clknet_leaf_19_clk),
    .D(net413),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1284_ (.CLK(clknet_leaf_19_clk),
    .D(net410),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1285_ (.CLK(clknet_leaf_19_clk),
    .D(\p8div.sa.div.genblk1[9].div_n.a_ge_b ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1286_ (.CLK(clknet_leaf_19_clk),
    .D(net229),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1287_ (.CLK(clknet_leaf_16_clk),
    .D(net372),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1288_ (.CLK(clknet_leaf_19_clk),
    .D(net260),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1289_ (.CLK(clknet_leaf_20_clk),
    .D(net250),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1290_ (.CLK(clknet_leaf_20_clk),
    .D(net251),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1291_ (.CLK(clknet_leaf_20_clk),
    .D(net242),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1292_ (.CLK(clknet_leaf_15_clk),
    .D(net164),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1293_ (.CLK(clknet_leaf_15_clk),
    .D(net142),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1294_ (.CLK(clknet_leaf_15_clk),
    .D(net280),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[10].div_n.Q_I[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1295_ (.CLK(clknet_leaf_18_clk),
    .D(_0054_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1296_ (.CLK(clknet_leaf_18_clk),
    .D(_0055_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1297_ (.CLK(clknet_leaf_18_clk),
    .D(_0056_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1298_ (.CLK(clknet_leaf_19_clk),
    .D(_0057_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1299_ (.CLK(clknet_leaf_19_clk),
    .D(_0058_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1300_ (.CLK(clknet_leaf_19_clk),
    .D(_0059_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1301_ (.CLK(clknet_leaf_18_clk),
    .D(net431),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1302_ (.CLK(clknet_leaf_18_clk),
    .D(net435),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1303_ (.CLK(clknet_leaf_18_clk),
    .D(net393),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1304_ (.CLK(clknet_leaf_19_clk),
    .D(net389),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1305_ (.CLK(clknet_leaf_19_clk),
    .D(net399),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1306_ (.CLK(clknet_leaf_19_clk),
    .D(net401),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1307_ (.CLK(clknet_leaf_19_clk),
    .D(\p8div.sa.div.genblk1[8].div_n.a_ge_b ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1308_ (.CLK(clknet_leaf_19_clk),
    .D(net227),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1309_ (.CLK(clknet_leaf_20_clk),
    .D(net320),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1310_ (.CLK(clknet_leaf_20_clk),
    .D(net237),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1311_ (.CLK(clknet_leaf_20_clk),
    .D(net301),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1312_ (.CLK(clknet_leaf_20_clk),
    .D(net274),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1313_ (.CLK(clknet_leaf_20_clk),
    .D(net350),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1314_ (.CLK(clknet_leaf_20_clk),
    .D(net233),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1315_ (.CLK(clknet_leaf_15_clk),
    .D(net125),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.Q_O[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1316_ (.CLK(clknet_leaf_18_clk),
    .D(_0048_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1317_ (.CLK(clknet_leaf_18_clk),
    .D(_0049_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1318_ (.CLK(clknet_leaf_18_clk),
    .D(_0050_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1319_ (.CLK(clknet_leaf_18_clk),
    .D(_0051_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1320_ (.CLK(clknet_leaf_19_clk),
    .D(_0052_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1321_ (.CLK(clknet_leaf_19_clk),
    .D(_0053_),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1322_ (.CLK(clknet_leaf_18_clk),
    .D(net437),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1323_ (.CLK(clknet_leaf_18_clk),
    .D(net434),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1324_ (.CLK(clknet_leaf_18_clk),
    .D(net400),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1325_ (.CLK(clknet_leaf_18_clk),
    .D(net380),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1326_ (.CLK(clknet_leaf_19_clk),
    .D(net414),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1327_ (.CLK(clknet_leaf_19_clk),
    .D(net394),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1328_ (.CLK(clknet_leaf_19_clk),
    .D(\p8div.sa.div.genblk1[7].div_n.a_ge_b ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1329_ (.CLK(clknet_leaf_20_clk),
    .D(net307),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1330_ (.CLK(clknet_leaf_20_clk),
    .D(net329),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1331_ (.CLK(clknet_leaf_20_clk),
    .D(net313),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1332_ (.CLK(clknet_leaf_20_clk),
    .D(net318),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1333_ (.CLK(clknet_leaf_20_clk),
    .D(net139),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1334_ (.CLK(clknet_leaf_20_clk),
    .D(net330),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1335_ (.CLK(clknet_leaf_9_clk),
    .D(net317),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.Q_O[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1336_ (.CLK(clknet_leaf_22_clk),
    .D(_0042_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1337_ (.CLK(clknet_leaf_22_clk),
    .D(_0043_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1338_ (.CLK(clknet_leaf_21_clk),
    .D(_0044_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1339_ (.CLK(clknet_leaf_21_clk),
    .D(_0045_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1340_ (.CLK(clknet_leaf_21_clk),
    .D(_0046_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1341_ (.CLK(clknet_leaf_20_clk),
    .D(_0047_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1342_ (.CLK(clknet_leaf_22_clk),
    .D(net403),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1343_ (.CLK(clknet_leaf_22_clk),
    .D(net402),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1344_ (.CLK(clknet_leaf_22_clk),
    .D(net396),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1345_ (.CLK(clknet_leaf_21_clk),
    .D(net386),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1346_ (.CLK(clknet_leaf_20_clk),
    .D(net388),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1347_ (.CLK(clknet_leaf_20_clk),
    .D(net408),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1348_ (.CLK(clknet_leaf_20_clk),
    .D(\p8div.sa.div.genblk1[6].div_n.a_ge_b ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1349_ (.CLK(clknet_leaf_20_clk),
    .D(net355),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1350_ (.CLK(clknet_leaf_20_clk),
    .D(net321),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1351_ (.CLK(clknet_leaf_1_clk),
    .D(net273),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1352_ (.CLK(clknet_leaf_2_clk),
    .D(net373),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1353_ (.CLK(clknet_leaf_1_clk),
    .D(net328),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1354_ (.CLK(clknet_leaf_2_clk),
    .D(net370),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.Q_O[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1355_ (.CLK(clknet_leaf_22_clk),
    .D(_0036_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1356_ (.CLK(clknet_leaf_22_clk),
    .D(_0037_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1357_ (.CLK(clknet_leaf_22_clk),
    .D(_0038_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1358_ (.CLK(clknet_leaf_21_clk),
    .D(_0039_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1359_ (.CLK(clknet_leaf_21_clk),
    .D(_0040_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1360_ (.CLK(clknet_leaf_21_clk),
    .D(_0041_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1361_ (.CLK(clknet_leaf_22_clk),
    .D(net404),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1362_ (.CLK(clknet_leaf_22_clk),
    .D(net415),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1363_ (.CLK(clknet_leaf_22_clk),
    .D(net391),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1364_ (.CLK(clknet_leaf_21_clk),
    .D(net420),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1365_ (.CLK(clknet_leaf_20_clk),
    .D(net379),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1366_ (.CLK(clknet_leaf_20_clk),
    .D(net398),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1367_ (.CLK(clknet_leaf_1_clk),
    .D(\p8div.sa.div.genblk1[5].div_n.a_ge_b ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1368_ (.CLK(clknet_leaf_1_clk),
    .D(net323),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1369_ (.CLK(clknet_leaf_1_clk),
    .D(net346),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1370_ (.CLK(clknet_leaf_1_clk),
    .D(net316),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.Q_O[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1371_ (.CLK(clknet_leaf_1_clk),
    .D(net341),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.Q_O[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1372_ (.CLK(clknet_leaf_1_clk),
    .D(net340),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.Q_O[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1373_ (.CLK(clknet_leaf_22_clk),
    .D(_0030_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1374_ (.CLK(clknet_leaf_22_clk),
    .D(_0031_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1375_ (.CLK(clknet_leaf_22_clk),
    .D(_0032_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1376_ (.CLK(clknet_leaf_22_clk),
    .D(_0033_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1377_ (.CLK(clknet_leaf_23_clk),
    .D(_0034_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1378_ (.CLK(clknet_leaf_23_clk),
    .D(_0035_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1379_ (.CLK(clknet_leaf_22_clk),
    .D(net439),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1380_ (.CLK(clknet_leaf_22_clk),
    .D(net438),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1381_ (.CLK(clknet_leaf_22_clk),
    .D(net436),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1382_ (.CLK(clknet_leaf_22_clk),
    .D(net407),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1383_ (.CLK(clknet_leaf_21_clk),
    .D(net425),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1384_ (.CLK(clknet_leaf_1_clk),
    .D(net424),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1385_ (.CLK(clknet_leaf_1_clk),
    .D(\p8div.sa.div.genblk1[4].div_n.a_ge_b ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1386_ (.CLK(clknet_leaf_1_clk),
    .D(net345),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1387_ (.CLK(clknet_leaf_1_clk),
    .D(net248),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1388_ (.CLK(clknet_leaf_1_clk),
    .D(net277),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.Q_O[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1389_ (.CLK(clknet_leaf_1_clk),
    .D(net138),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.Q_O[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1390_ (.CLK(clknet_leaf_23_clk),
    .D(_0024_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1391_ (.CLK(clknet_leaf_23_clk),
    .D(_0025_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1392_ (.CLK(clknet_leaf_23_clk),
    .D(_0026_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1393_ (.CLK(clknet_leaf_23_clk),
    .D(_0027_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1394_ (.CLK(clknet_leaf_23_clk),
    .D(_0028_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1395_ (.CLK(clknet_leaf_23_clk),
    .D(_0029_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1396_ (.CLK(clknet_leaf_1_clk),
    .D(net430),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1397_ (.CLK(clknet_leaf_1_clk),
    .D(net421),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1398_ (.CLK(clknet_leaf_1_clk),
    .D(net417),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1399_ (.CLK(clknet_leaf_23_clk),
    .D(net428),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1400_ (.CLK(clknet_leaf_1_clk),
    .D(net423),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1401_ (.CLK(clknet_leaf_23_clk),
    .D(net387),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1402_ (.CLK(clknet_leaf_1_clk),
    .D(\p8div.sa.div.genblk1[3].div_n.a_ge_b ),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1403_ (.CLK(clknet_leaf_1_clk),
    .D(net343),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1404_ (.CLK(clknet_leaf_1_clk),
    .D(net292),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1405_ (.CLK(clknet_leaf_2_clk),
    .D(net129),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.Q_O[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1406_ (.CLK(clknet_leaf_0_clk),
    .D(_0018_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1407_ (.CLK(clknet_leaf_0_clk),
    .D(_0019_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1408_ (.CLK(clknet_leaf_0_clk),
    .D(_0020_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1409_ (.CLK(clknet_leaf_0_clk),
    .D(_0021_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1410_ (.CLK(clknet_leaf_0_clk),
    .D(_0022_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1411_ (.CLK(clknet_leaf_0_clk),
    .D(_0023_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1412_ (.CLK(clknet_leaf_0_clk),
    .D(net411),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1413_ (.CLK(clknet_leaf_0_clk),
    .D(net382),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1414_ (.CLK(clknet_leaf_0_clk),
    .D(net422),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1415_ (.CLK(clknet_leaf_0_clk),
    .D(net416),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1416_ (.CLK(clknet_leaf_0_clk),
    .D(net392),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1417_ (.CLK(clknet_leaf_23_clk),
    .D(net429),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1418_ (.CLK(clknet_leaf_1_clk),
    .D(\p8div.sa.div.genblk1[2].div_n.a_ge_b ),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1419_ (.CLK(clknet_leaf_1_clk),
    .D(net331),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1420_ (.CLK(clknet_leaf_3_clk),
    .D(net351),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.Q_O[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1421_ (.CLK(clknet_leaf_0_clk),
    .D(_0012_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1422_ (.CLK(clknet_leaf_0_clk),
    .D(_0013_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1423_ (.CLK(clknet_leaf_0_clk),
    .D(_0014_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1424_ (.CLK(clknet_leaf_0_clk),
    .D(_0015_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1425_ (.CLK(clknet_leaf_0_clk),
    .D(_0016_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1426_ (.CLK(clknet_leaf_0_clk),
    .D(_0017_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1427_ (.CLK(clknet_leaf_0_clk),
    .D(net419),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1428_ (.CLK(clknet_leaf_3_clk),
    .D(net390),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1429_ (.CLK(clknet_leaf_0_clk),
    .D(net383),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1430_ (.CLK(clknet_leaf_3_clk),
    .D(net381),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1431_ (.CLK(clknet_leaf_4_clk),
    .D(net385),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1432_ (.CLK(clknet_leaf_0_clk),
    .D(net418),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1433_ (.CLK(clknet_leaf_0_clk),
    .D(\p8div.sa.div.genblk1[1].div_n.a_ge_b ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.Q_O[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1434_ (.CLK(clknet_leaf_3_clk),
    .D(net298),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.Q_O[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1435_ (.CLK(clknet_leaf_3_clk),
    .D(_0000_),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1436_ (.CLK(clknet_leaf_4_clk),
    .D(_0001_),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1437_ (.CLK(clknet_leaf_4_clk),
    .D(_0002_),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1438_ (.CLK(clknet_leaf_4_clk),
    .D(_0003_),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1439_ (.CLK(clknet_leaf_4_clk),
    .D(_0004_),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1440_ (.CLK(clknet_leaf_4_clk),
    .D(_0005_),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ));
 sky130_fd_sc_hd__dfrtp_1 _1441_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.B_decode.F[0] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1442_ (.CLK(clknet_leaf_4_clk),
    .D(\p8div.B_decode.F[1] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1443_ (.CLK(clknet_leaf_4_clk),
    .D(\p8div.B_decode.F[2] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1444_ (.CLK(clknet_leaf_4_clk),
    .D(\p8div.B_decode.F[3] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1445_ (.CLK(clknet_leaf_4_clk),
    .D(\p8div.B_decode.F[4] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1446_ (.CLK(clknet_leaf_0_clk),
    .D(net113),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.div.b[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1447_ (.CLK(clknet_leaf_8_clk),
    .D(net315),
    .RESET_B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1448_ (.CLK(clknet_leaf_2_clk),
    .D(net325),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1449_ (.CLK(clknet_leaf_2_clk),
    .D(net270),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1450_ (.CLK(clknet_leaf_2_clk),
    .D(net377),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1451_ (.CLK(clknet_leaf_2_clk),
    .D(net190),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1452_ (.CLK(clknet_leaf_2_clk),
    .D(net130),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1453_ (.CLK(clknet_leaf_2_clk),
    .D(net337),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1454_ (.CLK(clknet_leaf_2_clk),
    .D(net282),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1455_ (.CLK(clknet_leaf_2_clk),
    .D(net135),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1456_ (.CLK(clknet_leaf_2_clk),
    .D(net128),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1457_ (.CLK(clknet_leaf_8_clk),
    .D(net245),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1458_ (.CLK(clknet_leaf_8_clk),
    .D(net357),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1459_ (.CLK(clknet_leaf_2_clk),
    .D(net181),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1460_ (.CLK(clknet_leaf_1_clk),
    .D(net140),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1461_ (.CLK(clknet_leaf_2_clk),
    .D(net284),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1462_ (.CLK(clknet_leaf_8_clk),
    .D(net199),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1463_ (.CLK(clknet_leaf_8_clk),
    .D(net236),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1464_ (.CLK(clknet_leaf_8_clk),
    .D(net293),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1465_ (.CLK(clknet_leaf_2_clk),
    .D(net371),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1466_ (.CLK(clknet_leaf_2_clk),
    .D(net179),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1467_ (.CLK(clknet_leaf_2_clk),
    .D(net268),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1468_ (.CLK(clknet_leaf_2_clk),
    .D(net194),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1469_ (.CLK(clknet_leaf_2_clk),
    .D(net192),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1470_ (.CLK(clknet_leaf_1_clk),
    .D(net157),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1471_ (.CLK(clknet_leaf_2_clk),
    .D(net255),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1472_ (.CLK(clknet_leaf_9_clk),
    .D(net290),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1473_ (.CLK(clknet_leaf_9_clk),
    .D(net163),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1474_ (.CLK(clknet_leaf_9_clk),
    .D(net183),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1475_ (.CLK(clknet_leaf_2_clk),
    .D(net244),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1476_ (.CLK(clknet_leaf_8_clk),
    .D(net286),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1477_ (.CLK(clknet_leaf_3_clk),
    .D(net147),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1478_ (.CLK(clknet_leaf_2_clk),
    .D(net132),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1479_ (.CLK(clknet_leaf_2_clk),
    .D(net127),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1480_ (.CLK(clknet_leaf_3_clk),
    .D(net149),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1481_ (.CLK(clknet_leaf_3_clk),
    .D(net342),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1482_ (.CLK(clknet_leaf_9_clk),
    .D(net221),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1483_ (.CLK(clknet_leaf_9_clk),
    .D(net185),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1484_ (.CLK(clknet_leaf_15_clk),
    .D(net122),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1485_ (.CLK(clknet_leaf_15_clk),
    .D(net124),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1486_ (.CLK(clknet_leaf_15_clk),
    .D(net118),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1487_ (.CLK(clknet_leaf_15_clk),
    .D(net121),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1488_ (.CLK(clknet_leaf_15_clk),
    .D(net117),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1489_ (.CLK(clknet_leaf_15_clk),
    .D(net362),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1490_ (.CLK(clknet_leaf_15_clk),
    .D(net294),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1491_ (.CLK(clknet_leaf_15_clk),
    .D(net338),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[9][4] ));
 sky130_fd_sc_hd__dfrtp_4 _1492_ (.CLK(clknet_leaf_15_clk),
    .D(net304),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_scale[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1493_ (.CLK(clknet_leaf_15_clk),
    .D(net361),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_scale[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1494_ (.CLK(clknet_leaf_15_clk),
    .D(net354),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_scale[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1495_ (.CLK(clknet_leaf_15_clk),
    .D(net291),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_scale[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1496_ (.CLK(clknet_leaf_15_clk),
    .D(net288),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.c_scale[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1497_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_0_HCA.hca_stage_0.SUM ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _1498_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _1499_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _1500_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _1501_ (.CLK(clknet_leaf_3_clk),
    .D(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p8div.sa.pipe_scale_c.a_q[0][4] ));
 sky130_fd_sc_hd__conb_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa_114  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net114));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net97));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net98));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net99));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net100));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net101));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net102));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net103));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net104));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net105));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net106));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net107));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net108));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net109));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net110));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net111));
 sky130_fd_sc_hd__conb_1 tt_um_swangust3_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net112));
 sky130_fd_sc_hd__conb_1 _1446__113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net113));
 sky130_fd_sc_hd__fa_1 \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.add_frac_sum_a.C ),
    .SUM(\p8div.sa.add_frac_sum_a.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(net114),
    .B(net96),
    .CIN(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.div_0.sub_acc.C ),
    .SUM(\p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[10].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[2].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[3].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[4].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[5].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[6].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[7].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[8].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_0_HCA.hca_stage_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[1].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[2].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[3].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.SUM ));
 sky130_fd_sc_hd__fa_1 \p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa  (.A(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.A ),
    .B(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.B ),
    .CIN(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[4].fca_stage_n.C_OUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.C_OUT ),
    .SUM(\p8div.sa.div.genblk1[9].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.SUM ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(uio_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(uio_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(uio_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(uio_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(uio_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(uio_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(uio_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_1 max_cap18 (.A(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_1 max_cap19 (.A(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 wire20 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 wire21 (.A(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 wire22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 wire23 (.A(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(\p8div.c_decoded[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 fanout31 (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 fanout33 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout35 (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 fanout62 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 fanout68 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 fanout70 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__conb_1 \p8div.sa.div.div_0.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[5].fca_stage_n.G_SKY.fa_96  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net96));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_leaf_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_leaf_15_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_12 clkload3 (.A(clknet_leaf_16_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_leaf_17_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload5 (.A(clknet_leaf_18_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_leaf_19_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_20_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_12 clkload8 (.A(clknet_leaf_21_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_leaf_22_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_12 clkload10 (.A(clknet_leaf_23_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_leaf_3_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload12 (.A(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload13 (.A(clknet_leaf_5_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload14 (.A(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload15 (.A(clknet_leaf_7_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload16 (.A(clknet_leaf_8_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload17 (.A(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload18 (.A(clknet_leaf_10_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload19 (.A(clknet_leaf_11_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload21 (.A(clknet_leaf_14_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\p8div.pipe_A.a_q[4][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\p8div.pipe_sign.a_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\p8div.sa.pipe_scale_c.a_q[8][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\p8div.sa.pipe_scale_c.a_q[7][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\p8div.pipe_B.a_q[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\p8div.pipe_A.a_q[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\p8div.sa.pipe_scale_c.a_q[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\p8div.sa.pipe_scale_c.a_q[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\p8div.pipe_A.a_q[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\p8div.sa.pipe_scale_c.a_q[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\p8div.pipe_A.a_q[3][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\p8div.sa.pipe_scale_c.a_q[0][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\p8div.sa.pipe_scale_c.a_q[1][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\p8div.sa.div.genblk1[2].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\p8div.sa.pipe_scale_c.a_q[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\p8div.pipe_B.a_q[2][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\p8div.sa.pipe_scale_c.a_q[0][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\p8div.pipe_A.a_q[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\p8div.pipe_A.a_q[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\p8div.sa.pipe_scale_c.a_q[1][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\p8div.pipe_B.a_q[2][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\p8div.pipe_B.a_q[0][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\p8div.sa.div.genblk1[3].div_n.Q_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\p8div.sa.pipe_scale_c.a_q[4][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\p8div.pipe_sign.a_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\p8div.pipe_sign.a_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\p8div.pipe_A.a_q[3][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\p8div.pipe_B.a_q[1][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\p8div.sa.pipe_scale_c.a_q[0][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\p8div.pipe_B.a_q[0][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\p8div.sa.pipe_scale_c.a_q[0][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\p8div.pipe_A.a_q[3][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\p8div.pipe_A.a_q[7][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\p8div.pipe_B.a_q[8][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\p8div.pipe_B.a_q[4][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\p8div.pipe_B.a_q[3][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\p8div.pipe_B.a_q[0][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\p8div.sa.pipe_scale_c.a_q[2][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\p8div.pipe_B.a_q[4][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\p8div.pipe_B.a_q[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\p8div.pipe_A.a_q[6][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\p8div.pipe_B.a_q[1][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\p8div.pipe_A.a_q[0][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\p8div.sa.pipe_scale_c.a_q[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\p8div.pipe_A.a_q[2][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\p8div.pipe_B.a_q[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\p8div.pipe_B.a_q[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\p8div.pipe_A.a_q[0][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\p8div.pipe_sign.a_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\p8div.pipe_B.a_q[0][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\p8div.pipe_A.a_q[4][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\p8div.pipe_B.a_q[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\p8div.pipe_A.a_q[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\p8div.pipe_B.a_q[2][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\p8div.pipe_B.a_q[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\p8div.pipe_B.a_q[3][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\p8div.pipe_B.a_q[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\p8div.pipe_B.a_q[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\p8div.sa.pipe_scale_c.a_q[5][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\p8div.pipe_A.a_q[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\p8div.sa.pipe_scale_c.a_q[4][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\p8div.pipe_B.a_q[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\p8div.sa.pipe_scale_c.a_q[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\p8div.pipe_A.a_q[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\p8div.sa.pipe_scale_c.a_q[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\p8div.pipe_A.a_q[4][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\p8div.pipe_B.a_q[3][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\p8div.pipe_A.a_q[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\p8div.pipe_A.a_q[4][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\p8div.sa.pipe_scale_c.a_q[3][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\p8div.pipe_A.a_q[8][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\p8div.sa.pipe_scale_c.a_q[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\p8div.pipe_A.a_q[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\p8div.sa.pipe_scale_c.a_q[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\p8div.pipe_B.a_q[8][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\p8div.pipe_B.a_q[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\p8div.pipe_B.a_q[9][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\p8div.sa.pipe_scale_c.a_q[5][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\p8div.pipe_sign.a_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\p8div.pipe_A.a_q[0][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\p8div.pipe_A.a_q[4][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\p8div.pipe_B.a_q[5][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\p8div.pipe_B.a_q[2][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\p8div.pipe_A.a_q[7][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\p8div.pipe_A.a_q[5][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\p8div.pipe_B.a_q[4][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\p8div.pipe_sign.a_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\p8div.pipe_B.a_q[8][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\p8div.pipe_B.a_q[9][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\p8div.pipe_A.a_q[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\p8div.pipe_A.a_q[3][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\p8div.pipe_B.a_q[3][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\p8div.pipe_B.a_q[6][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\p8div.pipe_A.a_q[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\p8div.pipe_A.a_q[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\p8div.pipe_A.a_q[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\p8div.pipe_A.a_q[1][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\p8div.pipe_A.a_q[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\p8div.pipe_A.a_q[2][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\p8div.sa.pipe_scale_c.a_q[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\p8div.pipe_sign.a_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\p8div.pipe_A.a_q[7][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\p8div.pipe_B.a_q[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\p8div.pipe_A.a_q[0][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\p8div.pipe_A.a_q[8][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\p8div.pipe_A.a_q[5][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\p8div.pipe_A.a_q[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\p8div.pipe_B.a_q[9][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\p8div.pipe_A.a_q[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\p8div.pipe_A.a_q[7][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\p8div.pipe_B.a_q[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\p8div.sa.pipe_scale_c.a_q[5][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\p8div.pipe_B.a_q[1][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\p8div.pipe_B.a_q[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\p8div.pipe_A.a_q[8][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\p8div.pipe_B.a_q[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\p8div.pipe_A.a_q[0][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\p8div.sa.pipe_scale_c.a_q[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\p8div.sa.pipe_scale_c.a_q[4][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\p8div.pipe_sign.a_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\p8div.pipe_B.a_q[8][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\p8div.sa.div.genblk1[3].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\p8div.pipe_A.a_q[0][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\p8div.pipe_B.a_q[4][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\p8div.pipe_B.a_q[0][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\p8div.sa.pipe_scale_c.a_q[2][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\p8div.pipe_A.a_q[6][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\p8div.pipe_sign.a_q[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\p8div.pipe_B.a_q[1][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\p8div.pipe_B.a_q[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\p8div.pipe_B.a_q[6][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\p8div.pipe_B.a_q[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\p8div.pipe_A.a_q[5][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\p8div.pipe_A.a_q[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\p8div.pipe_A.a_q[2][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\p8div.pipe_A.a_q[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\p8div.pipe_B.a_q[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\p8div.sa.pipe_scale_c.a_q[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\p8div.pipe_B.a_q[5][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\p8div.sa.pipe_scale_c.a_q[3][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\p8div.pipe_A.a_q[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\p8div.pipe_A.a_q[6][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\p8div.sa.div.genblk1[5].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\p8div.pipe_B.a_q[4][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\p8div.pipe_A.a_q[6][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\p8div.sa.div.genblk1[3].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\p8div.pipe_B.a_q[7][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\p8div.pipe_B.a_q[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\p8div.pipe_B.a_q[7][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\p8div.sa.pipe_scale_c.a_q[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\p8div.pipe_B.a_q[6][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\p8div.sa.pipe_scale_c.a_q[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\p8div.pipe_A.a_q[4][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\p8div.sa.pipe_scale_c.a_q[6][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\p8div.pipe_A.a_q[9][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\p8div.sa.pipe_scale_c.a_q[9][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\p8div.sa.pipe_scale_c.a_q[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\p8div.sa.pipe_scale_c.a_q[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\p8div.sa.div.genblk1[2].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\p8div.sa.pipe_scale_c.a_q[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\p8div.sa.pipe_scale_c.a_q[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\p8div.pipe_A.a_q[8][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\p8div.pipe_B.a_q[5][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\p8div.sa.div.genblk1[1].div_n.Q_I ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\p8div.pipe_B.a_q[0][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\p8div.pipe_B.a_q[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\p8div.pipe_A.a_q[1][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\p8div.pipe_A.a_q[1][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\p8div.sa.pipe_scale_c.a_q[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\p8div.pipe_A.a_q[5][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\p8div.pipe_A.a_q[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\p8div.pipe_A.a_q[9][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\p8div.pipe_A.a_q[1][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\p8div.pipe_A.a_q[5][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\p8div.pipe_sign.a_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\p8div.pipe_A.a_q[4][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\p8div.pipe_A.a_q[9][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\p8div.sa.pipe_scale_c.a_q[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\p8div.sa.div.genblk1[4].div_n.Q_O[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\p8div.pipe_B.a_q[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\p8div.sa.div.genblk1[5].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\p8div.pipe_A.a_q[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\p8div.sa.div.genblk1[4].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\p8div.pipe_B.a_q[5][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\p8div.sa.pipe_scale_c.a_q[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\p8div.pipe_A.a_q[0][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\p8div.pipe_A.a_q[1][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\p8div.sa.div.genblk1[5].div_n.Q_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\p8div.sa.div.genblk1[6].div_n.Q_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\p8div.sa.div.genblk1[1].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\p8div.pipe_B.a_q[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\p8div.pipe_B.a_q[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\p8div.pipe_A.a_q[8][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\p8div.pipe_B.a_q[0][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\p8div.pipe_B.a_q[7][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\p8div.sa.pipe_scale_c.a_q[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\p8div.sa.pipe_scale_c.a_q[8][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\p8div.pipe_A.a_q[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\p8div.sa.div.genblk1[4].div_n.Q_O[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\p8div.sa.div.genblk1[4].div_n.Q_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\p8div.sa.pipe_scale_c.a_q[0][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\p8div.sa.div.genblk1[2].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\p8div.pipe_B.a_q[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\p8div.sa.div.genblk1[3].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\p8div.sa.div.genblk1[4].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\p8div.pipe_A.a_q[5][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\p8div.pipe_B.a_q[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\p8div.pipe_A.a_q[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\p8div.sa.div.genblk1[7].div_n.Q_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\p8div.sa.div.genblk1[1].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\p8div.pipe_B.a_q[4][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\p8div.pipe_B.a_q[5][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\p8div.sa.pipe_scale_c.a_q[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\p8div.sa.div.genblk1[5].div_n.Q_O[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\p8div.pipe_A.a_q[9][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\p8div.sa.pipe_scale_c.a_q[4][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\p8div.pipe_A.a_q[2][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\p8div.pipe_A.a_q[3][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\p8div.sa.pipe_scale_c.a_q[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\p8div.sa.pipe_scale_c.a_q[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\p8div.pipe_A.a_q[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\p8div.pipe_B.a_q[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\p8div.pipe_A.a_q[2][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\p8div.pipe_B.a_q[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\p8div.pipe_A.a_q[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\p8div.pipe_A.a_q[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\p8div.pipe_A.a_q[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\p8div.sa.div.genblk1[5].div_n.Q_O[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\p8div.sa.pipe_scale_c.a_q[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\p8div.sa.div.genblk1[8].div_n.Q_O[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\p8div.sa.div.genblk1[5].div_n.Q_O[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\p8div.sa.div.genblk1[10].div_n.Q_I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\p8div.sa.pipe_scale_c.a_q[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\p8div.pipe_A.a_q[0][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\p8div.sa.div.b[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\p8div.sa.div.b[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\p8div.sa.div.b[0][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\p8div.sa.div.b[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\p8div.sa.div.b[0][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\p8div.pipe_B.a_q[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\p8div.sa.div.b[0][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\p8div.sa.div.b[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\p8div.sa.div.b[2][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\p8div.sa.div.b[5][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\p8div.sa.div.b[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\p8div.sa.div.b[0][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\p8div.sa.div.b[4][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\p8div.sa.div.b[1][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\p8div.sa.div.b[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\p8div.sa.div.b[6][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\p8div.sa.div.b[9][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\p8div.sa.div.b[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\p8div.sa.div.b[8][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\p8div.sa.div.b[4][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\p8div.sa.div.b[7][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\p8div.sa.div.b[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\p8div.sa.div.b[7][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\p8div.sa.div.b[5][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\p8div.sa.div.b[5][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\p8div.sa.div.b[4][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\p8div.sa.div.b[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\p8div.sa.div.b[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\p8div.sa.div.b[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\p8div.sa.div.b[5][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\p8div.sa.div.b[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\p8div.sa.div.b[8][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\p8div.sa.div.b[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\p8div.sa.div.b[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\p8div.sa.div.b[8][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\p8div.sa.div.b[6][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\p8div.sa.div.b[4][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\p8div.sa.div.b[1][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\p8div.sa.div.b[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\p8div.sa.div.b[0][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\p8div.sa.div.b[0][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\p8div.sa.div.b[4][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\p8div.sa.div.b[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\p8div.sa.div.b[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\p8div.sa.div.b[2][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\p8div.sa.div.b[3][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\p8div.sa.div.b[3][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\p8div.sa.div.b[9][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\p8div.sa.div.b[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\p8div.sa.div.b[2][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\p8div.sa.div.b[1][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\p8div.sa.div.b[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\p8div.sa.div.b[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\p8div.sa.div.b[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\p8div.sa.div.b[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\p8div.sa.div.b[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\p8div.sa.div.b[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\p8div.sa.div.b[3][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\p8div.sa.div.b[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\p8div.sa.div.b[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\p8div.sa.div.b[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\p8div.sa.div.genblk1[1].div_n.sub_acc.G_RCA.RCA_0.G_N_FCA.SN[6].fca_stage_n.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\p8div.sa.div.b[5][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\p8div.pipe_A.a_q[7][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_2_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_164 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_223 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_295 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_304 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_7_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_7_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_8_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_9_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_9_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_187 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_10_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_10_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_202 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_11_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_12_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_132 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_308 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_13_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_14_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_14_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_14_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_15_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_15_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_302 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_314 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_16_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_16_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_133 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_17_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_180 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_192 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_17_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_18_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_282 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_18_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_18_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_19_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_258 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_20_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_296 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_21_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_78 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_300 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_312 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_102 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_266 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_278 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_22_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_23_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_24_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_191 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_58 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_26_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_163 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_211 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_26_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_26_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_284 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_296 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_26_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_27_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_66 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_28_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_120 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_28_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_29_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_47 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_63 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_31_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_31_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_31_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_31_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_32_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_235 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_32_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_32_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_32_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_260 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_34_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_180 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_34_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_34_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_34_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_35_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_36_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_36_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_36_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_245 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_37_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_303 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_37_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_38_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_38_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_38_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_38_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_39_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_39_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_86 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_39_98 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_39_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_304 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_39_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_39_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_40_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_41_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_41_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_41_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_41_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_42_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_283 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_42_295 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_42_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_42_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_42_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_28 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_43_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_43_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_43_297 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_43_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_43_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_43_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_44_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_274 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_44_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_45_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_45_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_45_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_40 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_46_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_46_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_46_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_47_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_47_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_47_300 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_47_312 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_47_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_269 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_48_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_48_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_48_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_49_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_49_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_50_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_213 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_50_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_50_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_23 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_51_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_307 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_51_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_51_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_52_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_296 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_52_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_52_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_52_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_53_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_78 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_53_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_53_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_53_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_210 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_53_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_53_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_303 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_54_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_296 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_55_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_55_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_55_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_178 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_55_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_55_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_56_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_47 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_56_59 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_56_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_56_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_56_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_266 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_56_286 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_56_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_57_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_57_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_57_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_57_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_57_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_58_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_89 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_58_101 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_58_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_58_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_59_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_59_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_59_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_59_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_59_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_60_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_60_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_60_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_60_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_60_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_60_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_60_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_60_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_61_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_61_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_61_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_260 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_61_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_62_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_62_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_49 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_72 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_128 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_62_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_62_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_62_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_63_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_87 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_63_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_64_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_105 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_117 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_64_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_65_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_65_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_65_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_70 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_66_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_67_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_67_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_68_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_69_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_70_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_96 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_71_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_71_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_71_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_72_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_73_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_73_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_74_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_70 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_74_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_74_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_75_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_75_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_83 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_75_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_75_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_76_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_77_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_77_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_78_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_78_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_78_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_78_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_79_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_79_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_79_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_79_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_80_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_80_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_80_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_80_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net97;
 assign uio_oe[1] = net98;
 assign uio_oe[2] = net99;
 assign uio_oe[3] = net100;
 assign uio_oe[4] = net101;
 assign uio_oe[5] = net102;
 assign uio_oe[6] = net103;
 assign uio_oe[7] = net104;
 assign uio_out[0] = net105;
 assign uio_out[1] = net106;
 assign uio_out[2] = net107;
 assign uio_out[3] = net108;
 assign uio_out[4] = net109;
 assign uio_out[5] = net110;
 assign uio_out[6] = net111;
 assign uio_out[7] = net112;
endmodule
