VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_jyblue1001_pll
  CLASS BLOCK ;
  FOREIGN tt_um_jyblue1001_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.705000 ;
    ANTENNADIFFAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 74.085 98.045 87.515 100.665 ;
      LAYER pwell ;
        RECT 66.200 96.050 66.600 97.450 ;
        RECT 56.250 95.285 62.950 96.050 ;
      LAYER nwell ;
        RECT 42.835 84.285 45.455 95.125 ;
        RECT 46.735 76.435 49.355 95.155 ;
        RECT 50.635 82.555 54.915 95.165 ;
      LAYER pwell ;
        RECT 56.250 90.115 57.015 95.285 ;
        RECT 62.185 90.115 62.950 95.285 ;
        RECT 56.250 89.350 62.950 90.115 ;
        RECT 63.050 95.285 69.750 96.050 ;
        RECT 63.050 90.115 63.815 95.285 ;
        RECT 68.985 90.115 69.750 95.285 ;
        RECT 63.050 89.350 69.750 90.115 ;
        RECT 69.850 95.285 76.550 96.050 ;
        RECT 69.850 90.115 70.615 95.285 ;
        RECT 75.785 90.115 76.550 95.285 ;
        RECT 69.850 89.350 76.550 90.115 ;
        RECT 56.250 88.485 62.950 89.250 ;
        RECT 56.250 83.315 57.015 88.485 ;
        RECT 62.185 83.315 62.950 88.485 ;
        RECT 56.250 82.550 62.950 83.315 ;
        RECT 63.050 88.485 69.750 89.250 ;
        RECT 63.050 83.315 63.815 88.485 ;
        RECT 68.985 83.315 69.750 88.485 ;
        RECT 63.050 82.550 69.750 83.315 ;
        RECT 69.850 88.485 76.550 89.250 ;
        RECT 69.850 83.315 70.615 88.485 ;
        RECT 75.785 83.315 76.550 88.485 ;
        RECT 69.850 82.550 76.550 83.315 ;
      LAYER nwell ;
        RECT 77.235 82.555 81.515 95.165 ;
      LAYER pwell ;
        RECT 56.250 81.685 62.950 82.450 ;
        RECT 56.250 76.515 57.015 81.685 ;
        RECT 62.185 76.515 62.950 81.685 ;
        RECT 56.250 75.750 62.950 76.515 ;
        RECT 63.050 81.685 69.750 82.450 ;
        RECT 63.050 76.515 63.815 81.685 ;
        RECT 68.985 76.515 69.750 81.685 ;
        RECT 63.050 75.750 69.750 76.515 ;
        RECT 69.850 81.685 76.550 82.450 ;
        RECT 69.850 76.515 70.615 81.685 ;
        RECT 75.785 76.515 76.550 81.685 ;
      LAYER nwell ;
        RECT 82.785 80.885 85.405 95.155 ;
        RECT 86.735 84.285 89.355 95.125 ;
      LAYER pwell ;
        RECT 69.850 75.750 76.550 76.515 ;
      LAYER nwell ;
        RECT 56.835 72.585 75.945 75.205 ;
        RECT 96.500 59.450 113.700 66.000 ;
        RECT 52.000 57.900 65.650 59.300 ;
        RECT 67.150 57.900 80.800 59.300 ;
        RECT 114.985 59.135 117.605 70.955 ;
        RECT 57.500 50.100 75.300 53.500 ;
        RECT 76.800 51.100 80.650 52.500 ;
        RECT 57.550 47.100 65.750 48.500 ;
        RECT 67.050 47.100 75.250 48.500 ;
        RECT 114.985 47.785 117.605 57.855 ;
        RECT 65.650 32.350 90.550 38.550 ;
        RECT 96.950 32.500 113.050 35.400 ;
        RECT 61.300 16.950 113.850 18.000 ;
        RECT 115.250 16.700 126.800 27.850 ;
      LAYER pwell ;
        RECT 115.250 9.200 125.850 16.300 ;
      LAYER li1 ;
        RECT 80.600 100.485 81.000 100.500 ;
        RECT 74.265 100.315 87.335 100.485 ;
        RECT 74.265 98.395 74.435 100.315 ;
        RECT 80.600 100.100 81.000 100.315 ;
        RECT 74.960 99.180 77.120 99.530 ;
        RECT 84.480 99.180 86.640 99.530 ;
        RECT 87.165 98.395 87.335 100.315 ;
        RECT 74.265 98.225 87.335 98.395 ;
        RECT 62.800 95.920 63.200 95.950 ;
        RECT 66.200 95.920 66.600 97.450 ;
        RECT 69.600 95.920 70.000 95.950 ;
        RECT 56.380 95.425 76.420 95.920 ;
        RECT 43.950 94.945 44.350 95.050 ;
        RECT 47.850 94.975 48.250 95.100 ;
        RECT 53.400 94.985 53.800 95.150 ;
        RECT 43.015 94.775 45.275 94.945 ;
        RECT 43.015 84.635 43.185 94.775 ;
        RECT 43.950 94.650 44.350 94.775 ;
        RECT 43.800 92.090 44.490 94.250 ;
        RECT 43.800 85.160 44.490 87.320 ;
        RECT 45.105 84.635 45.275 94.775 ;
        RECT 43.015 84.465 45.275 84.635 ;
        RECT 46.915 94.805 49.175 94.975 ;
        RECT 46.915 76.785 47.085 94.805 ;
        RECT 47.850 94.700 48.250 94.805 ;
        RECT 47.870 92.120 48.220 94.280 ;
        RECT 47.870 77.310 48.220 79.470 ;
        RECT 49.005 76.785 49.175 94.805 ;
        RECT 50.815 94.815 54.735 94.985 ;
        RECT 50.815 82.905 50.985 94.815 ;
        RECT 53.400 94.750 53.800 94.815 ;
        RECT 53.430 92.130 53.780 94.290 ;
        RECT 51.770 83.430 52.120 85.590 ;
        RECT 54.565 82.905 54.735 94.815 ;
        RECT 56.380 90.700 56.875 95.425 ;
        RECT 57.195 94.745 62.005 95.105 ;
        RECT 57.195 90.700 57.555 94.745 ;
        RECT 57.865 90.965 61.335 94.435 ;
        RECT 61.645 90.700 62.005 94.745 ;
        RECT 62.325 90.700 63.675 95.425 ;
        RECT 63.995 94.745 68.805 95.105 ;
        RECT 63.995 90.700 64.355 94.745 ;
        RECT 64.665 90.965 68.135 94.435 ;
        RECT 68.445 90.700 68.805 94.745 ;
        RECT 69.125 90.700 70.475 95.425 ;
        RECT 70.795 94.745 75.605 95.105 ;
        RECT 70.795 90.700 71.155 94.745 ;
        RECT 71.465 90.965 74.935 94.435 ;
        RECT 75.245 90.700 75.605 94.745 ;
        RECT 75.925 90.700 76.420 95.425 ;
        RECT 78.350 94.985 78.750 95.150 ;
        RECT 77.415 94.815 81.335 94.985 ;
        RECT 83.900 94.975 84.300 95.150 ;
        RECT 56.350 89.450 76.450 90.700 ;
        RECT 62.800 89.120 63.200 89.450 ;
        RECT 69.600 89.120 70.000 89.450 ;
        RECT 56.380 88.625 76.420 89.120 ;
        RECT 56.380 83.900 56.875 88.625 ;
        RECT 57.195 87.945 62.005 88.305 ;
        RECT 57.195 83.900 57.555 87.945 ;
        RECT 57.865 84.165 61.335 87.635 ;
        RECT 61.645 83.900 62.005 87.945 ;
        RECT 62.325 83.900 63.675 88.625 ;
        RECT 63.995 87.945 68.805 88.305 ;
        RECT 63.995 83.900 64.355 87.945 ;
        RECT 64.665 84.165 68.135 87.635 ;
        RECT 68.445 83.900 68.805 87.945 ;
        RECT 69.125 83.900 70.475 88.625 ;
        RECT 70.795 87.945 75.605 88.305 ;
        RECT 70.795 83.900 71.155 87.945 ;
        RECT 71.465 84.165 74.935 87.635 ;
        RECT 75.245 83.900 75.605 87.945 ;
        RECT 75.925 83.900 76.420 88.625 ;
        RECT 50.815 82.735 54.735 82.905 ;
        RECT 56.350 82.650 76.450 83.900 ;
        RECT 77.415 82.905 77.585 94.815 ;
        RECT 78.350 94.750 78.750 94.815 ;
        RECT 78.370 92.130 78.720 94.290 ;
        RECT 80.030 83.430 80.380 85.590 ;
        RECT 81.165 82.905 81.335 94.815 ;
        RECT 77.415 82.735 81.335 82.905 ;
        RECT 82.965 94.805 85.225 94.975 ;
        RECT 87.850 94.945 88.250 95.050 ;
        RECT 62.800 82.320 63.200 82.650 ;
        RECT 69.600 82.320 70.000 82.650 ;
        RECT 56.380 81.825 76.420 82.320 ;
        RECT 56.380 77.100 56.875 81.825 ;
        RECT 57.195 81.145 62.005 81.505 ;
        RECT 57.195 77.100 57.555 81.145 ;
        RECT 57.865 77.365 61.335 80.835 ;
        RECT 61.645 77.100 62.005 81.145 ;
        RECT 62.325 77.100 63.675 81.825 ;
        RECT 63.995 81.145 68.805 81.505 ;
        RECT 63.995 77.100 64.355 81.145 ;
        RECT 64.665 77.365 68.135 80.835 ;
        RECT 68.445 77.100 68.805 81.145 ;
        RECT 69.125 77.100 70.475 81.825 ;
        RECT 70.795 81.145 75.605 81.505 ;
        RECT 70.795 77.100 71.155 81.145 ;
        RECT 71.465 77.365 74.935 80.835 ;
        RECT 75.245 77.100 75.605 81.145 ;
        RECT 75.925 77.100 76.420 81.825 ;
        RECT 82.965 81.235 83.135 94.805 ;
        RECT 83.900 94.750 84.300 94.805 ;
        RECT 83.920 92.120 84.270 94.280 ;
        RECT 83.920 81.760 84.270 83.920 ;
        RECT 85.055 81.235 85.225 94.805 ;
        RECT 86.915 94.775 89.175 94.945 ;
        RECT 86.915 84.635 87.085 94.775 ;
        RECT 87.850 94.650 88.250 94.775 ;
        RECT 87.700 92.090 88.390 94.250 ;
        RECT 87.700 85.160 88.390 87.320 ;
        RECT 89.005 84.635 89.175 94.775 ;
        RECT 86.915 84.465 89.175 84.635 ;
        RECT 82.965 81.065 85.225 81.235 ;
        RECT 46.915 76.615 49.175 76.785 ;
        RECT 56.350 75.850 76.450 77.100 ;
        RECT 57.015 74.855 75.765 75.025 ;
        RECT 57.015 72.935 57.185 74.855 ;
        RECT 57.710 73.720 59.870 74.070 ;
        RECT 72.910 73.720 75.070 74.070 ;
        RECT 75.595 73.550 75.765 74.855 ;
        RECT 75.500 73.150 75.900 73.550 ;
        RECT 75.595 72.935 75.765 73.150 ;
        RECT 57.015 72.765 75.765 72.935 ;
        RECT 55.850 71.100 56.150 71.350 ;
        RECT 55.400 70.700 56.150 71.100 ;
        RECT 55.850 70.450 56.150 70.700 ;
        RECT 66.250 70.450 66.550 71.350 ;
        RECT 76.650 71.300 77.350 71.350 ;
        RECT 76.650 70.500 77.750 71.300 ;
        RECT 115.165 70.605 117.425 70.775 ;
        RECT 76.650 70.450 77.350 70.500 ;
        RECT 55.900 70.250 56.100 70.450 ;
        RECT 66.300 70.250 66.500 70.450 ;
        RECT 55.800 69.850 56.200 70.250 ;
        RECT 56.600 69.850 57.000 70.250 ;
        RECT 57.400 69.850 57.800 70.250 ;
        RECT 58.200 69.850 58.600 70.250 ;
        RECT 59.000 69.850 59.400 70.250 ;
        RECT 59.800 69.850 60.200 70.250 ;
        RECT 60.600 69.850 61.000 70.250 ;
        RECT 61.400 69.850 61.800 70.250 ;
        RECT 62.200 69.850 62.600 70.250 ;
        RECT 63.000 69.850 63.400 70.250 ;
        RECT 63.800 69.850 64.200 70.250 ;
        RECT 64.600 69.850 65.000 70.250 ;
        RECT 65.400 69.850 65.800 70.250 ;
        RECT 66.200 69.850 66.600 70.250 ;
        RECT 67.000 69.850 67.400 70.250 ;
        RECT 67.800 69.850 68.200 70.250 ;
        RECT 68.600 69.850 69.000 70.250 ;
        RECT 69.400 69.850 69.800 70.250 ;
        RECT 70.200 69.850 70.600 70.250 ;
        RECT 71.000 69.850 71.400 70.250 ;
        RECT 71.800 69.850 72.200 70.250 ;
        RECT 72.600 69.850 73.000 70.250 ;
        RECT 73.400 69.850 73.800 70.250 ;
        RECT 74.200 69.850 74.600 70.250 ;
        RECT 75.000 69.850 75.400 70.250 ;
        RECT 75.800 69.850 76.200 70.250 ;
        RECT 59.500 68.300 59.900 68.900 ;
        RECT 72.900 68.300 73.300 68.900 ;
        RECT 53.750 65.900 54.050 68.300 ;
        RECT 59.150 65.900 60.250 68.300 ;
        RECT 53.700 65.500 54.100 65.900 ;
        RECT 54.600 65.300 55.000 65.700 ;
        RECT 55.800 65.300 56.200 65.700 ;
        RECT 57.000 65.300 57.400 65.700 ;
        RECT 58.200 65.300 58.600 65.700 ;
        RECT 61.400 65.300 61.800 65.700 ;
        RECT 62.600 65.300 63.000 65.700 ;
        RECT 63.800 65.300 64.200 65.700 ;
        RECT 65.350 65.450 65.650 68.300 ;
        RECT 67.150 65.450 67.450 68.300 ;
        RECT 72.550 65.900 73.650 68.300 ;
        RECT 78.750 65.900 79.050 68.300 ;
        RECT 115.165 67.950 115.335 70.605 ;
        RECT 115.050 67.550 115.450 67.950 ;
        RECT 116.120 67.920 116.470 70.080 ;
        RECT 68.600 65.300 69.000 65.700 ;
        RECT 69.800 65.300 70.200 65.700 ;
        RECT 71.000 65.300 71.400 65.700 ;
        RECT 74.200 65.300 74.600 65.700 ;
        RECT 75.400 65.300 75.800 65.700 ;
        RECT 76.600 65.300 77.000 65.700 ;
        RECT 77.800 65.300 78.200 65.700 ;
        RECT 101.600 65.600 102.000 66.000 ;
        RECT 103.600 65.600 104.000 66.000 ;
        RECT 57.155 63.450 57.445 63.800 ;
        RECT 58.955 63.450 59.245 63.800 ;
        RECT 59.555 63.450 59.845 63.800 ;
        RECT 61.355 63.450 61.645 63.800 ;
        RECT 61.955 63.450 62.245 63.800 ;
        RECT 56.850 62.850 57.150 63.250 ;
        RECT 57.450 62.850 57.750 63.250 ;
        RECT 58.050 62.850 58.350 63.250 ;
        RECT 58.650 62.850 58.950 63.250 ;
        RECT 59.250 62.850 59.550 63.250 ;
        RECT 59.850 62.850 60.150 63.250 ;
        RECT 60.450 62.850 60.750 63.250 ;
        RECT 61.050 62.850 61.350 63.250 ;
        RECT 61.650 62.850 61.950 63.250 ;
        RECT 62.250 62.850 62.550 63.250 ;
        RECT 62.850 62.850 63.150 63.250 ;
        RECT 57.660 62.300 57.950 62.650 ;
        RECT 58.450 62.300 58.740 62.650 ;
        RECT 60.070 62.300 60.360 62.650 ;
        RECT 60.840 62.300 61.130 62.650 ;
        RECT 62.460 62.300 62.750 62.650 ;
        RECT 64.000 62.500 64.400 63.700 ;
        RECT 68.400 62.500 68.800 63.700 ;
        RECT 70.555 63.450 70.845 63.800 ;
        RECT 71.155 63.450 71.445 63.800 ;
        RECT 72.955 63.450 73.245 63.800 ;
        RECT 73.555 63.450 73.845 63.800 ;
        RECT 75.355 63.450 75.645 63.800 ;
        RECT 69.650 62.850 69.950 63.250 ;
        RECT 70.250 62.850 70.550 63.250 ;
        RECT 70.850 62.850 71.150 63.250 ;
        RECT 71.450 62.850 71.750 63.250 ;
        RECT 72.050 62.850 72.350 63.250 ;
        RECT 72.650 62.850 72.950 63.250 ;
        RECT 73.250 62.850 73.550 63.250 ;
        RECT 73.850 62.850 74.150 63.250 ;
        RECT 74.450 62.850 74.750 63.250 ;
        RECT 75.050 62.850 75.350 63.250 ;
        RECT 75.650 62.850 75.950 63.250 ;
        RECT 97.100 63.000 98.000 65.400 ;
        RECT 98.600 63.000 99.000 65.400 ;
        RECT 99.600 63.000 100.000 65.400 ;
        RECT 100.600 63.000 101.000 65.400 ;
        RECT 101.600 63.000 102.000 65.400 ;
        RECT 102.600 63.000 103.000 65.400 ;
        RECT 103.600 63.000 104.000 65.400 ;
        RECT 104.600 63.000 105.000 65.400 ;
        RECT 105.600 63.000 106.000 65.400 ;
        RECT 106.600 63.000 107.000 65.400 ;
        RECT 107.600 63.000 108.500 65.400 ;
        RECT 70.050 62.300 70.340 62.650 ;
        RECT 71.670 62.300 71.960 62.650 ;
        RECT 72.440 62.300 72.730 62.650 ;
        RECT 74.060 62.300 74.350 62.650 ;
        RECT 74.850 62.300 75.140 62.650 ;
        RECT 97.600 62.400 98.000 63.000 ;
        RECT 107.600 62.400 108.000 62.800 ;
        RECT 105.000 61.600 105.400 62.000 ;
        RECT 110.600 61.600 111.000 62.000 ;
        RECT 97.550 61.050 97.950 61.250 ;
        RECT 99.600 61.050 100.000 61.450 ;
        RECT 100.850 61.050 101.250 61.250 ;
        RECT 103.250 61.050 103.650 61.250 ;
        RECT 105.000 61.050 105.200 61.600 ;
        RECT 106.550 61.050 106.950 61.250 ;
        RECT 108.950 61.050 109.350 61.250 ;
        RECT 110.700 61.050 110.900 61.600 ;
        RECT 112.250 61.050 112.650 61.250 ;
        RECT 97.350 60.850 101.450 61.050 ;
        RECT 97.350 60.650 97.550 60.850 ;
        RECT 98.000 60.650 98.200 60.850 ;
        RECT 99.300 60.650 99.500 60.850 ;
        RECT 100.600 60.650 100.800 60.850 ;
        RECT 101.250 60.650 101.450 60.850 ;
        RECT 103.050 60.850 107.150 61.050 ;
        RECT 103.050 60.650 103.250 60.850 ;
        RECT 103.700 60.650 103.900 60.850 ;
        RECT 105.000 60.650 105.200 60.850 ;
        RECT 106.300 60.650 106.500 60.850 ;
        RECT 106.950 60.650 107.150 60.850 ;
        RECT 108.750 60.850 112.850 61.050 ;
        RECT 108.750 60.650 108.950 60.850 ;
        RECT 109.400 60.650 109.600 60.850 ;
        RECT 110.700 60.650 110.900 60.850 ;
        RECT 112.000 60.650 112.200 60.850 ;
        RECT 112.650 60.650 112.850 60.850 ;
        RECT 97.250 59.750 97.650 60.650 ;
        RECT 97.900 59.750 98.300 60.650 ;
        RECT 98.550 59.750 98.950 60.650 ;
        RECT 99.200 59.750 99.600 60.650 ;
        RECT 99.850 59.750 100.250 60.650 ;
        RECT 100.500 59.750 100.950 60.650 ;
        RECT 101.150 59.750 101.550 60.650 ;
        RECT 102.450 59.750 103.350 60.650 ;
        RECT 103.600 59.750 104.000 60.650 ;
        RECT 104.250 59.750 104.650 60.650 ;
        RECT 104.900 59.750 105.300 60.650 ;
        RECT 105.550 59.750 105.950 60.650 ;
        RECT 106.200 59.750 106.600 60.650 ;
        RECT 106.850 59.750 107.750 60.650 ;
        RECT 108.150 59.750 109.050 60.650 ;
        RECT 109.300 59.750 109.700 60.650 ;
        RECT 109.950 59.750 110.350 60.650 ;
        RECT 110.600 59.750 111.000 60.650 ;
        RECT 111.250 59.750 111.650 60.650 ;
        RECT 111.900 59.750 112.300 60.650 ;
        RECT 112.550 59.750 113.450 60.650 ;
        RECT 53.550 59.300 53.850 59.700 ;
        RECT 54.400 59.250 54.800 59.650 ;
        RECT 56.850 59.250 57.150 59.650 ;
        RECT 58.000 59.250 58.400 59.650 ;
        RECT 60.450 59.250 60.750 59.650 ;
        RECT 61.600 59.250 62.000 59.650 ;
        RECT 63.750 59.250 64.050 59.650 ;
        RECT 68.750 59.250 69.050 59.650 ;
        RECT 70.800 59.250 71.200 59.650 ;
        RECT 72.050 59.250 72.350 59.650 ;
        RECT 74.400 59.250 74.800 59.650 ;
        RECT 75.650 59.250 75.950 59.650 ;
        RECT 78.000 59.250 78.400 59.650 ;
        RECT 78.950 59.300 79.250 59.700 ;
        RECT 98.100 59.150 98.500 59.550 ;
        RECT 100.300 59.150 100.700 59.550 ;
        RECT 104.250 59.100 104.650 59.500 ;
        RECT 109.500 59.150 109.900 59.550 ;
        RECT 52.250 58.150 52.950 59.050 ;
        RECT 53.250 58.150 53.550 59.050 ;
        RECT 53.850 58.150 54.150 59.050 ;
        RECT 54.450 58.150 54.750 59.050 ;
        RECT 55.050 58.150 55.350 59.050 ;
        RECT 55.650 58.150 55.950 59.050 ;
        RECT 56.250 58.150 56.550 59.050 ;
        RECT 56.850 58.150 57.150 59.050 ;
        RECT 57.450 58.150 57.750 59.050 ;
        RECT 58.050 58.150 58.350 59.050 ;
        RECT 58.650 58.150 58.950 59.050 ;
        RECT 59.250 58.150 59.550 59.050 ;
        RECT 59.850 58.150 60.150 59.050 ;
        RECT 60.450 58.150 60.750 59.050 ;
        RECT 61.050 58.150 61.350 59.050 ;
        RECT 61.650 58.150 61.950 59.050 ;
        RECT 62.250 58.150 62.550 59.050 ;
        RECT 62.850 58.150 63.150 59.050 ;
        RECT 63.450 58.150 63.750 59.050 ;
        RECT 64.050 58.150 64.350 59.050 ;
        RECT 64.650 58.150 65.350 59.050 ;
        RECT 67.450 58.150 68.150 59.050 ;
        RECT 68.450 58.150 68.750 59.050 ;
        RECT 69.050 58.150 69.350 59.050 ;
        RECT 69.650 58.150 69.950 59.050 ;
        RECT 70.250 58.150 70.550 59.050 ;
        RECT 70.850 58.150 71.150 59.050 ;
        RECT 71.450 58.150 71.750 59.050 ;
        RECT 72.050 58.150 72.350 59.050 ;
        RECT 72.650 58.150 72.950 59.050 ;
        RECT 73.250 58.150 73.550 59.050 ;
        RECT 73.850 58.150 74.150 59.050 ;
        RECT 74.450 58.150 74.750 59.050 ;
        RECT 75.050 58.150 75.350 59.050 ;
        RECT 75.650 58.150 75.950 59.050 ;
        RECT 76.250 58.150 76.550 59.050 ;
        RECT 76.850 58.150 77.150 59.050 ;
        RECT 77.450 58.150 77.750 59.050 ;
        RECT 78.050 58.150 78.350 59.050 ;
        RECT 78.650 58.150 78.950 59.050 ;
        RECT 79.250 58.150 79.550 59.050 ;
        RECT 79.850 58.150 80.550 59.050 ;
        RECT 110.150 58.700 110.350 59.750 ;
        RECT 111.250 58.700 111.450 59.750 ;
        RECT 113.700 59.150 114.100 59.550 ;
        RECT 115.165 59.485 115.335 67.550 ;
        RECT 116.120 60.010 116.470 62.170 ;
        RECT 117.255 59.485 117.425 70.605 ;
        RECT 115.165 59.315 117.425 59.485 ;
        RECT 109.500 58.050 109.900 58.450 ;
        RECT 110.150 58.300 110.550 58.700 ;
        RECT 111.150 58.300 111.550 58.700 ;
        RECT 117.800 58.300 118.200 58.700 ;
        RECT 52.650 57.550 52.950 57.950 ;
        RECT 64.650 57.550 64.950 57.950 ;
        RECT 67.850 57.550 68.150 57.950 ;
        RECT 79.850 57.550 80.150 57.950 ;
        RECT 98.550 57.450 98.950 57.850 ;
        RECT 103.800 57.450 104.200 57.850 ;
        RECT 106.000 57.450 106.400 57.850 ;
        RECT 110.150 57.250 110.350 58.300 ;
        RECT 111.250 57.250 111.450 58.300 ;
        RECT 113.700 57.450 114.100 57.850 ;
        RECT 115.165 57.505 117.425 57.675 ;
        RECT 96.750 56.850 97.650 57.250 ;
        RECT 97.900 56.850 98.300 57.250 ;
        RECT 98.550 56.850 98.950 57.250 ;
        RECT 99.200 56.850 99.600 57.250 ;
        RECT 99.850 56.850 100.250 57.250 ;
        RECT 100.500 56.850 100.900 57.250 ;
        RECT 101.150 56.850 102.050 57.250 ;
        RECT 102.950 56.850 103.350 57.250 ;
        RECT 103.600 56.850 104.000 57.250 ;
        RECT 104.250 56.850 104.650 57.250 ;
        RECT 104.900 56.850 105.300 57.250 ;
        RECT 105.550 56.850 105.950 57.250 ;
        RECT 106.200 56.850 106.600 57.250 ;
        RECT 106.850 56.850 107.250 57.250 ;
        RECT 108.150 56.850 109.050 57.250 ;
        RECT 109.300 56.850 109.700 57.250 ;
        RECT 109.950 56.850 110.350 57.250 ;
        RECT 110.600 56.850 111.000 57.250 ;
        RECT 111.250 56.850 111.650 57.250 ;
        RECT 111.900 56.850 112.300 57.250 ;
        RECT 112.550 56.850 113.450 57.250 ;
        RECT 97.350 56.650 97.550 56.850 ;
        RECT 98.000 56.650 98.200 56.850 ;
        RECT 99.300 56.650 99.500 56.850 ;
        RECT 100.600 56.650 100.800 56.850 ;
        RECT 101.250 56.650 101.450 56.850 ;
        RECT 97.350 56.450 101.450 56.650 ;
        RECT 103.050 56.650 103.250 56.850 ;
        RECT 103.700 56.650 103.900 56.850 ;
        RECT 105.000 56.650 105.200 56.850 ;
        RECT 106.300 56.650 106.500 56.850 ;
        RECT 106.950 56.650 107.150 56.850 ;
        RECT 103.050 56.450 107.150 56.650 ;
        RECT 108.750 56.650 108.950 56.850 ;
        RECT 109.400 56.650 109.600 56.850 ;
        RECT 110.700 56.650 110.900 56.850 ;
        RECT 112.000 56.650 112.200 56.850 ;
        RECT 112.650 56.650 112.850 56.850 ;
        RECT 97.550 56.200 98.000 56.450 ;
        RECT 99.300 55.900 99.500 56.450 ;
        RECT 100.800 56.200 101.250 56.450 ;
        RECT 103.250 56.250 103.650 56.450 ;
        RECT 104.900 56.050 105.300 56.450 ;
        RECT 106.550 56.250 106.950 56.450 ;
        RECT 108.750 56.400 112.850 56.650 ;
        RECT 108.950 56.250 109.350 56.400 ;
        RECT 110.700 55.900 110.900 56.400 ;
        RECT 112.250 56.250 112.650 56.400 ;
        RECT 99.200 55.500 99.600 55.900 ;
        RECT 110.600 55.500 111.000 55.900 ;
        RECT 97.000 54.750 97.400 55.150 ;
        RECT 104.900 54.950 105.300 55.350 ;
        RECT 99.100 54.750 105.300 54.950 ;
        RECT 107.000 54.750 107.400 55.150 ;
        RECT 97.100 54.550 97.300 54.750 ;
        RECT 99.100 54.550 99.300 54.750 ;
        RECT 105.100 54.550 105.300 54.750 ;
        RECT 107.100 54.550 107.300 54.750 ;
        RECT 59.500 53.450 59.850 53.850 ;
        RECT 60.350 53.450 60.750 53.850 ;
        RECT 61.250 53.450 61.650 53.850 ;
        RECT 62.150 53.450 62.550 53.850 ;
        RECT 63.050 53.450 63.450 53.850 ;
        RECT 63.950 53.450 64.350 53.850 ;
        RECT 64.850 53.450 65.250 53.850 ;
        RECT 65.750 53.450 66.100 53.850 ;
        RECT 66.700 53.450 67.050 53.850 ;
        RECT 67.550 53.450 67.950 53.850 ;
        RECT 68.450 53.450 68.850 53.850 ;
        RECT 69.350 53.450 69.750 53.850 ;
        RECT 70.250 53.450 70.650 53.850 ;
        RECT 71.150 53.450 71.550 53.850 ;
        RECT 72.050 53.450 72.450 53.850 ;
        RECT 72.950 53.450 73.300 53.850 ;
        RECT 96.500 53.400 97.400 54.550 ;
        RECT 98.000 53.400 98.400 54.550 ;
        RECT 99.000 53.400 99.400 54.550 ;
        RECT 100.000 53.400 100.400 54.550 ;
        RECT 101.000 53.400 101.400 54.550 ;
        RECT 102.000 53.400 102.400 54.550 ;
        RECT 103.000 53.400 103.400 54.550 ;
        RECT 104.000 53.400 104.400 54.550 ;
        RECT 105.000 53.400 105.400 54.550 ;
        RECT 106.000 53.400 106.400 54.550 ;
        RECT 107.000 53.400 107.900 54.550 ;
        RECT 57.750 50.350 58.450 53.250 ;
        RECT 59.050 50.350 59.350 53.250 ;
        RECT 59.950 50.350 60.250 53.250 ;
        RECT 60.850 50.350 61.150 53.250 ;
        RECT 61.750 50.350 62.050 53.250 ;
        RECT 62.650 50.350 62.950 53.250 ;
        RECT 63.550 50.350 63.850 53.250 ;
        RECT 64.450 50.350 64.750 53.250 ;
        RECT 65.350 50.350 65.650 53.250 ;
        RECT 66.250 50.350 66.550 53.250 ;
        RECT 67.150 50.350 67.450 53.250 ;
        RECT 68.050 50.350 68.350 53.250 ;
        RECT 68.950 50.350 69.250 53.250 ;
        RECT 69.850 50.350 70.150 53.250 ;
        RECT 70.750 50.350 71.050 53.250 ;
        RECT 71.650 50.350 71.950 53.250 ;
        RECT 72.550 50.350 72.850 53.250 ;
        RECT 73.450 50.350 73.750 53.250 ;
        RECT 74.350 50.350 75.050 53.250 ;
        RECT 101.100 53.200 101.300 53.400 ;
        RECT 103.100 53.200 103.300 53.400 ;
        RECT 77.950 52.450 78.350 52.850 ;
        RECT 78.550 52.450 78.950 52.850 ;
        RECT 79.150 52.450 79.550 52.850 ;
        RECT 101.000 52.800 103.400 53.200 ;
        RECT 77.050 51.350 77.800 52.250 ;
        RECT 78.050 51.350 78.350 52.250 ;
        RECT 78.600 51.350 78.900 52.250 ;
        RECT 79.150 51.350 79.450 52.250 ;
        RECT 79.700 51.350 80.400 52.250 ;
        RECT 95.700 52.200 96.300 52.250 ;
        RECT 102.950 52.200 103.400 52.800 ;
        RECT 95.700 51.870 96.470 52.200 ;
        RECT 102.670 51.870 103.400 52.200 ;
        RECT 95.700 51.850 96.300 51.870 ;
        RECT 102.800 51.850 103.400 51.870 ;
        RECT 77.450 50.750 77.850 51.150 ;
        RECT 78.550 50.750 78.950 51.150 ;
        RECT 79.700 50.750 80.000 51.150 ;
        RECT 58.200 50.150 58.400 50.350 ;
        RECT 60.000 50.150 60.200 50.350 ;
        RECT 61.800 50.150 62.000 50.350 ;
        RECT 63.600 50.150 63.800 50.350 ;
        RECT 65.400 50.150 65.600 50.350 ;
        RECT 67.200 50.150 67.400 50.350 ;
        RECT 69.000 50.150 69.200 50.350 ;
        RECT 70.800 50.150 71.000 50.350 ;
        RECT 72.600 50.150 72.800 50.350 ;
        RECT 74.400 50.150 74.600 50.350 ;
        RECT 115.165 50.300 115.335 57.505 ;
        RECT 116.120 54.820 116.470 56.980 ;
        RECT 58.100 49.750 58.500 50.150 ;
        RECT 59.900 49.750 60.300 50.150 ;
        RECT 61.700 49.750 62.100 50.150 ;
        RECT 63.500 49.750 63.900 50.150 ;
        RECT 65.300 49.750 65.700 50.150 ;
        RECT 67.100 49.750 67.500 50.150 ;
        RECT 68.900 49.750 69.300 50.150 ;
        RECT 70.700 49.750 71.100 50.150 ;
        RECT 72.500 49.750 72.900 50.150 ;
        RECT 74.300 49.750 74.700 50.150 ;
        RECT 115.050 49.900 115.450 50.300 ;
        RECT 59.030 48.450 59.320 48.800 ;
        RECT 59.580 48.450 59.870 48.800 ;
        RECT 60.130 48.450 60.420 48.800 ;
        RECT 60.680 48.450 60.970 48.800 ;
        RECT 61.230 48.450 61.520 48.800 ;
        RECT 61.780 48.450 62.070 48.800 ;
        RECT 62.330 48.450 62.620 48.800 ;
        RECT 62.880 48.450 63.170 48.800 ;
        RECT 63.430 48.450 63.720 48.800 ;
        RECT 63.980 48.450 64.270 48.800 ;
        RECT 68.530 48.450 68.820 48.800 ;
        RECT 69.080 48.450 69.370 48.800 ;
        RECT 69.630 48.450 69.920 48.800 ;
        RECT 70.180 48.450 70.470 48.800 ;
        RECT 70.730 48.450 71.020 48.800 ;
        RECT 71.280 48.450 71.570 48.800 ;
        RECT 71.830 48.450 72.120 48.800 ;
        RECT 72.380 48.450 72.670 48.800 ;
        RECT 72.930 48.450 73.220 48.800 ;
        RECT 73.480 48.450 73.770 48.800 ;
        RECT 57.800 47.350 58.500 48.250 ;
        RECT 58.750 47.350 59.050 48.250 ;
        RECT 59.300 47.350 59.600 48.250 ;
        RECT 59.850 47.350 60.150 48.250 ;
        RECT 60.400 47.350 60.700 48.250 ;
        RECT 60.950 47.350 61.250 48.250 ;
        RECT 61.500 47.350 61.800 48.250 ;
        RECT 62.050 47.350 62.350 48.250 ;
        RECT 62.600 47.350 62.900 48.250 ;
        RECT 63.150 47.350 63.450 48.250 ;
        RECT 63.700 47.350 64.000 48.250 ;
        RECT 64.250 47.350 64.550 48.250 ;
        RECT 64.800 47.350 65.500 48.250 ;
        RECT 67.300 47.350 68.000 48.250 ;
        RECT 68.250 47.350 68.550 48.250 ;
        RECT 68.800 47.350 69.100 48.250 ;
        RECT 69.350 47.350 69.650 48.250 ;
        RECT 69.900 47.350 70.200 48.250 ;
        RECT 70.450 47.350 70.750 48.250 ;
        RECT 71.000 47.350 71.300 48.250 ;
        RECT 71.550 47.350 71.850 48.250 ;
        RECT 72.100 47.350 72.400 48.250 ;
        RECT 72.650 47.350 72.950 48.250 ;
        RECT 73.200 47.350 73.500 48.250 ;
        RECT 73.750 47.350 74.050 48.250 ;
        RECT 74.300 47.350 75.000 48.250 ;
        RECT 115.165 48.135 115.335 49.900 ;
        RECT 116.120 48.660 116.470 50.820 ;
        RECT 117.255 48.135 117.425 57.505 ;
        RECT 115.165 47.965 117.425 48.135 ;
        RECT 58.150 46.750 58.550 47.150 ;
        RECT 64.750 46.750 65.150 47.150 ;
        RECT 67.650 46.750 68.050 47.150 ;
        RECT 74.250 46.750 74.650 47.150 ;
        RECT 66.250 41.150 66.650 41.550 ;
        RECT 67.350 41.150 67.750 41.550 ;
        RECT 68.850 41.150 69.250 41.550 ;
        RECT 70.000 41.150 70.400 41.550 ;
        RECT 70.750 41.150 71.150 41.550 ;
        RECT 71.850 41.150 72.250 41.550 ;
        RECT 73.350 41.150 73.750 41.550 ;
        RECT 74.450 41.150 74.850 41.550 ;
        RECT 76.450 41.150 76.850 41.550 ;
        RECT 78.100 41.150 78.500 41.550 ;
        RECT 79.750 41.150 80.150 41.550 ;
        RECT 81.950 41.150 82.350 41.550 ;
        RECT 85.850 41.150 86.250 41.550 ;
        RECT 89.250 41.150 89.650 41.550 ;
        RECT 115.450 41.450 116.000 42.000 ;
        RECT 66.350 40.400 66.550 41.150 ;
        RECT 67.450 40.400 67.650 41.150 ;
        RECT 68.950 40.400 69.150 41.150 ;
        RECT 70.100 40.400 70.300 41.150 ;
        RECT 70.850 40.400 71.050 41.150 ;
        RECT 71.950 40.400 72.150 41.150 ;
        RECT 73.450 40.400 73.650 41.150 ;
        RECT 74.550 40.400 74.750 41.150 ;
        RECT 76.550 40.400 76.750 41.150 ;
        RECT 78.200 40.400 78.400 41.150 ;
        RECT 79.850 40.400 80.050 41.150 ;
        RECT 82.050 40.400 82.250 41.150 ;
        RECT 84.500 40.600 84.900 41.000 ;
        RECT 85.950 40.400 86.150 41.150 ;
        RECT 87.650 40.600 88.050 41.000 ;
        RECT 89.350 40.400 89.550 41.150 ;
        RECT 65.900 39.500 66.600 40.400 ;
        RECT 66.850 39.500 67.150 40.400 ;
        RECT 67.400 39.500 67.700 40.400 ;
        RECT 68.900 39.500 69.200 40.400 ;
        RECT 69.450 39.500 69.750 40.400 ;
        RECT 70.000 39.500 71.100 40.400 ;
        RECT 71.350 39.500 71.650 40.400 ;
        RECT 71.900 39.500 72.200 40.400 ;
        RECT 73.400 39.500 73.700 40.400 ;
        RECT 73.950 39.500 74.250 40.400 ;
        RECT 74.500 39.500 75.200 40.400 ;
        RECT 75.950 39.500 76.250 40.400 ;
        RECT 76.500 39.500 77.200 40.400 ;
        RECT 77.600 39.500 77.900 40.400 ;
        RECT 78.150 39.500 78.850 40.400 ;
        RECT 79.250 39.500 79.550 40.400 ;
        RECT 79.800 39.500 80.500 40.400 ;
        RECT 81.450 39.500 82.350 40.400 ;
        RECT 82.600 39.500 83.000 40.400 ;
        RECT 83.900 39.500 84.300 40.400 ;
        RECT 84.550 39.500 84.950 40.400 ;
        RECT 85.350 39.500 86.250 40.400 ;
        RECT 86.500 39.500 86.900 40.400 ;
        RECT 87.300 39.500 87.700 40.400 ;
        RECT 87.950 39.500 88.350 40.400 ;
        RECT 88.750 39.500 89.650 40.400 ;
        RECT 89.900 39.500 90.300 40.400 ;
        RECT 96.700 40.350 97.100 40.750 ;
        RECT 111.900 40.350 112.300 40.750 ;
        RECT 65.650 38.700 66.050 39.100 ;
        RECT 66.850 38.700 67.050 39.500 ;
        RECT 67.300 39.100 67.700 39.300 ;
        RECT 67.300 38.900 68.700 39.100 ;
        RECT 66.850 38.500 67.650 38.700 ;
        RECT 67.450 38.300 67.650 38.500 ;
        RECT 65.900 36.400 66.600 38.300 ;
        RECT 66.850 36.400 67.150 38.300 ;
        RECT 67.400 36.650 67.700 38.300 ;
        RECT 67.900 36.650 68.300 36.800 ;
        RECT 67.400 36.400 68.300 36.650 ;
        RECT 68.500 36.600 68.700 38.900 ;
        RECT 69.500 38.700 69.700 39.500 ;
        RECT 68.950 38.500 69.700 38.700 ;
        RECT 69.900 38.700 70.300 38.900 ;
        RECT 71.350 38.700 71.550 39.500 ;
        RECT 71.800 39.100 72.200 39.300 ;
        RECT 71.800 38.900 73.200 39.100 ;
        RECT 69.900 38.500 72.150 38.700 ;
        RECT 68.950 38.300 69.150 38.500 ;
        RECT 71.950 38.300 72.150 38.500 ;
        RECT 68.900 36.600 69.200 38.300 ;
        RECT 68.500 36.400 69.200 36.600 ;
        RECT 69.450 36.400 69.750 38.300 ;
        RECT 70.000 36.400 71.100 38.300 ;
        RECT 71.350 36.400 71.650 38.300 ;
        RECT 71.900 36.650 72.200 38.300 ;
        RECT 72.400 36.650 72.800 36.800 ;
        RECT 71.900 36.400 72.800 36.650 ;
        RECT 73.000 36.600 73.200 38.900 ;
        RECT 74.000 38.700 74.200 39.500 ;
        RECT 75.950 39.050 76.150 39.500 ;
        RECT 77.600 39.050 77.800 39.500 ;
        RECT 79.250 39.050 79.450 39.500 ;
        RECT 73.450 38.500 74.200 38.700 ;
        RECT 75.250 38.650 76.150 39.050 ;
        RECT 77.300 38.650 77.800 39.050 ;
        RECT 78.950 38.650 79.450 39.050 ;
        RECT 80.400 38.650 80.800 39.050 ;
        RECT 81.150 38.700 81.550 39.100 ;
        RECT 82.700 38.700 82.900 39.500 ;
        RECT 84.000 38.700 84.200 39.500 ;
        RECT 73.450 38.300 73.650 38.500 ;
        RECT 75.950 38.300 76.150 38.650 ;
        RECT 77.600 38.300 77.800 38.650 ;
        RECT 79.250 38.300 79.450 38.650 ;
        RECT 82.700 38.500 84.200 38.700 ;
        RECT 82.700 38.300 82.900 38.500 ;
        RECT 84.000 38.300 84.200 38.500 ;
        RECT 84.650 38.950 84.850 39.500 ;
        RECT 86.700 39.350 86.900 39.500 ;
        RECT 86.700 39.000 87.100 39.350 ;
        RECT 84.650 38.550 85.150 38.950 ;
        RECT 84.650 38.300 84.850 38.550 ;
        RECT 86.700 38.300 86.900 39.000 ;
        RECT 87.400 38.300 87.600 39.500 ;
        RECT 88.050 39.100 88.250 39.500 ;
        RECT 90.000 39.300 90.200 39.500 ;
        RECT 90.000 39.100 90.400 39.300 ;
        RECT 88.050 38.900 90.400 39.100 ;
        RECT 88.050 38.300 88.250 38.900 ;
        RECT 73.400 36.600 73.700 38.300 ;
        RECT 73.000 36.400 73.700 36.600 ;
        RECT 73.950 36.400 74.250 38.300 ;
        RECT 74.500 36.400 75.200 38.300 ;
        RECT 75.950 36.400 76.250 38.300 ;
        RECT 76.500 36.400 77.200 38.300 ;
        RECT 77.600 36.400 77.900 38.300 ;
        RECT 78.150 36.400 78.850 38.300 ;
        RECT 79.250 36.400 79.550 38.300 ;
        RECT 79.800 36.400 80.500 38.300 ;
        RECT 81.450 36.400 82.350 38.300 ;
        RECT 82.600 36.400 83.000 38.300 ;
        RECT 83.900 36.400 84.300 38.300 ;
        RECT 84.550 36.400 84.950 38.300 ;
        RECT 85.350 36.400 86.250 38.300 ;
        RECT 86.500 36.400 86.900 38.300 ;
        RECT 87.300 36.400 87.700 38.300 ;
        RECT 87.950 36.400 88.350 38.300 ;
        RECT 96.200 38.250 97.100 40.150 ;
        RECT 97.800 38.250 98.200 40.150 ;
        RECT 98.900 37.700 99.300 40.150 ;
        RECT 100.000 38.250 100.400 40.150 ;
        RECT 101.100 38.250 102.500 40.150 ;
        RECT 103.200 38.250 103.600 40.150 ;
        RECT 104.300 38.250 104.700 40.150 ;
        RECT 105.400 38.250 105.800 40.150 ;
        RECT 106.500 38.250 107.900 40.150 ;
        RECT 108.600 38.250 109.000 40.150 ;
        RECT 109.700 38.250 110.100 40.150 ;
        RECT 110.800 38.250 111.200 40.150 ;
        RECT 111.900 38.250 112.800 40.150 ;
        RECT 101.600 37.650 102.000 38.250 ;
        RECT 107.000 37.650 107.400 38.250 ;
        RECT 109.050 37.500 109.450 37.900 ;
        RECT 110.350 37.500 110.750 37.900 ;
        RECT 113.700 37.500 114.250 38.050 ;
        RECT 66.350 35.650 66.550 36.400 ;
        RECT 68.500 36.200 68.700 36.400 ;
        RECT 68.500 35.800 68.900 36.200 ;
        RECT 70.050 35.650 70.250 36.400 ;
        RECT 70.850 35.650 71.050 36.400 ;
        RECT 74.550 35.650 74.750 36.400 ;
        RECT 76.650 35.650 76.850 36.400 ;
        RECT 78.200 35.650 78.400 36.400 ;
        RECT 79.850 35.650 80.050 36.400 ;
        RECT 82.050 35.650 82.250 36.400 ;
        RECT 84.100 35.850 84.500 36.200 ;
        RECT 85.950 35.650 86.150 36.400 ;
        RECT 87.400 36.200 87.600 36.400 ;
        RECT 87.300 35.800 87.700 36.200 ;
        RECT 66.250 35.250 66.650 35.650 ;
        RECT 69.950 35.250 70.350 35.650 ;
        RECT 70.750 35.250 71.150 35.650 ;
        RECT 74.450 35.250 74.850 35.650 ;
        RECT 75.700 35.250 76.100 35.650 ;
        RECT 76.650 35.250 77.450 35.650 ;
        RECT 78.100 35.250 78.500 35.650 ;
        RECT 79.750 35.250 80.150 35.650 ;
        RECT 81.950 35.250 82.350 35.650 ;
        RECT 83.900 35.250 84.300 35.650 ;
        RECT 85.850 35.250 86.250 35.650 ;
        RECT 89.250 35.250 89.650 35.650 ;
        RECT 66.350 34.500 66.550 35.250 ;
        RECT 70.050 34.500 70.250 35.250 ;
        RECT 70.850 34.500 71.050 35.250 ;
        RECT 74.550 34.500 74.750 35.250 ;
        RECT 75.800 34.500 76.000 35.250 ;
        RECT 76.250 34.700 76.650 35.050 ;
        RECT 77.150 34.500 77.350 35.250 ;
        RECT 78.250 34.500 78.450 35.250 ;
        RECT 79.900 34.500 80.100 35.250 ;
        RECT 82.050 34.500 82.250 35.250 ;
        RECT 84.000 34.500 84.200 35.250 ;
        RECT 85.950 34.500 86.150 35.250 ;
        RECT 89.350 34.500 89.550 35.250 ;
        RECT 101.000 34.850 101.400 35.250 ;
        RECT 104.800 34.650 105.200 35.250 ;
        RECT 106.850 35.000 107.250 35.400 ;
        RECT 110.350 35.000 110.750 35.400 ;
        RECT 113.700 34.850 114.250 35.400 ;
        RECT 65.900 32.600 66.600 34.500 ;
        RECT 66.850 32.600 67.150 34.500 ;
        RECT 67.400 34.250 68.300 34.500 ;
        RECT 67.400 32.600 67.700 34.250 ;
        RECT 67.900 34.100 68.300 34.250 ;
        RECT 68.500 34.300 69.200 34.500 ;
        RECT 67.450 32.400 67.650 32.600 ;
        RECT 66.850 32.200 67.650 32.400 ;
        RECT 65.650 31.800 66.050 32.200 ;
        RECT 66.850 31.400 67.050 32.200 ;
        RECT 68.500 32.000 68.700 34.300 ;
        RECT 68.900 32.600 69.200 34.300 ;
        RECT 69.450 32.600 69.750 34.500 ;
        RECT 70.000 32.600 71.100 34.500 ;
        RECT 71.350 32.600 71.650 34.500 ;
        RECT 71.900 34.250 72.800 34.500 ;
        RECT 71.900 32.600 72.200 34.250 ;
        RECT 72.400 34.100 72.800 34.250 ;
        RECT 73.000 34.300 73.700 34.500 ;
        RECT 68.950 32.400 69.150 32.600 ;
        RECT 71.950 32.400 72.150 32.600 ;
        RECT 68.950 32.200 69.700 32.400 ;
        RECT 67.300 31.800 68.700 32.000 ;
        RECT 67.300 31.600 67.700 31.800 ;
        RECT 65.900 30.500 66.600 31.400 ;
        RECT 66.850 30.500 67.150 31.400 ;
        RECT 67.400 30.500 67.700 31.400 ;
        RECT 66.350 29.750 66.550 30.500 ;
        RECT 67.450 29.750 67.650 30.500 ;
        RECT 68.500 30.300 68.700 31.800 ;
        RECT 69.500 31.400 69.700 32.200 ;
        RECT 69.900 32.200 72.150 32.400 ;
        RECT 69.900 32.000 70.300 32.200 ;
        RECT 71.350 31.400 71.550 32.200 ;
        RECT 73.000 32.000 73.200 34.300 ;
        RECT 73.400 32.600 73.700 34.300 ;
        RECT 73.950 32.600 74.250 34.500 ;
        RECT 74.500 32.600 75.200 34.500 ;
        RECT 75.600 32.600 76.300 34.500 ;
        RECT 76.550 32.600 76.850 34.500 ;
        RECT 77.100 32.600 77.400 34.500 ;
        RECT 77.800 32.600 78.500 34.500 ;
        RECT 78.750 32.600 79.050 34.500 ;
        RECT 79.450 32.600 80.150 34.500 ;
        RECT 80.400 32.600 80.700 34.500 ;
        RECT 81.450 32.600 82.350 34.500 ;
        RECT 82.600 32.600 83.000 34.500 ;
        RECT 83.400 32.600 84.300 34.500 ;
        RECT 84.550 32.600 84.950 34.500 ;
        RECT 85.350 32.600 86.250 34.500 ;
        RECT 86.500 32.600 86.900 34.500 ;
        RECT 87.300 32.600 87.700 34.500 ;
        RECT 87.950 32.600 88.350 34.500 ;
        RECT 88.750 32.600 89.650 34.500 ;
        RECT 89.900 32.600 90.300 34.500 ;
        RECT 97.200 32.750 98.100 34.650 ;
        RECT 98.800 32.750 99.200 34.650 ;
        RECT 99.900 32.750 100.300 34.650 ;
        RECT 101.000 32.750 101.400 34.650 ;
        RECT 102.100 32.750 102.500 34.650 ;
        RECT 103.200 32.750 103.600 34.650 ;
        RECT 104.300 32.750 105.700 34.650 ;
        RECT 106.400 32.750 106.800 34.650 ;
        RECT 107.500 32.750 107.900 34.650 ;
        RECT 108.600 32.750 109.000 34.650 ;
        RECT 109.700 32.750 110.100 34.650 ;
        RECT 110.800 32.750 111.200 34.650 ;
        RECT 111.900 32.750 112.800 34.650 ;
        RECT 73.450 32.400 73.650 32.600 ;
        RECT 73.450 32.200 74.200 32.400 ;
        RECT 71.800 31.800 73.200 32.000 ;
        RECT 71.800 31.600 72.200 31.800 ;
        RECT 74.000 31.400 74.200 32.200 ;
        RECT 76.600 32.250 76.800 32.600 ;
        RECT 78.850 32.250 79.050 32.600 ;
        RECT 80.500 32.250 80.700 32.600 ;
        RECT 76.600 32.050 77.700 32.250 ;
        RECT 75.150 31.650 75.550 32.050 ;
        RECT 77.150 31.850 77.700 32.050 ;
        RECT 78.850 31.850 79.350 32.250 ;
        RECT 80.500 31.850 81.000 32.250 ;
        RECT 82.800 32.150 83.000 32.600 ;
        RECT 84.100 32.150 84.500 32.250 ;
        RECT 77.150 31.400 77.350 31.850 ;
        RECT 78.850 31.400 79.050 31.850 ;
        RECT 80.500 31.400 80.700 31.850 ;
        RECT 81.250 31.700 81.650 32.100 ;
        RECT 82.800 31.950 84.500 32.150 ;
        RECT 82.800 31.400 83.000 31.950 ;
        RECT 84.100 31.850 84.500 31.950 ;
        RECT 84.750 32.000 84.950 32.600 ;
        RECT 86.700 32.400 86.900 32.600 ;
        RECT 86.700 32.000 87.100 32.400 ;
        RECT 84.750 31.800 86.450 32.000 ;
        RECT 84.750 31.400 84.950 31.800 ;
        RECT 86.050 31.600 86.450 31.800 ;
        RECT 86.700 31.400 86.900 32.000 ;
        RECT 87.400 31.400 87.600 32.600 ;
        RECT 88.050 31.800 88.250 32.600 ;
        RECT 88.450 32.000 88.850 32.400 ;
        RECT 90.000 32.000 90.200 32.600 ;
        RECT 97.700 32.150 98.100 32.550 ;
        RECT 111.900 32.150 112.300 32.550 ;
        RECT 90.000 31.800 90.400 32.000 ;
        RECT 88.050 31.600 90.400 31.800 ;
        RECT 88.050 31.400 88.250 31.600 ;
        RECT 68.900 30.500 69.200 31.400 ;
        RECT 69.450 30.500 69.750 31.400 ;
        RECT 70.000 30.500 71.100 31.400 ;
        RECT 71.350 30.500 71.650 31.400 ;
        RECT 71.900 30.500 72.200 31.400 ;
        RECT 73.400 30.500 73.700 31.400 ;
        RECT 73.950 30.500 74.250 31.400 ;
        RECT 74.500 30.500 75.200 31.400 ;
        RECT 75.600 30.500 76.300 31.400 ;
        RECT 76.550 30.500 76.850 31.400 ;
        RECT 77.100 30.500 77.400 31.400 ;
        RECT 77.800 30.500 78.500 31.400 ;
        RECT 78.750 30.500 79.050 31.400 ;
        RECT 79.450 30.500 80.150 31.400 ;
        RECT 80.400 30.500 80.700 31.400 ;
        RECT 81.550 30.500 82.350 31.400 ;
        RECT 82.600 30.500 83.000 31.400 ;
        RECT 83.500 30.500 84.300 31.400 ;
        RECT 84.550 30.500 84.950 31.400 ;
        RECT 85.450 30.500 86.250 31.400 ;
        RECT 86.500 30.500 86.900 31.400 ;
        RECT 87.300 30.500 87.700 31.400 ;
        RECT 87.950 30.500 88.350 31.400 ;
        RECT 68.300 29.900 68.700 30.300 ;
        RECT 68.950 29.750 69.150 30.500 ;
        RECT 70.050 29.750 70.250 30.500 ;
        RECT 70.850 29.750 71.050 30.500 ;
        RECT 71.950 29.750 72.150 30.500 ;
        RECT 73.450 29.750 73.650 30.500 ;
        RECT 74.550 29.750 74.750 30.500 ;
        RECT 76.050 29.750 76.250 30.500 ;
        RECT 76.900 29.900 77.300 30.300 ;
        RECT 78.250 29.750 78.450 30.500 ;
        RECT 79.900 29.750 80.100 30.500 ;
        RECT 82.050 29.750 82.250 30.500 ;
        RECT 84.000 29.750 84.200 30.500 ;
        RECT 85.950 29.750 86.150 30.500 ;
        RECT 87.400 30.300 87.600 30.500 ;
        RECT 87.300 29.900 87.700 30.300 ;
        RECT 66.250 29.350 66.650 29.750 ;
        RECT 67.350 29.350 67.750 29.750 ;
        RECT 68.850 29.350 69.250 29.750 ;
        RECT 69.950 29.350 70.350 29.750 ;
        RECT 70.750 29.350 71.150 29.750 ;
        RECT 71.850 29.350 72.250 29.750 ;
        RECT 73.350 29.350 73.750 29.750 ;
        RECT 74.450 29.350 74.850 29.750 ;
        RECT 75.950 29.350 76.350 29.750 ;
        RECT 78.150 29.350 78.550 29.750 ;
        RECT 79.800 29.350 80.200 29.750 ;
        RECT 81.950 29.350 82.350 29.750 ;
        RECT 83.900 29.350 84.300 29.750 ;
        RECT 85.850 29.350 86.250 29.750 ;
        RECT 114.900 28.950 115.450 29.500 ;
        RECT 117.900 27.650 118.300 27.750 ;
        RECT 120.500 27.650 120.900 27.750 ;
        RECT 123.100 27.650 123.500 27.750 ;
        RECT 125.700 27.650 126.100 27.750 ;
        RECT 115.450 27.450 126.600 27.650 ;
        RECT 63.300 18.350 63.700 18.750 ;
        RECT 65.400 18.350 65.800 18.750 ;
        RECT 68.750 18.350 69.150 18.750 ;
        RECT 71.600 18.350 72.000 18.750 ;
        RECT 75.350 18.350 75.750 18.750 ;
        RECT 77.500 18.350 77.900 18.750 ;
        RECT 79.700 18.350 80.100 18.750 ;
        RECT 80.950 18.350 81.350 18.750 ;
        RECT 82.050 18.350 82.450 18.750 ;
        RECT 84.400 18.350 84.800 18.750 ;
        RECT 86.600 18.350 87.000 18.750 ;
        RECT 89.700 18.350 90.100 18.750 ;
        RECT 91.400 18.350 91.800 18.750 ;
        RECT 93.200 18.350 93.600 18.750 ;
        RECT 96.200 18.350 96.600 18.750 ;
        RECT 97.900 18.350 98.300 18.750 ;
        RECT 99.700 18.350 100.100 18.750 ;
        RECT 102.700 18.350 103.100 18.750 ;
        RECT 104.400 18.350 104.800 18.750 ;
        RECT 106.200 18.350 106.600 18.750 ;
        RECT 109.200 18.350 109.600 18.750 ;
        RECT 110.900 18.350 111.300 18.750 ;
        RECT 112.700 18.350 113.100 18.750 ;
        RECT 63.400 17.600 63.600 18.350 ;
        RECT 64.900 17.800 65.300 18.200 ;
        RECT 65.500 17.600 65.700 18.350 ;
        RECT 65.900 17.800 66.250 18.200 ;
        RECT 66.050 17.600 66.250 17.800 ;
        RECT 66.450 17.700 66.850 18.100 ;
        RECT 68.850 17.600 69.050 18.350 ;
        RECT 70.500 17.800 70.900 18.200 ;
        RECT 71.200 17.800 71.500 18.200 ;
        RECT 71.700 17.600 71.900 18.350 ;
        RECT 75.450 17.600 75.650 18.350 ;
        RECT 77.000 17.800 77.400 18.200 ;
        RECT 77.600 17.600 77.800 18.350 ;
        RECT 78.100 17.800 78.500 18.200 ;
        RECT 78.100 17.600 78.300 17.800 ;
        RECT 79.800 17.600 80.000 18.350 ;
        RECT 81.050 17.600 81.250 18.350 ;
        RECT 82.150 17.600 82.350 18.350 ;
        RECT 83.750 17.850 84.150 18.200 ;
        RECT 83.950 17.600 84.150 17.850 ;
        RECT 84.500 17.600 84.700 18.350 ;
        RECT 85.800 17.850 86.200 18.200 ;
        RECT 86.700 17.600 86.900 18.350 ;
        RECT 89.800 17.600 90.000 18.350 ;
        RECT 91.500 17.600 91.700 18.350 ;
        RECT 93.300 17.600 93.500 18.350 ;
        RECT 95.550 17.800 95.950 18.200 ;
        RECT 95.750 17.600 95.950 17.800 ;
        RECT 96.300 17.600 96.500 18.350 ;
        RECT 98.000 17.600 98.200 18.350 ;
        RECT 98.450 17.800 98.850 18.200 ;
        RECT 99.800 17.600 100.000 18.350 ;
        RECT 102.050 17.800 102.450 18.200 ;
        RECT 102.250 17.600 102.450 17.800 ;
        RECT 102.800 17.600 103.000 18.350 ;
        RECT 104.500 17.600 104.700 18.350 ;
        RECT 104.950 17.800 105.350 18.200 ;
        RECT 106.300 17.600 106.500 18.350 ;
        RECT 108.550 17.800 108.950 18.200 ;
        RECT 108.750 17.600 108.950 17.800 ;
        RECT 109.300 17.600 109.500 18.350 ;
        RECT 111.000 17.600 111.200 18.350 ;
        RECT 111.450 17.800 111.850 18.200 ;
        RECT 112.800 17.600 113.000 18.350 ;
        RECT 61.500 17.500 61.900 17.600 ;
        RECT 62.800 17.500 63.100 17.600 ;
        RECT 61.500 17.300 63.100 17.500 ;
        RECT 61.500 17.200 61.900 17.300 ;
        RECT 62.800 17.200 63.100 17.300 ;
        RECT 63.350 17.200 64.050 17.600 ;
        RECT 64.900 17.500 65.200 17.600 ;
        RECT 64.250 17.300 65.200 17.500 ;
        RECT 61.600 16.750 61.800 17.200 ;
        RECT 61.200 16.350 61.800 16.750 ;
        RECT 61.600 16.000 61.800 16.350 ;
        RECT 62.250 16.400 62.650 16.600 ;
        RECT 64.250 16.400 64.450 17.300 ;
        RECT 64.900 17.200 65.200 17.300 ;
        RECT 65.450 17.200 65.750 17.600 ;
        RECT 66.000 17.200 66.300 17.600 ;
        RECT 68.250 17.500 68.550 17.600 ;
        RECT 67.150 17.300 68.550 17.500 ;
        RECT 66.050 17.000 66.250 17.200 ;
        RECT 62.250 16.200 64.450 16.400 ;
        RECT 63.150 16.000 63.350 16.200 ;
        RECT 64.250 16.000 64.450 16.200 ;
        RECT 64.700 16.800 66.250 17.000 ;
        RECT 64.700 16.000 64.900 16.800 ;
        RECT 67.150 16.600 67.350 17.300 ;
        RECT 68.250 17.200 68.550 17.300 ;
        RECT 68.800 17.200 69.100 17.600 ;
        RECT 69.350 17.200 69.650 17.600 ;
        RECT 70.450 17.200 70.750 17.600 ;
        RECT 71.000 17.200 71.300 17.600 ;
        RECT 71.550 17.200 71.900 17.600 ;
        RECT 72.100 17.200 72.400 17.600 ;
        RECT 73.650 17.500 74.050 17.600 ;
        RECT 74.850 17.500 75.150 17.600 ;
        RECT 73.650 17.300 75.150 17.500 ;
        RECT 73.650 17.200 74.050 17.300 ;
        RECT 74.850 17.200 75.150 17.300 ;
        RECT 75.400 17.200 76.100 17.600 ;
        RECT 76.950 17.500 77.250 17.600 ;
        RECT 76.300 17.300 77.250 17.500 ;
        RECT 67.850 16.600 68.250 17.000 ;
        RECT 65.150 16.500 65.550 16.600 ;
        RECT 66.850 16.500 67.350 16.600 ;
        RECT 65.150 16.300 67.350 16.500 ;
        RECT 65.150 16.200 65.550 16.300 ;
        RECT 66.850 16.200 67.350 16.300 ;
        RECT 68.050 16.400 68.250 16.600 ;
        RECT 69.350 16.400 69.550 17.200 ;
        RECT 69.850 17.000 70.250 17.200 ;
        RECT 70.500 17.000 70.700 17.200 ;
        RECT 72.150 17.000 72.350 17.200 ;
        RECT 69.850 16.800 73.150 17.000 ;
        RECT 68.050 16.200 69.550 16.400 ;
        RECT 69.750 16.200 70.150 16.550 ;
        RECT 70.500 16.200 71.800 16.400 ;
        RECT 72.350 16.200 72.750 16.550 ;
        RECT 67.150 16.000 67.350 16.200 ;
        RECT 68.250 16.000 68.450 16.200 ;
        RECT 69.350 16.000 69.550 16.200 ;
        RECT 70.500 16.000 70.700 16.200 ;
        RECT 71.600 16.000 71.800 16.200 ;
        RECT 72.950 16.000 73.150 16.800 ;
        RECT 61.600 15.600 62.300 16.000 ;
        RECT 62.550 15.600 62.850 16.000 ;
        RECT 63.100 15.600 63.400 16.000 ;
        RECT 63.650 15.600 63.950 16.000 ;
        RECT 64.200 15.600 64.500 16.000 ;
        RECT 64.700 15.700 65.200 16.000 ;
        RECT 64.900 15.600 65.200 15.700 ;
        RECT 65.450 15.600 65.750 16.000 ;
        RECT 66.000 15.600 66.300 16.000 ;
        RECT 67.150 15.600 67.450 16.000 ;
        RECT 67.700 15.600 68.000 16.000 ;
        RECT 68.250 15.600 68.550 16.000 ;
        RECT 68.800 15.600 69.100 16.000 ;
        RECT 69.350 15.600 69.650 16.000 ;
        RECT 70.450 15.600 70.750 16.000 ;
        RECT 71.000 15.600 71.300 16.000 ;
        RECT 71.550 15.600 71.850 16.000 ;
        RECT 72.100 15.600 72.400 16.000 ;
        RECT 72.650 15.700 73.150 16.000 ;
        RECT 73.850 16.000 74.050 17.200 ;
        RECT 74.300 16.400 74.700 16.550 ;
        RECT 76.300 16.400 76.500 17.300 ;
        RECT 76.950 17.200 77.250 17.300 ;
        RECT 77.500 17.200 77.800 17.600 ;
        RECT 78.050 17.200 78.350 17.600 ;
        RECT 79.200 17.200 79.500 17.600 ;
        RECT 79.750 17.200 80.050 17.600 ;
        RECT 80.300 17.200 80.600 17.600 ;
        RECT 81.000 17.200 81.300 17.600 ;
        RECT 81.550 17.200 81.850 17.600 ;
        RECT 82.100 17.200 82.400 17.600 ;
        RECT 83.900 17.500 84.200 17.600 ;
        RECT 82.800 17.300 84.200 17.500 ;
        RECT 78.100 17.000 78.300 17.200 ;
        RECT 74.300 16.200 76.500 16.400 ;
        RECT 75.200 16.000 75.400 16.200 ;
        RECT 76.300 16.000 76.500 16.200 ;
        RECT 76.750 16.800 78.300 17.000 ;
        RECT 78.550 17.000 78.950 17.200 ;
        RECT 79.250 17.000 79.450 17.200 ;
        RECT 80.350 17.000 80.550 17.200 ;
        RECT 78.550 16.800 80.550 17.000 ;
        RECT 76.750 16.000 76.950 16.800 ;
        RECT 77.200 16.500 77.600 16.600 ;
        RECT 78.250 16.500 78.650 16.550 ;
        RECT 77.200 16.300 78.650 16.500 ;
        RECT 77.200 16.200 77.600 16.300 ;
        RECT 78.250 16.200 78.650 16.300 ;
        RECT 73.850 15.700 74.350 16.000 ;
        RECT 72.650 15.600 72.950 15.700 ;
        RECT 74.050 15.600 74.350 15.700 ;
        RECT 74.600 15.600 74.900 16.000 ;
        RECT 75.150 15.600 75.450 16.000 ;
        RECT 75.700 15.600 76.000 16.000 ;
        RECT 76.250 15.600 76.550 16.000 ;
        RECT 76.750 15.700 77.250 16.000 ;
        RECT 76.950 15.600 77.250 15.700 ;
        RECT 77.500 15.600 77.800 16.000 ;
        RECT 78.050 15.600 78.750 16.000 ;
        RECT 78.950 15.900 79.150 16.800 ;
        RECT 81.600 16.650 81.800 17.200 ;
        RECT 82.800 16.850 83.000 17.300 ;
        RECT 83.900 17.200 84.200 17.300 ;
        RECT 84.450 17.200 84.750 17.600 ;
        RECT 85.000 17.200 85.300 17.600 ;
        RECT 86.100 17.200 86.400 17.600 ;
        RECT 86.650 17.200 86.950 17.600 ;
        RECT 87.200 17.500 87.500 17.600 ;
        RECT 88.450 17.500 88.850 17.600 ;
        RECT 89.200 17.500 89.500 17.600 ;
        RECT 87.200 17.300 88.250 17.500 ;
        RECT 87.200 17.200 87.500 17.300 ;
        RECT 81.150 16.600 81.800 16.650 ;
        RECT 79.450 16.400 81.800 16.600 ;
        RECT 82.500 16.450 83.000 16.850 ;
        RECT 83.500 16.600 83.900 17.000 ;
        RECT 79.450 16.200 79.850 16.400 ;
        RECT 81.150 16.250 81.800 16.400 ;
        RECT 81.600 16.000 81.800 16.250 ;
        RECT 82.800 16.000 83.000 16.450 ;
        RECT 83.700 16.400 83.900 16.600 ;
        RECT 85.000 16.400 85.200 17.200 ;
        RECT 85.500 17.000 85.900 17.200 ;
        RECT 86.150 17.000 86.350 17.200 ;
        RECT 87.250 17.000 87.450 17.200 ;
        RECT 85.500 16.800 87.450 17.000 ;
        RECT 83.700 16.200 85.200 16.400 ;
        RECT 85.650 16.500 86.050 16.550 ;
        RECT 87.450 16.500 87.850 16.550 ;
        RECT 85.650 16.300 87.850 16.500 ;
        RECT 85.650 16.200 86.050 16.300 ;
        RECT 87.450 16.200 87.850 16.300 ;
        RECT 83.900 16.000 84.100 16.200 ;
        RECT 85.000 16.000 85.200 16.200 ;
        RECT 88.050 16.000 88.250 17.300 ;
        RECT 88.450 17.300 89.500 17.500 ;
        RECT 88.450 17.200 88.850 17.300 ;
        RECT 89.200 17.200 89.500 17.300 ;
        RECT 89.750 17.200 90.450 17.600 ;
        RECT 90.750 17.200 91.200 17.600 ;
        RECT 91.450 17.200 91.750 17.600 ;
        RECT 92.000 17.200 92.300 17.600 ;
        RECT 92.700 17.200 93.000 17.600 ;
        RECT 93.250 17.200 93.550 17.600 ;
        RECT 93.800 17.200 94.100 17.600 ;
        RECT 95.700 17.500 96.000 17.600 ;
        RECT 95.150 17.300 96.000 17.500 ;
        RECT 79.750 15.900 80.050 16.000 ;
        RECT 78.950 15.700 80.050 15.900 ;
        RECT 79.750 15.600 80.050 15.700 ;
        RECT 80.300 15.600 80.600 16.000 ;
        RECT 81.550 15.600 81.850 16.000 ;
        RECT 82.100 15.600 82.400 16.000 ;
        RECT 82.800 15.600 83.100 16.000 ;
        RECT 83.350 15.600 83.650 16.000 ;
        RECT 83.900 15.600 84.200 16.000 ;
        RECT 84.450 15.600 84.750 16.000 ;
        RECT 85.000 15.600 85.300 16.000 ;
        RECT 85.700 15.600 86.400 16.000 ;
        RECT 86.650 15.600 86.950 16.000 ;
        RECT 87.200 15.600 87.500 16.000 ;
        RECT 87.750 15.700 88.250 16.000 ;
        RECT 88.650 16.000 88.850 17.200 ;
        RECT 89.100 16.400 89.500 16.550 ;
        RECT 90.750 16.400 90.950 17.200 ;
        RECT 92.050 17.000 92.250 17.200 ;
        RECT 91.150 16.800 92.250 17.000 ;
        RECT 91.150 16.600 91.750 16.800 ;
        RECT 89.100 16.200 91.300 16.400 ;
        RECT 90.000 16.000 90.200 16.200 ;
        RECT 91.100 16.000 91.300 16.200 ;
        RECT 91.550 16.000 91.750 16.600 ;
        RECT 92.000 16.400 92.400 16.600 ;
        RECT 92.750 16.400 92.950 17.200 ;
        RECT 93.850 16.400 94.050 17.200 ;
        RECT 95.150 16.700 95.350 17.300 ;
        RECT 95.700 17.200 96.000 17.300 ;
        RECT 96.250 17.200 96.950 17.600 ;
        RECT 97.250 17.200 97.700 17.600 ;
        RECT 97.950 17.200 98.250 17.600 ;
        RECT 98.500 17.200 98.800 17.600 ;
        RECT 99.200 17.200 99.500 17.600 ;
        RECT 99.750 17.200 100.050 17.600 ;
        RECT 100.300 17.200 100.600 17.600 ;
        RECT 102.200 17.500 102.500 17.600 ;
        RECT 101.650 17.300 102.500 17.500 ;
        RECT 92.000 16.200 94.050 16.400 ;
        RECT 94.350 16.500 95.350 16.700 ;
        RECT 94.350 16.300 94.750 16.500 ;
        RECT 93.850 16.000 94.050 16.200 ;
        RECT 88.650 15.700 89.150 16.000 ;
        RECT 87.750 15.600 88.050 15.700 ;
        RECT 88.850 15.600 89.150 15.700 ;
        RECT 89.400 15.600 89.700 16.000 ;
        RECT 89.950 15.600 90.250 16.000 ;
        RECT 90.500 15.600 90.800 16.000 ;
        RECT 91.050 15.600 91.350 16.000 ;
        RECT 91.550 15.800 92.450 16.000 ;
        RECT 92.150 15.600 92.450 15.800 ;
        RECT 92.700 15.600 93.000 16.000 ;
        RECT 93.250 15.600 93.600 16.000 ;
        RECT 93.800 15.600 94.100 16.000 ;
        RECT 61.600 15.400 61.800 15.600 ;
        RECT 61.500 15.000 61.900 15.400 ;
        RECT 62.600 14.850 62.800 15.600 ;
        RECT 63.700 14.850 63.900 15.600 ;
        RECT 66.050 14.850 66.250 15.600 ;
        RECT 66.450 15.100 66.850 15.500 ;
        RECT 67.200 15.400 67.400 15.600 ;
        RECT 67.100 15.050 67.500 15.400 ;
        RECT 67.750 14.850 67.950 15.600 ;
        RECT 68.850 14.850 69.050 15.600 ;
        RECT 71.050 14.850 71.250 15.600 ;
        RECT 71.800 15.050 72.200 15.400 ;
        RECT 73.350 15.150 73.650 15.550 ;
        RECT 73.400 14.850 73.600 15.150 ;
        RECT 74.650 14.850 74.850 15.600 ;
        RECT 75.750 14.850 75.950 15.600 ;
        RECT 78.100 14.850 78.300 15.600 ;
        RECT 79.800 15.050 80.200 15.400 ;
        RECT 80.400 14.850 80.600 15.600 ;
        RECT 82.150 14.850 82.350 15.600 ;
        RECT 83.400 14.850 83.600 15.600 ;
        RECT 84.500 14.850 84.700 15.600 ;
        RECT 86.150 14.850 86.350 15.600 ;
        RECT 89.450 14.850 89.650 15.600 ;
        RECT 90.550 14.850 90.750 15.600 ;
        RECT 92.870 15.000 93.200 15.400 ;
        RECT 93.400 14.850 93.600 15.600 ;
        RECT 95.150 15.550 95.350 16.500 ;
        RECT 95.600 15.950 96.000 16.150 ;
        RECT 97.250 15.950 97.450 17.200 ;
        RECT 98.550 17.000 98.750 17.200 ;
        RECT 97.650 16.800 98.750 17.000 ;
        RECT 97.650 16.600 98.250 16.800 ;
        RECT 95.600 15.750 97.800 15.950 ;
        RECT 96.500 15.550 96.700 15.750 ;
        RECT 97.600 15.550 97.800 15.750 ;
        RECT 98.050 15.550 98.250 16.600 ;
        RECT 98.500 15.950 98.900 16.150 ;
        RECT 99.250 15.950 99.450 17.200 ;
        RECT 100.350 15.950 100.550 17.200 ;
        RECT 101.650 16.700 101.850 17.300 ;
        RECT 102.200 17.200 102.500 17.300 ;
        RECT 102.750 17.200 103.450 17.600 ;
        RECT 103.750 17.200 104.200 17.600 ;
        RECT 104.450 17.200 104.750 17.600 ;
        RECT 105.000 17.200 105.300 17.600 ;
        RECT 105.700 17.200 106.000 17.600 ;
        RECT 106.250 17.200 106.550 17.600 ;
        RECT 106.800 17.200 107.100 17.600 ;
        RECT 108.700 17.500 109.000 17.600 ;
        RECT 108.150 17.300 109.000 17.500 ;
        RECT 100.850 16.500 101.850 16.700 ;
        RECT 100.850 16.300 101.250 16.500 ;
        RECT 98.500 15.750 100.550 15.950 ;
        RECT 100.350 15.550 100.550 15.750 ;
        RECT 101.650 15.550 101.850 16.500 ;
        RECT 102.100 15.950 102.500 16.150 ;
        RECT 103.750 15.950 103.950 17.200 ;
        RECT 105.050 17.000 105.250 17.200 ;
        RECT 104.150 16.800 105.250 17.000 ;
        RECT 104.150 16.600 104.750 16.800 ;
        RECT 102.100 15.750 104.300 15.950 ;
        RECT 103.000 15.550 103.200 15.750 ;
        RECT 104.100 15.550 104.300 15.750 ;
        RECT 104.550 15.550 104.750 16.600 ;
        RECT 105.000 15.950 105.400 16.150 ;
        RECT 105.750 15.950 105.950 17.200 ;
        RECT 106.850 15.950 107.050 17.200 ;
        RECT 108.150 16.700 108.350 17.300 ;
        RECT 108.700 17.200 109.000 17.300 ;
        RECT 109.250 17.200 109.950 17.600 ;
        RECT 110.250 17.200 110.700 17.600 ;
        RECT 110.950 17.200 111.250 17.600 ;
        RECT 111.500 17.200 111.800 17.600 ;
        RECT 112.200 17.200 112.500 17.600 ;
        RECT 112.750 17.200 113.050 17.600 ;
        RECT 113.300 17.200 113.600 17.600 ;
        RECT 107.350 16.500 108.350 16.700 ;
        RECT 107.350 16.300 107.750 16.500 ;
        RECT 105.000 15.750 107.050 15.950 ;
        RECT 106.850 15.550 107.050 15.750 ;
        RECT 108.150 15.550 108.350 16.500 ;
        RECT 108.600 15.950 109.000 16.150 ;
        RECT 110.250 15.950 110.450 17.200 ;
        RECT 111.550 17.000 111.750 17.200 ;
        RECT 110.650 16.800 111.750 17.000 ;
        RECT 110.650 16.600 111.250 16.800 ;
        RECT 108.600 15.750 110.800 15.950 ;
        RECT 109.500 15.550 109.700 15.750 ;
        RECT 110.600 15.550 110.800 15.750 ;
        RECT 111.050 15.550 111.250 16.600 ;
        RECT 111.500 15.950 111.900 16.150 ;
        RECT 112.250 15.950 112.450 17.200 ;
        RECT 113.350 15.950 113.550 17.200 ;
        RECT 115.450 17.100 115.650 27.450 ;
        RECT 117.900 27.350 118.300 27.450 ;
        RECT 120.500 27.350 120.900 27.450 ;
        RECT 123.100 27.350 123.500 27.450 ;
        RECT 125.700 27.350 126.100 27.450 ;
        RECT 116.050 25.200 116.350 27.100 ;
        RECT 117.950 25.200 118.250 27.100 ;
        RECT 118.650 25.200 118.950 27.100 ;
        RECT 120.550 25.200 120.850 27.100 ;
        RECT 121.250 25.200 121.550 27.100 ;
        RECT 123.150 25.200 123.450 27.100 ;
        RECT 123.850 25.200 124.150 27.100 ;
        RECT 125.750 25.200 126.050 27.100 ;
        RECT 116.950 24.600 117.350 25.000 ;
        RECT 119.550 24.600 119.950 25.000 ;
        RECT 122.150 24.600 122.550 25.000 ;
        RECT 124.800 24.600 125.100 25.000 ;
        RECT 116.050 20.750 116.350 23.650 ;
        RECT 116.600 20.750 116.900 23.650 ;
        RECT 118.650 20.750 118.950 23.650 ;
        RECT 119.200 20.750 119.500 23.650 ;
        RECT 121.250 20.750 121.550 23.650 ;
        RECT 121.800 20.750 122.100 23.650 ;
        RECT 116.400 20.200 116.690 20.550 ;
        RECT 119.000 20.200 119.290 20.550 ;
        RECT 121.600 20.200 121.890 20.550 ;
        RECT 116.040 17.850 116.340 19.750 ;
        RECT 116.600 17.850 116.900 19.750 ;
        RECT 118.640 17.850 118.940 19.750 ;
        RECT 119.200 17.850 119.500 19.750 ;
        RECT 121.240 17.850 121.540 19.750 ;
        RECT 121.800 17.850 122.100 19.750 ;
        RECT 116.260 17.300 116.550 17.650 ;
        RECT 118.860 17.300 119.150 17.650 ;
        RECT 121.460 17.300 121.750 17.650 ;
        RECT 126.400 17.100 126.600 27.450 ;
        RECT 115.450 16.900 126.600 17.100 ;
        RECT 113.760 16.300 114.050 16.700 ;
        RECT 111.500 15.750 113.550 15.950 ;
        RECT 113.350 15.550 113.550 15.750 ;
        RECT 115.450 15.900 125.650 16.100 ;
        RECT 94.650 15.150 94.950 15.550 ;
        RECT 95.150 15.250 95.650 15.550 ;
        RECT 95.350 15.150 95.650 15.250 ;
        RECT 95.900 15.150 96.200 15.550 ;
        RECT 96.450 15.150 96.750 15.550 ;
        RECT 97.000 15.150 97.300 15.550 ;
        RECT 97.550 15.150 97.850 15.550 ;
        RECT 98.050 15.350 98.950 15.550 ;
        RECT 98.650 15.150 98.950 15.350 ;
        RECT 99.200 15.150 99.500 15.550 ;
        RECT 99.750 15.150 100.050 15.550 ;
        RECT 100.300 15.150 100.600 15.550 ;
        RECT 101.150 15.150 101.450 15.550 ;
        RECT 101.650 15.250 102.150 15.550 ;
        RECT 101.850 15.150 102.150 15.250 ;
        RECT 102.400 15.150 102.700 15.550 ;
        RECT 102.950 15.150 103.250 15.550 ;
        RECT 103.500 15.150 103.800 15.550 ;
        RECT 104.050 15.150 104.350 15.550 ;
        RECT 104.550 15.350 105.450 15.550 ;
        RECT 105.150 15.150 105.450 15.350 ;
        RECT 105.700 15.150 106.000 15.550 ;
        RECT 106.250 15.150 106.550 15.550 ;
        RECT 106.800 15.150 107.100 15.550 ;
        RECT 107.650 15.150 107.950 15.550 ;
        RECT 108.150 15.250 108.650 15.550 ;
        RECT 108.350 15.150 108.650 15.250 ;
        RECT 108.900 15.150 109.200 15.550 ;
        RECT 109.450 15.150 109.750 15.550 ;
        RECT 110.000 15.150 110.300 15.550 ;
        RECT 110.550 15.150 110.850 15.550 ;
        RECT 111.050 15.350 111.950 15.550 ;
        RECT 111.650 15.150 111.950 15.350 ;
        RECT 112.200 15.150 112.500 15.550 ;
        RECT 112.750 15.150 113.050 15.550 ;
        RECT 113.300 15.150 113.600 15.550 ;
        RECT 94.700 14.850 94.900 15.150 ;
        RECT 95.950 14.850 96.150 15.150 ;
        RECT 97.050 14.850 97.250 15.150 ;
        RECT 99.800 14.850 100.000 15.150 ;
        RECT 101.200 14.850 101.400 15.150 ;
        RECT 102.450 14.850 102.650 15.150 ;
        RECT 103.550 14.850 103.750 15.150 ;
        RECT 106.300 14.850 106.500 15.150 ;
        RECT 107.700 14.850 107.900 15.150 ;
        RECT 108.950 14.850 109.150 15.150 ;
        RECT 110.050 14.850 110.250 15.150 ;
        RECT 112.800 14.850 113.000 15.150 ;
        RECT 62.500 14.450 62.900 14.850 ;
        RECT 63.600 14.450 64.000 14.850 ;
        RECT 65.950 14.450 66.350 14.850 ;
        RECT 67.650 14.450 68.050 14.850 ;
        RECT 68.750 14.450 69.150 14.850 ;
        RECT 70.950 14.450 71.350 14.850 ;
        RECT 73.300 14.450 73.700 14.850 ;
        RECT 74.550 14.450 74.950 14.850 ;
        RECT 75.650 14.450 76.050 14.850 ;
        RECT 78.000 14.450 78.400 14.850 ;
        RECT 80.300 14.450 80.700 14.850 ;
        RECT 82.050 14.450 82.450 14.850 ;
        RECT 83.300 14.450 83.700 14.850 ;
        RECT 84.400 14.450 84.800 14.850 ;
        RECT 86.050 14.450 86.450 14.850 ;
        RECT 89.350 14.450 89.750 14.850 ;
        RECT 90.450 14.450 90.850 14.850 ;
        RECT 93.300 14.450 93.700 14.850 ;
        RECT 94.600 14.450 95.000 14.850 ;
        RECT 95.850 14.450 96.250 14.850 ;
        RECT 96.950 14.450 97.350 14.850 ;
        RECT 99.700 14.450 100.100 14.850 ;
        RECT 101.100 14.450 101.500 14.850 ;
        RECT 102.350 14.450 102.750 14.850 ;
        RECT 103.450 14.450 103.850 14.850 ;
        RECT 106.200 14.450 106.600 14.850 ;
        RECT 107.600 14.450 108.000 14.850 ;
        RECT 108.850 14.450 109.250 14.850 ;
        RECT 109.950 14.450 110.350 14.850 ;
        RECT 112.700 14.450 113.100 14.850 ;
        RECT 115.450 9.600 115.650 15.900 ;
        RECT 116.260 15.350 116.550 15.700 ;
        RECT 118.860 15.350 119.150 15.700 ;
        RECT 121.460 15.350 121.750 15.700 ;
        RECT 116.040 14.250 116.340 15.150 ;
        RECT 116.600 14.250 116.900 15.150 ;
        RECT 118.640 14.250 118.940 15.150 ;
        RECT 119.200 14.250 119.500 15.150 ;
        RECT 121.240 14.250 121.540 15.150 ;
        RECT 121.800 14.250 122.100 15.150 ;
        RECT 116.400 13.450 116.690 13.800 ;
        RECT 119.000 13.450 119.290 13.800 ;
        RECT 121.600 13.450 121.890 13.800 ;
        RECT 116.050 11.850 116.350 13.250 ;
        RECT 116.600 11.850 116.900 13.250 ;
        RECT 118.650 11.850 118.950 13.250 ;
        RECT 119.200 11.850 119.500 13.250 ;
        RECT 121.250 11.850 121.550 13.250 ;
        RECT 121.800 11.850 122.100 13.250 ;
        RECT 116.330 11.050 116.620 11.400 ;
        RECT 118.930 11.050 119.220 11.400 ;
        RECT 121.530 11.050 121.820 11.400 ;
        RECT 124.370 11.050 124.660 11.400 ;
        RECT 116.050 9.950 116.350 10.850 ;
        RECT 116.600 9.950 116.900 10.850 ;
        RECT 118.650 9.950 118.950 10.850 ;
        RECT 119.200 9.950 119.500 10.850 ;
        RECT 121.250 9.950 121.550 10.850 ;
        RECT 121.800 9.950 122.100 10.850 ;
        RECT 124.250 9.950 124.550 10.850 ;
        RECT 124.800 9.950 125.100 10.850 ;
        RECT 116.550 9.600 116.950 9.700 ;
        RECT 119.150 9.600 119.550 9.700 ;
        RECT 121.750 9.600 122.150 9.700 ;
        RECT 124.200 9.600 124.600 9.700 ;
        RECT 125.450 9.600 125.650 15.900 ;
        RECT 115.450 9.400 125.650 9.600 ;
        RECT 116.550 9.300 116.950 9.400 ;
        RECT 119.150 9.300 119.550 9.400 ;
        RECT 121.750 9.300 122.150 9.400 ;
        RECT 124.200 9.300 124.600 9.400 ;
      LAYER met1 ;
        RECT 80.600 100.100 81.000 100.500 ;
        RECT 129.950 99.550 130.450 99.600 ;
        RECT 74.950 99.150 77.100 99.550 ;
        RECT 84.500 99.150 86.650 99.550 ;
        RECT 129.950 99.100 132.400 99.550 ;
        RECT 43.950 94.650 44.350 97.450 ;
        RECT 43.850 92.115 44.440 94.220 ;
        RECT 45.850 92.150 46.250 98.000 ;
        RECT 47.850 92.100 48.250 97.450 ;
        RECT 53.400 92.150 53.800 97.450 ;
        RECT 43.850 85.190 44.440 87.295 ;
        RECT 43.950 48.450 44.350 85.190 ;
        RECT 47.300 55.100 47.700 71.100 ;
        RECT 47.850 55.650 48.250 79.500 ;
        RECT 51.750 75.250 52.150 85.600 ;
        RECT 48.400 46.200 48.800 72.500 ;
        RECT 53.100 60.250 53.500 71.950 ;
        RECT 55.150 71.550 55.550 98.000 ;
        RECT 66.200 96.250 66.600 97.450 ;
        RECT 57.850 90.950 74.950 94.450 ;
        RECT 78.350 92.150 78.750 97.450 ;
        RECT 83.900 92.150 84.300 97.450 ;
        RECT 87.850 94.650 88.250 97.450 ;
        RECT 90.950 95.900 91.350 98.000 ;
        RECT 83.970 92.145 84.220 92.150 ;
        RECT 87.750 92.115 88.340 94.220 ;
        RECT 55.700 73.700 56.100 86.100 ;
        RECT 57.850 80.850 61.350 90.950 ;
        RECT 64.650 84.150 68.150 87.650 ;
        RECT 71.450 80.850 74.950 90.950 ;
        RECT 57.850 77.350 74.950 80.850 ;
        RECT 76.700 75.650 77.100 86.100 ;
        RECT 80.000 75.650 80.400 85.600 ;
        RECT 87.750 85.190 88.340 87.295 ;
        RECT 81.200 75.650 81.600 76.050 ;
        RECT 57.700 73.700 59.900 74.100 ;
        RECT 72.900 73.700 75.100 75.650 ;
        RECT 80.750 73.700 81.150 74.100 ;
        RECT 75.500 73.150 75.900 73.550 ;
        RECT 55.400 70.700 55.800 71.100 ;
        RECT 77.350 70.500 77.750 71.300 ;
        RECT 78.550 70.500 78.950 73.550 ;
        RECT 55.800 69.850 56.200 70.250 ;
        RECT 56.600 69.850 57.000 70.250 ;
        RECT 57.400 69.850 57.800 70.250 ;
        RECT 58.200 69.850 58.600 70.250 ;
        RECT 59.000 69.850 59.400 70.250 ;
        RECT 59.800 69.850 60.200 70.250 ;
        RECT 60.600 69.850 61.000 70.250 ;
        RECT 61.400 69.850 61.800 70.250 ;
        RECT 62.200 69.850 62.600 70.250 ;
        RECT 63.000 69.850 63.400 70.250 ;
        RECT 63.800 69.850 64.200 70.250 ;
        RECT 64.600 69.850 65.000 70.250 ;
        RECT 65.400 69.850 65.800 70.250 ;
        RECT 66.200 69.850 66.600 70.250 ;
        RECT 67.000 69.850 67.400 70.250 ;
        RECT 67.800 69.850 68.200 70.250 ;
        RECT 68.600 69.850 69.000 70.250 ;
        RECT 69.400 69.850 69.800 70.250 ;
        RECT 70.200 69.850 70.600 70.250 ;
        RECT 71.000 69.850 71.400 70.250 ;
        RECT 71.800 69.850 72.200 70.250 ;
        RECT 72.600 69.850 73.000 70.250 ;
        RECT 73.400 69.850 73.800 70.250 ;
        RECT 74.200 69.850 74.600 70.250 ;
        RECT 75.000 69.850 75.400 70.250 ;
        RECT 75.800 69.850 76.200 70.250 ;
        RECT 59.500 68.500 59.900 69.700 ;
        RECT 53.700 63.950 54.100 65.900 ;
        RECT 54.600 64.500 55.000 65.700 ;
        RECT 55.800 64.500 56.200 65.700 ;
        RECT 57.000 64.500 57.400 65.700 ;
        RECT 58.200 64.500 58.600 65.700 ;
        RECT 61.400 64.500 61.800 65.700 ;
        RECT 62.600 64.500 63.000 65.700 ;
        RECT 63.800 64.500 64.200 65.700 ;
        RECT 57.450 63.950 57.850 64.350 ;
        RECT 58.550 63.950 58.950 64.350 ;
        RECT 59.850 63.950 60.250 64.350 ;
        RECT 60.950 63.950 61.350 64.350 ;
        RECT 62.250 63.950 62.650 64.350 ;
        RECT 57.155 63.450 57.445 63.800 ;
        RECT 57.600 63.250 57.750 63.950 ;
        RECT 58.650 63.250 58.800 63.950 ;
        RECT 58.955 63.450 59.245 63.800 ;
        RECT 59.555 63.450 59.845 63.800 ;
        RECT 60.000 63.250 60.150 63.950 ;
        RECT 61.050 63.250 61.200 63.950 ;
        RECT 61.355 63.450 61.645 63.800 ;
        RECT 61.955 63.450 62.245 63.800 ;
        RECT 62.400 63.250 62.550 63.950 ;
        RECT 56.850 61.600 57.150 63.250 ;
        RECT 57.450 62.850 57.750 63.250 ;
        RECT 58.050 62.850 58.350 63.250 ;
        RECT 58.650 62.850 58.950 63.250 ;
        RECT 59.250 62.850 59.550 63.250 ;
        RECT 59.850 62.850 60.150 63.250 ;
        RECT 60.450 62.850 60.750 63.250 ;
        RECT 61.050 62.850 61.350 63.250 ;
        RECT 61.650 62.850 61.950 63.250 ;
        RECT 62.250 62.850 62.550 63.250 ;
        RECT 62.850 62.850 63.150 63.250 ;
        RECT 57.660 62.300 57.950 62.650 ;
        RECT 58.100 62.150 58.300 62.850 ;
        RECT 58.450 62.300 58.740 62.650 ;
        RECT 53.100 59.850 53.900 60.250 ;
        RECT 55.600 59.850 56.000 60.250 ;
        RECT 56.800 59.850 57.200 61.600 ;
        RECT 53.550 59.300 53.850 59.850 ;
        RECT 54.400 59.250 54.800 59.650 ;
        RECT 52.650 57.400 52.950 59.050 ;
        RECT 53.250 57.950 53.550 59.050 ;
        RECT 53.200 57.550 53.600 57.950 ;
        RECT 53.850 57.400 54.150 59.050 ;
        RECT 54.450 58.150 54.750 59.250 ;
        RECT 55.050 57.400 55.350 59.050 ;
        RECT 55.650 58.150 55.950 59.850 ;
        RECT 56.850 59.250 57.150 59.850 ;
        RECT 58.000 59.250 58.400 62.150 ;
        RECT 59.300 61.600 59.500 62.850 ;
        RECT 60.070 62.300 60.360 62.650 ;
        RECT 60.500 62.150 60.700 62.850 ;
        RECT 60.840 62.300 61.130 62.650 ;
        RECT 60.400 61.750 60.800 62.150 ;
        RECT 61.700 61.600 61.900 62.850 ;
        RECT 62.460 62.300 62.750 62.650 ;
        RECT 62.900 62.150 63.100 62.850 ;
        RECT 64.000 62.500 64.400 63.700 ;
        RECT 62.800 61.750 63.200 62.150 ;
        RECT 59.200 61.200 59.600 61.600 ;
        RECT 61.600 61.200 62.000 61.600 ;
        RECT 59.200 59.850 59.600 60.250 ;
        RECT 60.400 59.850 60.800 60.250 ;
        RECT 62.800 59.850 63.200 60.250 ;
        RECT 63.700 59.850 64.100 60.250 ;
        RECT 56.250 57.400 56.550 59.050 ;
        RECT 56.850 57.950 57.150 59.050 ;
        RECT 56.800 57.550 57.200 57.950 ;
        RECT 57.450 57.400 57.750 59.050 ;
        RECT 58.050 58.150 58.350 59.250 ;
        RECT 58.650 57.400 58.950 59.050 ;
        RECT 59.250 58.150 59.550 59.850 ;
        RECT 60.450 59.250 60.750 59.850 ;
        RECT 61.600 59.250 62.000 59.650 ;
        RECT 59.850 57.400 60.150 59.050 ;
        RECT 60.450 57.950 60.750 59.050 ;
        RECT 60.400 57.550 60.800 57.950 ;
        RECT 61.050 57.400 61.350 59.050 ;
        RECT 61.650 58.150 61.950 59.250 ;
        RECT 62.250 57.400 62.550 59.050 ;
        RECT 62.850 58.150 63.150 59.850 ;
        RECT 63.750 59.250 64.050 59.850 ;
        RECT 63.450 57.400 63.750 59.050 ;
        RECT 64.050 57.950 64.350 59.050 ;
        RECT 64.000 57.550 64.400 57.950 ;
        RECT 64.650 57.400 64.950 59.050 ;
        RECT 65.350 57.950 65.650 65.850 ;
        RECT 65.800 62.500 67.000 69.700 ;
        RECT 72.900 68.500 73.300 69.700 ;
        RECT 67.150 57.950 67.450 65.850 ;
        RECT 68.600 64.500 69.000 65.700 ;
        RECT 69.800 64.500 70.200 65.700 ;
        RECT 71.000 64.500 71.400 65.700 ;
        RECT 74.200 64.500 74.600 65.700 ;
        RECT 75.400 64.500 75.800 65.700 ;
        RECT 76.600 64.500 77.000 65.700 ;
        RECT 77.800 64.500 78.200 65.700 ;
        RECT 78.750 64.350 79.050 68.300 ;
        RECT 70.150 63.950 70.550 64.350 ;
        RECT 71.450 63.950 71.850 64.350 ;
        RECT 72.550 63.950 72.950 64.350 ;
        RECT 73.850 63.950 74.250 64.350 ;
        RECT 74.950 63.950 75.350 64.350 ;
        RECT 78.700 63.950 79.100 64.350 ;
        RECT 68.400 62.500 68.800 63.700 ;
        RECT 70.250 63.250 70.400 63.950 ;
        RECT 70.555 63.450 70.845 63.800 ;
        RECT 71.155 63.450 71.445 63.800 ;
        RECT 71.600 63.250 71.750 63.950 ;
        RECT 72.650 63.250 72.800 63.950 ;
        RECT 72.955 63.450 73.245 63.800 ;
        RECT 73.555 63.450 73.845 63.800 ;
        RECT 74.000 63.250 74.150 63.950 ;
        RECT 75.050 63.250 75.200 63.950 ;
        RECT 80.850 63.800 81.050 73.700 ;
        RECT 75.355 63.450 75.645 63.800 ;
        RECT 80.750 63.400 81.150 63.800 ;
        RECT 69.650 62.850 69.950 63.250 ;
        RECT 70.250 62.850 70.550 63.250 ;
        RECT 70.850 62.850 71.150 63.250 ;
        RECT 71.450 62.850 71.750 63.250 ;
        RECT 72.050 62.850 72.350 63.250 ;
        RECT 72.650 62.850 72.950 63.250 ;
        RECT 73.250 62.850 73.550 63.250 ;
        RECT 73.850 62.850 74.150 63.250 ;
        RECT 74.450 62.850 74.750 63.250 ;
        RECT 75.050 62.850 75.350 63.250 ;
        RECT 69.700 62.150 69.900 62.850 ;
        RECT 70.050 62.300 70.340 62.650 ;
        RECT 69.600 61.750 70.000 62.150 ;
        RECT 70.900 61.600 71.100 62.850 ;
        RECT 71.670 62.300 71.960 62.650 ;
        RECT 72.100 62.150 72.300 62.850 ;
        RECT 72.440 62.300 72.730 62.650 ;
        RECT 72.000 61.750 72.400 62.150 ;
        RECT 73.300 61.600 73.500 62.850 ;
        RECT 74.060 62.300 74.350 62.650 ;
        RECT 74.500 62.150 74.700 62.850 ;
        RECT 74.850 62.300 75.140 62.650 ;
        RECT 70.800 61.200 71.200 61.600 ;
        RECT 73.200 61.200 73.600 61.600 ;
        RECT 68.700 59.850 69.100 61.050 ;
        RECT 69.600 59.850 70.000 61.050 ;
        RECT 70.800 59.850 71.200 61.050 ;
        RECT 72.000 59.850 72.400 61.050 ;
        RECT 73.200 59.850 73.600 61.050 ;
        RECT 68.750 59.250 69.050 59.850 ;
        RECT 65.300 57.550 65.700 57.950 ;
        RECT 52.600 56.200 53.000 57.400 ;
        RECT 53.800 56.200 54.200 57.400 ;
        RECT 55.000 56.200 55.400 57.400 ;
        RECT 56.200 56.200 56.600 57.400 ;
        RECT 57.400 56.200 57.800 57.400 ;
        RECT 58.600 56.200 59.000 57.400 ;
        RECT 59.800 56.200 60.200 57.400 ;
        RECT 61.000 56.200 61.400 57.400 ;
        RECT 62.200 56.200 62.600 57.400 ;
        RECT 63.400 56.200 63.800 57.400 ;
        RECT 64.600 56.200 65.000 57.400 ;
        RECT 59.000 55.650 59.400 56.050 ;
        RECT 66.200 55.650 66.600 56.050 ;
        RECT 58.150 50.350 58.450 53.250 ;
        RECT 59.050 50.350 59.350 55.650 ;
        RECT 60.800 55.100 61.200 55.500 ;
        RECT 59.500 53.450 59.850 53.850 ;
        RECT 60.350 53.450 60.750 53.850 ;
        RECT 60.900 53.250 61.100 55.100 ;
        RECT 62.600 54.550 63.000 54.950 ;
        RECT 61.250 53.450 61.650 53.850 ;
        RECT 62.150 53.450 62.550 53.850 ;
        RECT 62.700 53.250 62.900 54.550 ;
        RECT 64.400 54.000 64.800 54.400 ;
        RECT 63.050 53.450 63.450 53.850 ;
        RECT 63.950 53.450 64.350 53.850 ;
        RECT 64.500 53.250 64.700 54.000 ;
        RECT 64.850 53.450 65.250 53.850 ;
        RECT 65.750 53.450 66.100 53.850 ;
        RECT 59.950 50.350 60.250 53.250 ;
        RECT 60.850 50.350 61.150 53.250 ;
        RECT 61.750 50.350 62.050 53.250 ;
        RECT 62.650 50.350 62.950 53.250 ;
        RECT 63.550 50.350 63.850 53.250 ;
        RECT 64.450 50.350 64.750 53.250 ;
        RECT 65.350 50.350 65.650 53.250 ;
        RECT 66.250 50.350 66.550 55.650 ;
        RECT 67.100 53.850 67.500 57.950 ;
        RECT 67.850 57.400 68.150 59.050 ;
        RECT 68.450 57.950 68.750 59.050 ;
        RECT 68.400 57.550 68.800 57.950 ;
        RECT 69.050 57.400 69.350 59.050 ;
        RECT 69.650 58.150 69.950 59.850 ;
        RECT 70.800 59.250 71.200 59.650 ;
        RECT 72.050 59.250 72.350 59.850 ;
        RECT 70.250 57.400 70.550 59.050 ;
        RECT 70.850 58.150 71.150 59.250 ;
        RECT 71.450 57.400 71.750 59.050 ;
        RECT 72.050 57.950 72.350 59.050 ;
        RECT 72.000 57.550 72.400 57.950 ;
        RECT 72.650 57.400 72.950 59.050 ;
        RECT 73.250 58.150 73.550 59.850 ;
        RECT 74.400 59.250 74.800 62.150 ;
        RECT 75.650 61.600 75.950 63.250 ;
        RECT 75.600 59.850 76.000 61.600 ;
        RECT 76.800 59.850 77.200 61.050 ;
        RECT 78.900 59.850 79.300 61.050 ;
        RECT 75.650 59.250 75.950 59.850 ;
        RECT 73.850 57.400 74.150 59.050 ;
        RECT 74.450 58.150 74.750 59.250 ;
        RECT 75.050 57.400 75.350 59.050 ;
        RECT 75.650 57.950 75.950 59.050 ;
        RECT 75.600 57.550 76.000 57.950 ;
        RECT 76.250 57.400 76.550 59.050 ;
        RECT 76.850 58.150 77.150 59.850 ;
        RECT 78.000 59.250 78.400 59.650 ;
        RECT 78.950 59.300 79.250 59.850 ;
        RECT 77.450 57.400 77.750 59.050 ;
        RECT 78.050 58.150 78.350 59.250 ;
        RECT 78.650 57.400 78.950 59.050 ;
        RECT 79.250 57.950 79.550 59.050 ;
        RECT 67.800 56.200 68.200 57.400 ;
        RECT 69.000 56.200 69.400 57.400 ;
        RECT 70.200 56.200 70.600 57.400 ;
        RECT 71.400 56.200 71.800 57.400 ;
        RECT 72.600 56.200 73.000 57.400 ;
        RECT 73.800 56.200 74.200 57.400 ;
        RECT 75.000 56.200 75.400 57.400 ;
        RECT 76.200 56.200 76.600 57.400 ;
        RECT 77.400 56.200 77.800 57.400 ;
        RECT 78.600 56.200 79.000 57.400 ;
        RECT 73.400 55.650 73.800 56.050 ;
        RECT 71.600 55.100 72.000 55.500 ;
        RECT 69.800 54.550 70.200 54.950 ;
        RECT 68.000 54.000 68.400 54.400 ;
        RECT 66.700 53.450 67.950 53.850 ;
        RECT 68.100 53.250 68.300 54.000 ;
        RECT 68.450 53.450 68.850 53.850 ;
        RECT 69.350 53.450 69.750 53.850 ;
        RECT 69.900 53.250 70.100 54.550 ;
        RECT 70.250 53.450 70.650 53.850 ;
        RECT 71.150 53.450 71.550 53.850 ;
        RECT 71.700 53.250 71.900 55.100 ;
        RECT 72.050 53.450 72.450 53.850 ;
        RECT 72.950 53.450 73.300 53.850 ;
        RECT 67.150 50.350 67.450 53.250 ;
        RECT 68.050 50.350 68.350 53.250 ;
        RECT 68.950 50.350 69.250 53.250 ;
        RECT 69.850 50.350 70.150 53.250 ;
        RECT 70.750 50.350 71.050 53.250 ;
        RECT 71.650 50.350 71.950 53.250 ;
        RECT 72.550 50.350 72.850 53.250 ;
        RECT 73.450 50.350 73.750 55.650 ;
        RECT 76.200 54.550 76.600 54.950 ;
        RECT 74.350 50.350 74.650 53.250 ;
        RECT 76.300 51.150 76.500 54.550 ;
        RECT 77.950 52.450 78.350 52.850 ;
        RECT 78.550 52.450 78.950 55.500 ;
        RECT 79.200 52.850 79.600 57.950 ;
        RECT 79.850 57.400 80.150 59.050 ;
        RECT 79.800 56.200 80.200 57.400 ;
        RECT 80.850 54.400 81.050 63.400 ;
        RECT 81.300 62.650 81.500 75.650 ;
        RECT 81.200 62.250 81.600 62.650 ;
        RECT 81.300 54.950 81.500 62.250 ;
        RECT 81.750 59.850 82.950 78.850 ;
        RECT 83.900 72.100 84.300 83.950 ;
        RECT 87.850 57.550 88.250 85.190 ;
        RECT 89.750 81.900 90.150 94.300 ;
        RECT 93.200 92.350 93.700 92.850 ;
        RECT 90.600 67.200 91.000 89.300 ;
        RECT 93.250 71.550 93.650 92.350 ;
        RECT 93.900 85.350 94.400 85.850 ;
        RECT 93.900 78.350 94.400 78.850 ;
        RECT 116.170 69.650 116.420 70.050 ;
        RECT 116.050 69.150 116.550 69.650 ;
        RECT 115.050 67.550 115.450 67.950 ;
        RECT 116.170 67.945 116.420 69.150 ;
        RECT 90.200 66.700 91.400 67.200 ;
        RECT 81.200 54.550 81.600 54.950 ;
        RECT 80.750 54.000 81.150 54.400 ;
        RECT 79.150 52.450 79.550 52.850 ;
        RECT 77.500 51.150 77.800 52.250 ;
        RECT 78.050 51.350 78.350 52.450 ;
        RECT 78.600 51.150 78.900 52.250 ;
        RECT 79.150 51.350 79.450 52.450 ;
        RECT 79.700 51.150 80.000 52.250 ;
        RECT 76.200 50.750 76.600 51.150 ;
        RECT 77.450 50.750 77.850 51.150 ;
        RECT 78.550 50.750 78.950 51.150 ;
        RECT 79.650 50.750 80.050 51.150 ;
        RECT 77.500 50.150 77.800 50.750 ;
        RECT 79.700 50.150 80.000 50.750 ;
        RECT 58.100 48.950 58.500 50.150 ;
        RECT 59.900 48.950 60.300 50.150 ;
        RECT 61.700 48.950 62.100 50.150 ;
        RECT 63.500 48.950 63.900 50.150 ;
        RECT 65.300 48.950 65.700 50.150 ;
        RECT 67.100 48.950 67.500 50.150 ;
        RECT 68.900 48.950 69.300 50.150 ;
        RECT 70.700 48.950 71.100 50.150 ;
        RECT 72.500 48.950 72.900 50.150 ;
        RECT 74.300 48.950 74.700 50.150 ;
        RECT 77.450 48.950 77.850 50.150 ;
        RECT 79.650 48.950 80.050 50.150 ;
        RECT 59.030 48.450 59.320 48.800 ;
        RECT 59.580 48.450 59.870 48.800 ;
        RECT 60.130 48.450 60.420 48.800 ;
        RECT 60.680 48.450 60.970 48.800 ;
        RECT 61.230 48.450 61.520 48.800 ;
        RECT 61.780 48.450 62.070 48.800 ;
        RECT 62.330 48.450 62.620 48.800 ;
        RECT 62.880 48.450 63.170 48.800 ;
        RECT 63.430 48.450 63.720 48.800 ;
        RECT 63.980 48.450 64.270 48.800 ;
        RECT 68.530 48.450 68.820 48.800 ;
        RECT 69.080 48.450 69.370 48.800 ;
        RECT 69.630 48.450 69.920 48.800 ;
        RECT 70.180 48.450 70.470 48.800 ;
        RECT 70.730 48.450 71.020 48.800 ;
        RECT 71.280 48.450 71.570 48.800 ;
        RECT 71.830 48.450 72.120 48.800 ;
        RECT 72.380 48.450 72.670 48.800 ;
        RECT 72.930 48.450 73.220 48.800 ;
        RECT 73.480 48.450 73.770 48.800 ;
        RECT 57.800 47.350 58.500 48.250 ;
        RECT 58.200 47.150 58.500 47.350 ;
        RECT 58.150 46.750 58.550 47.150 ;
        RECT 58.750 46.600 59.050 48.250 ;
        RECT 59.300 47.150 59.600 48.250 ;
        RECT 59.250 46.750 59.650 47.150 ;
        RECT 59.850 46.600 60.150 48.250 ;
        RECT 60.400 47.150 60.700 48.250 ;
        RECT 60.350 46.750 60.750 47.150 ;
        RECT 60.950 46.600 61.250 48.250 ;
        RECT 61.500 47.150 61.800 48.250 ;
        RECT 61.450 46.750 61.850 47.150 ;
        RECT 62.050 46.600 62.350 48.250 ;
        RECT 62.600 47.150 62.900 48.250 ;
        RECT 62.550 46.750 62.950 47.150 ;
        RECT 63.150 46.600 63.450 48.250 ;
        RECT 63.700 47.150 64.000 48.250 ;
        RECT 63.650 46.750 64.050 47.150 ;
        RECT 64.250 46.600 64.550 48.250 ;
        RECT 64.800 47.350 65.500 48.250 ;
        RECT 67.300 47.350 68.000 48.250 ;
        RECT 64.800 47.150 65.100 47.350 ;
        RECT 67.700 47.150 68.000 47.350 ;
        RECT 64.750 46.750 65.150 47.150 ;
        RECT 67.650 46.750 68.050 47.150 ;
        RECT 58.700 46.200 59.100 46.600 ;
        RECT 59.800 46.200 60.200 46.600 ;
        RECT 60.900 46.200 61.300 46.600 ;
        RECT 62.000 46.200 62.400 46.600 ;
        RECT 63.100 46.200 63.500 46.600 ;
        RECT 64.200 46.200 64.600 46.600 ;
        RECT 68.250 46.550 68.550 48.250 ;
        RECT 68.800 47.150 69.100 48.250 ;
        RECT 68.750 46.750 69.150 47.150 ;
        RECT 69.350 46.550 69.650 48.250 ;
        RECT 69.900 47.150 70.200 48.250 ;
        RECT 69.850 46.750 70.250 47.150 ;
        RECT 70.450 46.550 70.750 48.250 ;
        RECT 71.000 47.150 71.300 48.250 ;
        RECT 70.950 46.750 71.350 47.150 ;
        RECT 71.550 46.550 71.850 48.250 ;
        RECT 72.100 47.150 72.400 48.250 ;
        RECT 72.050 46.750 72.450 47.150 ;
        RECT 72.650 46.550 72.950 48.250 ;
        RECT 73.200 47.150 73.500 48.250 ;
        RECT 73.150 46.750 73.550 47.150 ;
        RECT 73.750 46.550 74.050 48.250 ;
        RECT 74.300 47.350 75.000 48.250 ;
        RECT 74.300 47.150 74.600 47.350 ;
        RECT 74.250 46.750 74.650 47.150 ;
        RECT 68.200 45.350 68.600 46.550 ;
        RECT 69.300 45.350 69.700 46.550 ;
        RECT 70.400 45.350 70.800 46.550 ;
        RECT 71.500 45.350 71.900 46.550 ;
        RECT 72.600 45.350 73.000 46.550 ;
        RECT 73.700 45.350 74.100 46.550 ;
        RECT 66.250 41.150 66.650 41.550 ;
        RECT 67.350 41.150 67.750 41.550 ;
        RECT 68.850 41.150 69.250 41.550 ;
        RECT 70.000 41.150 70.400 41.550 ;
        RECT 70.750 41.150 71.150 41.550 ;
        RECT 71.850 41.150 72.250 41.550 ;
        RECT 73.350 41.150 73.750 41.550 ;
        RECT 74.450 41.150 74.850 41.550 ;
        RECT 76.450 41.150 76.850 41.550 ;
        RECT 78.100 41.150 78.500 41.550 ;
        RECT 79.750 41.150 80.150 41.550 ;
        RECT 81.950 41.150 82.350 41.550 ;
        RECT 83.250 41.150 83.650 41.550 ;
        RECT 85.850 41.150 86.250 41.550 ;
        RECT 89.250 41.150 89.650 41.550 ;
        RECT 59.700 6.300 60.100 32.200 ;
        RECT 60.250 16.350 60.650 39.100 ;
        RECT 65.650 38.700 66.050 39.100 ;
        RECT 75.250 38.650 75.650 39.050 ;
        RECT 80.400 38.650 81.000 39.050 ;
        RECT 68.500 35.800 68.900 36.200 ;
        RECT 66.250 35.250 66.650 35.650 ;
        RECT 69.950 35.250 70.350 35.650 ;
        RECT 70.750 35.250 71.150 35.650 ;
        RECT 74.450 35.250 74.850 35.650 ;
        RECT 65.650 31.800 66.050 32.200 ;
        RECT 75.350 32.050 75.550 38.650 ;
        RECT 76.150 35.800 76.550 36.200 ;
        RECT 75.700 35.250 76.100 35.650 ;
        RECT 76.250 35.050 76.450 35.800 ;
        RECT 76.650 35.250 77.450 35.650 ;
        RECT 78.100 35.250 78.500 35.650 ;
        RECT 79.750 35.250 80.150 35.650 ;
        RECT 76.250 34.700 76.650 35.050 ;
        RECT 80.800 32.250 81.000 38.650 ;
        RECT 81.150 38.700 81.550 39.100 ;
        RECT 81.150 36.250 81.350 38.700 ;
        RECT 81.150 35.850 81.550 36.250 ;
        RECT 83.350 36.150 83.550 41.150 ;
        RECT 84.500 40.600 85.250 41.000 ;
        RECT 87.650 40.600 88.050 41.000 ;
        RECT 90.500 40.600 90.900 41.900 ;
        RECT 83.250 35.850 83.650 36.150 ;
        RECT 84.100 35.850 84.500 36.200 ;
        RECT 85.050 35.650 85.250 40.600 ;
        RECT 90.000 38.900 90.400 39.300 ;
        RECT 90.900 37.100 91.300 39.300 ;
        RECT 87.300 35.800 87.700 36.200 ;
        RECT 90.900 35.800 91.300 36.950 ;
        RECT 93.250 36.550 94.450 46.550 ;
        RECT 81.950 35.250 82.350 35.650 ;
        RECT 83.900 35.250 84.300 35.650 ;
        RECT 84.950 35.250 85.350 35.650 ;
        RECT 85.850 35.250 86.250 35.650 ;
        RECT 89.250 35.250 89.650 35.650 ;
        RECT 75.150 31.650 75.550 32.050 ;
        RECT 80.600 31.850 81.000 32.250 ;
        RECT 81.250 31.700 81.650 32.100 ;
        RECT 81.250 30.400 81.450 31.700 ;
        RECT 68.300 29.900 68.700 30.300 ;
        RECT 76.900 29.900 77.300 30.300 ;
        RECT 81.150 30.000 81.550 30.400 ;
        RECT 87.300 29.900 87.700 30.300 ;
        RECT 66.250 29.350 66.650 29.750 ;
        RECT 67.350 29.350 67.750 29.750 ;
        RECT 68.850 29.350 69.250 29.750 ;
        RECT 69.950 29.350 70.350 29.750 ;
        RECT 70.750 29.350 71.150 29.750 ;
        RECT 71.850 29.350 72.250 29.750 ;
        RECT 73.350 29.350 73.750 29.750 ;
        RECT 74.450 29.350 74.850 29.750 ;
        RECT 75.950 29.350 76.350 29.750 ;
        RECT 78.150 29.350 78.550 29.750 ;
        RECT 79.800 29.350 80.200 29.750 ;
        RECT 81.950 29.350 82.350 29.750 ;
        RECT 83.900 29.350 84.300 29.750 ;
        RECT 85.850 29.350 86.250 29.750 ;
        RECT 88.450 29.050 88.850 32.400 ;
        RECT 90.000 31.600 90.400 32.000 ;
        RECT 91.450 31.600 91.850 36.400 ;
        RECT 92.000 29.900 92.400 35.850 ;
        RECT 94.600 34.850 95.000 58.300 ;
        RECT 95.150 42.700 95.550 59.100 ;
        RECT 95.700 51.850 96.100 66.000 ;
        RECT 97.600 63.000 98.000 65.400 ;
        RECT 97.600 61.600 98.000 62.800 ;
        RECT 98.600 61.600 99.000 65.400 ;
        RECT 99.600 61.050 100.000 65.400 ;
        RECT 100.600 61.600 101.000 65.400 ;
        RECT 101.600 63.000 102.000 66.000 ;
        RECT 102.600 61.600 103.000 65.400 ;
        RECT 103.600 63.000 104.000 66.000 ;
        RECT 104.600 62.000 105.000 65.400 ;
        RECT 105.600 62.300 106.000 65.400 ;
        RECT 104.600 61.600 105.400 62.000 ;
        RECT 106.600 61.600 107.000 65.400 ;
        RECT 107.600 61.600 108.000 65.400 ;
        RECT 110.600 61.600 111.000 62.000 ;
        RECT 97.250 59.750 97.650 60.650 ;
        RECT 97.900 59.750 98.300 60.650 ;
        RECT 98.550 59.750 98.950 60.650 ;
        RECT 99.200 59.750 99.600 60.650 ;
        RECT 99.850 59.750 100.250 60.650 ;
        RECT 100.500 59.750 100.900 60.650 ;
        RECT 101.150 59.750 101.550 60.650 ;
        RECT 102.950 59.750 103.350 60.650 ;
        RECT 103.600 59.750 104.000 60.650 ;
        RECT 98.100 59.150 98.500 59.550 ;
        RECT 98.650 57.850 98.850 59.750 ;
        RECT 99.950 58.650 100.150 59.750 ;
        RECT 100.300 59.150 100.700 59.550 ;
        RECT 99.850 58.350 100.250 58.650 ;
        RECT 97.250 56.850 97.650 57.250 ;
        RECT 97.900 56.850 98.300 57.250 ;
        RECT 98.550 56.850 98.950 57.850 ;
        RECT 99.950 57.450 100.150 58.350 ;
        RECT 100.400 58.200 100.600 59.150 ;
        RECT 104.250 59.100 104.650 60.650 ;
        RECT 104.900 59.750 105.300 60.650 ;
        RECT 105.550 59.750 105.950 60.650 ;
        RECT 106.200 59.750 106.600 60.650 ;
        RECT 106.850 59.750 107.250 60.650 ;
        RECT 105.650 59.450 105.850 59.750 ;
        RECT 103.600 58.750 104.000 59.050 ;
        RECT 100.300 57.800 100.700 58.200 ;
        RECT 103.800 57.850 104.000 58.750 ;
        RECT 103.800 57.450 104.200 57.850 ;
        RECT 99.200 56.850 99.600 57.250 ;
        RECT 99.850 56.850 100.250 57.450 ;
        RECT 104.350 57.250 104.550 59.100 ;
        RECT 105.650 59.050 106.050 59.450 ;
        RECT 109.500 59.150 109.900 59.550 ;
        RECT 113.700 59.150 114.100 59.550 ;
        RECT 116.100 59.150 116.500 62.200 ;
        RECT 105.650 57.250 105.850 59.050 ;
        RECT 109.500 58.050 109.900 58.450 ;
        RECT 110.150 58.300 110.550 58.700 ;
        RECT 111.150 58.300 111.550 58.700 ;
        RECT 106.000 57.450 106.400 57.850 ;
        RECT 113.700 57.450 114.100 57.850 ;
        RECT 100.500 56.850 100.900 57.250 ;
        RECT 101.150 56.850 101.550 57.250 ;
        RECT 102.950 56.850 103.350 57.250 ;
        RECT 103.600 56.850 104.000 57.250 ;
        RECT 104.250 56.850 104.650 57.250 ;
        RECT 104.900 56.850 105.300 57.250 ;
        RECT 105.550 56.850 105.950 57.250 ;
        RECT 106.200 56.850 106.600 57.250 ;
        RECT 106.850 56.850 107.250 57.250 ;
        RECT 97.000 54.750 97.400 55.900 ;
        RECT 98.000 53.400 98.400 55.900 ;
        RECT 99.200 55.500 99.600 55.900 ;
        RECT 100.000 53.400 100.400 55.900 ;
        RECT 102.000 53.400 102.400 55.900 ;
        RECT 104.000 53.400 104.400 55.900 ;
        RECT 104.900 54.950 105.300 56.450 ;
        RECT 106.000 53.400 106.400 55.900 ;
        RECT 107.000 54.750 107.400 55.900 ;
        RECT 110.600 55.500 111.000 55.900 ;
        RECT 116.100 54.850 116.500 57.850 ;
        RECT 117.700 56.900 118.250 60.000 ;
        RECT 116.170 54.845 116.420 54.850 ;
        RECT 115.050 49.900 115.450 50.300 ;
        RECT 116.050 47.300 116.550 50.800 ;
        RECT 95.700 35.450 96.100 42.550 ;
        RECT 115.450 41.450 116.000 42.000 ;
        RECT 96.700 38.250 97.100 41.200 ;
        RECT 97.800 38.250 98.200 41.200 ;
        RECT 98.900 38.250 99.300 40.150 ;
        RECT 100.000 38.250 100.400 41.200 ;
        RECT 101.600 40.150 102.000 41.200 ;
        RECT 101.100 38.250 102.500 40.150 ;
        RECT 103.200 38.250 103.600 41.200 ;
        RECT 98.900 36.550 99.300 38.100 ;
        RECT 97.700 31.600 98.100 34.650 ;
        RECT 98.800 31.600 99.200 34.650 ;
        RECT 99.900 32.750 100.300 35.250 ;
        RECT 101.000 34.850 101.400 35.850 ;
        RECT 101.000 31.600 101.400 34.650 ;
        RECT 102.100 32.750 102.500 35.250 ;
        RECT 104.300 34.850 104.700 40.150 ;
        RECT 105.400 38.250 105.800 41.200 ;
        RECT 107.000 40.150 107.400 41.200 ;
        RECT 106.500 38.250 107.900 40.150 ;
        RECT 108.600 38.250 109.000 41.200 ;
        RECT 109.050 37.500 109.450 37.900 ;
        RECT 106.850 35.000 107.250 36.400 ;
        RECT 103.200 31.600 103.600 34.650 ;
        RECT 104.300 32.750 105.700 34.650 ;
        RECT 104.800 31.600 105.200 32.750 ;
        RECT 106.400 31.600 106.800 34.650 ;
        RECT 107.500 32.750 107.900 35.250 ;
        RECT 108.600 31.600 109.000 34.650 ;
        RECT 109.700 32.750 110.100 40.150 ;
        RECT 110.800 38.250 111.200 41.200 ;
        RECT 111.900 38.250 112.300 41.200 ;
        RECT 110.350 37.500 110.750 37.900 ;
        RECT 113.700 37.500 114.250 38.050 ;
        RECT 110.350 35.000 110.750 35.400 ;
        RECT 113.700 34.850 114.250 35.400 ;
        RECT 110.800 31.600 111.200 34.650 ;
        RECT 111.900 31.600 112.300 34.650 ;
        RECT 114.900 28.950 115.450 29.500 ;
        RECT 117.900 27.350 118.300 28.250 ;
        RECT 120.500 27.350 120.900 28.250 ;
        RECT 123.100 27.350 123.500 28.250 ;
        RECT 125.700 27.350 126.100 28.250 ;
        RECT 116.050 20.750 116.350 27.100 ;
        RECT 116.950 24.600 117.350 25.000 ;
        RECT 117.950 24.100 118.250 27.350 ;
        RECT 116.550 23.700 116.950 24.100 ;
        RECT 117.900 23.700 118.300 24.100 ;
        RECT 116.600 20.750 116.900 23.700 ;
        RECT 117.050 20.750 117.450 21.150 ;
        RECT 116.050 19.750 116.250 20.750 ;
        RECT 116.400 20.200 116.690 20.550 ;
        RECT 63.300 18.350 63.700 18.750 ;
        RECT 65.400 18.350 65.800 18.750 ;
        RECT 68.750 18.350 69.150 18.750 ;
        RECT 71.600 18.350 72.000 18.750 ;
        RECT 75.350 18.350 75.750 18.750 ;
        RECT 77.500 18.350 77.900 18.750 ;
        RECT 79.700 18.350 80.100 18.750 ;
        RECT 80.950 18.350 81.350 18.750 ;
        RECT 82.050 18.350 82.450 18.750 ;
        RECT 84.400 18.350 84.800 18.750 ;
        RECT 86.600 18.350 87.000 18.750 ;
        RECT 89.700 18.350 90.100 18.750 ;
        RECT 91.400 18.350 91.800 18.750 ;
        RECT 93.200 18.350 93.600 18.750 ;
        RECT 96.200 18.350 96.600 18.750 ;
        RECT 97.900 18.350 98.300 18.750 ;
        RECT 99.700 18.350 100.100 18.750 ;
        RECT 102.700 18.350 103.100 18.750 ;
        RECT 104.400 18.350 104.800 18.750 ;
        RECT 106.200 18.350 106.600 18.750 ;
        RECT 109.200 18.350 109.600 18.750 ;
        RECT 110.900 18.350 111.300 18.750 ;
        RECT 112.700 18.350 113.100 18.750 ;
        RECT 64.900 18.000 65.300 18.200 ;
        RECT 65.900 18.000 66.250 18.200 ;
        RECT 64.900 17.800 66.250 18.000 ;
        RECT 66.450 18.000 66.850 18.100 ;
        RECT 70.500 18.000 70.900 18.200 ;
        RECT 66.450 17.800 70.900 18.000 ;
        RECT 71.200 18.000 71.500 18.200 ;
        RECT 77.000 18.000 77.400 18.200 ;
        RECT 78.100 18.000 78.500 18.200 ;
        RECT 71.200 17.800 73.850 18.000 ;
        RECT 77.000 17.800 78.500 18.000 ;
        RECT 83.750 18.050 84.150 18.200 ;
        RECT 85.800 18.050 86.200 18.200 ;
        RECT 83.750 17.850 86.200 18.050 ;
        RECT 95.550 18.000 95.950 18.200 ;
        RECT 98.450 18.000 98.850 18.200 ;
        RECT 95.550 17.800 98.850 18.000 ;
        RECT 102.050 18.000 102.450 18.200 ;
        RECT 104.950 18.000 105.350 18.200 ;
        RECT 102.050 17.800 105.350 18.000 ;
        RECT 108.550 18.000 108.950 18.200 ;
        RECT 111.450 18.000 111.850 18.200 ;
        RECT 108.550 17.800 111.850 18.000 ;
        RECT 116.040 17.850 116.340 19.750 ;
        RECT 116.600 17.800 116.900 19.750 ;
        RECT 66.450 17.700 66.850 17.800 ;
        RECT 73.650 17.600 73.850 17.800 ;
        RECT 95.750 17.600 95.950 17.800 ;
        RECT 102.250 17.600 102.450 17.800 ;
        RECT 108.750 17.600 108.950 17.800 ;
        RECT 73.650 17.200 74.050 17.600 ;
        RECT 116.260 17.300 116.550 17.650 ;
        RECT 116.300 17.100 116.550 17.300 ;
        RECT 61.200 16.350 61.600 16.750 ;
        RECT 114.050 16.700 115.250 17.100 ;
        RECT 69.750 16.350 72.750 16.550 ;
        RECT 69.750 16.200 70.150 16.350 ;
        RECT 72.350 16.200 72.750 16.350 ;
        RECT 81.150 16.250 81.550 16.650 ;
        RECT 113.760 16.300 115.250 16.700 ;
        RECT 61.500 15.300 61.900 15.400 ;
        RECT 66.450 15.300 66.850 15.500 ;
        RECT 81.150 15.400 81.350 16.250 ;
        RECT 61.500 15.100 66.850 15.300 ;
        RECT 67.100 15.250 67.500 15.400 ;
        RECT 71.800 15.250 72.200 15.400 ;
        RECT 79.800 15.250 80.200 15.400 ;
        RECT 61.500 15.000 61.900 15.100 ;
        RECT 67.100 15.050 80.200 15.250 ;
        RECT 81.150 15.200 93.200 15.400 ;
        RECT 92.870 15.000 93.200 15.200 ;
        RECT 62.500 14.450 62.900 14.850 ;
        RECT 63.600 14.450 64.000 14.850 ;
        RECT 65.950 14.450 66.350 14.850 ;
        RECT 67.650 14.450 68.050 14.850 ;
        RECT 68.750 14.450 69.150 14.850 ;
        RECT 70.950 14.450 71.350 14.850 ;
        RECT 73.300 14.450 73.700 14.850 ;
        RECT 74.550 14.450 74.950 14.850 ;
        RECT 75.650 14.450 76.050 14.850 ;
        RECT 78.000 14.450 78.400 14.850 ;
        RECT 80.300 14.450 80.700 14.850 ;
        RECT 82.050 14.450 82.450 14.850 ;
        RECT 83.300 14.450 83.700 14.850 ;
        RECT 84.400 14.450 84.800 14.850 ;
        RECT 86.050 14.450 86.450 14.850 ;
        RECT 89.350 14.450 89.750 14.850 ;
        RECT 90.450 14.450 90.850 14.850 ;
        RECT 93.300 14.450 93.700 14.850 ;
        RECT 94.600 14.450 95.000 14.850 ;
        RECT 95.850 14.450 96.250 14.850 ;
        RECT 96.950 14.450 97.350 14.850 ;
        RECT 99.700 14.450 100.100 14.850 ;
        RECT 101.100 14.450 101.500 14.850 ;
        RECT 102.350 14.450 102.750 14.850 ;
        RECT 103.450 14.450 103.850 14.850 ;
        RECT 106.200 14.450 106.600 14.850 ;
        RECT 107.600 14.450 108.000 14.850 ;
        RECT 108.850 14.450 109.250 14.850 ;
        RECT 109.950 14.450 110.350 14.850 ;
        RECT 112.700 14.450 113.100 14.850 ;
        RECT 114.050 8.000 115.250 16.300 ;
        RECT 116.250 15.900 116.550 17.100 ;
        RECT 116.300 15.700 116.550 15.900 ;
        RECT 116.260 15.350 116.550 15.700 ;
        RECT 116.700 17.100 116.900 17.800 ;
        RECT 116.700 15.900 117.000 17.100 ;
        RECT 116.700 15.150 116.900 15.900 ;
        RECT 115.850 14.250 116.340 15.150 ;
        RECT 116.600 14.250 116.900 15.150 ;
        RECT 115.850 14.000 116.060 14.250 ;
        RECT 115.850 13.250 116.050 14.000 ;
        RECT 117.150 13.850 117.450 20.750 ;
        RECT 118.650 20.750 118.950 27.100 ;
        RECT 119.550 24.600 119.950 25.000 ;
        RECT 120.550 24.100 120.850 27.350 ;
        RECT 119.150 23.700 119.550 24.100 ;
        RECT 120.500 23.700 120.900 24.100 ;
        RECT 119.200 20.750 119.500 23.700 ;
        RECT 119.650 20.750 120.050 21.150 ;
        RECT 116.400 13.450 116.690 13.800 ;
        RECT 117.050 13.450 117.450 13.850 ;
        RECT 115.850 11.850 116.350 13.250 ;
        RECT 116.600 11.850 117.100 13.250 ;
        RECT 117.600 12.850 118.000 20.550 ;
        RECT 118.650 19.750 118.850 20.750 ;
        RECT 119.000 20.200 119.290 20.550 ;
        RECT 118.640 17.850 118.940 19.750 ;
        RECT 119.200 17.800 119.500 19.750 ;
        RECT 118.860 17.300 119.150 17.650 ;
        RECT 118.900 17.100 119.150 17.300 ;
        RECT 118.850 15.900 119.150 17.100 ;
        RECT 118.900 15.700 119.150 15.900 ;
        RECT 118.860 15.350 119.150 15.700 ;
        RECT 119.300 17.100 119.500 17.800 ;
        RECT 119.300 15.900 119.600 17.100 ;
        RECT 119.300 15.150 119.500 15.900 ;
        RECT 118.450 14.250 118.940 15.150 ;
        RECT 119.200 14.250 119.500 15.150 ;
        RECT 118.450 14.000 118.660 14.250 ;
        RECT 118.450 13.250 118.650 14.000 ;
        RECT 119.750 13.850 120.050 20.750 ;
        RECT 121.250 20.750 121.550 27.100 ;
        RECT 122.150 24.600 122.550 25.000 ;
        RECT 123.150 24.100 123.450 27.350 ;
        RECT 123.850 24.600 124.150 27.100 ;
        RECT 125.750 25.200 126.050 27.350 ;
        RECT 121.750 23.700 122.150 24.100 ;
        RECT 123.100 23.700 123.500 24.100 ;
        RECT 121.800 20.750 122.100 23.700 ;
        RECT 122.250 20.750 122.650 21.150 ;
        RECT 119.000 13.450 119.290 13.800 ;
        RECT 119.650 13.450 120.050 13.850 ;
        RECT 115.850 10.850 116.050 11.850 ;
        RECT 116.330 11.050 116.620 11.400 ;
        RECT 116.900 10.850 117.100 11.850 ;
        RECT 115.850 9.950 116.350 10.850 ;
        RECT 116.600 9.950 117.100 10.850 ;
        RECT 118.450 11.850 118.950 13.250 ;
        RECT 119.200 11.850 119.700 13.250 ;
        RECT 120.200 12.850 120.600 20.550 ;
        RECT 121.250 19.750 121.450 20.750 ;
        RECT 121.600 20.200 121.890 20.550 ;
        RECT 121.240 17.850 121.540 19.750 ;
        RECT 121.800 17.800 122.100 19.750 ;
        RECT 121.460 17.300 121.750 17.650 ;
        RECT 121.500 17.100 121.750 17.300 ;
        RECT 121.450 15.900 121.750 17.100 ;
        RECT 121.500 15.700 121.750 15.900 ;
        RECT 121.460 15.350 121.750 15.700 ;
        RECT 121.900 17.100 122.100 17.800 ;
        RECT 121.900 15.900 122.200 17.100 ;
        RECT 121.900 15.150 122.100 15.900 ;
        RECT 121.050 14.250 121.540 15.150 ;
        RECT 121.800 14.250 122.100 15.150 ;
        RECT 121.050 14.000 121.260 14.250 ;
        RECT 121.050 13.250 121.250 14.000 ;
        RECT 122.350 13.850 122.650 20.750 ;
        RECT 121.600 13.450 121.890 13.800 ;
        RECT 122.250 13.450 122.650 13.850 ;
        RECT 118.450 10.850 118.650 11.850 ;
        RECT 118.930 11.050 119.220 11.400 ;
        RECT 119.500 10.850 119.700 11.850 ;
        RECT 118.450 9.950 118.950 10.850 ;
        RECT 119.200 9.950 119.700 10.850 ;
        RECT 121.050 11.850 121.550 13.250 ;
        RECT 121.800 11.850 122.300 13.250 ;
        RECT 122.800 12.850 123.200 20.550 ;
        RECT 121.050 10.850 121.250 11.850 ;
        RECT 121.530 11.050 121.820 11.400 ;
        RECT 122.100 10.850 122.300 11.850 ;
        RECT 124.370 11.050 124.660 11.400 ;
        RECT 121.050 9.950 121.550 10.850 ;
        RECT 121.800 9.950 122.300 10.850 ;
        RECT 116.600 9.700 116.900 9.950 ;
        RECT 119.200 9.700 119.500 9.950 ;
        RECT 121.800 9.700 122.100 9.950 ;
        RECT 124.250 9.700 124.550 10.850 ;
        RECT 124.800 9.950 125.100 25.000 ;
        RECT 116.550 7.450 116.950 9.700 ;
        RECT 119.150 7.450 119.550 9.700 ;
        RECT 121.750 7.450 122.150 9.700 ;
        RECT 124.200 7.450 124.600 9.700 ;
        RECT 125.850 8.000 127.050 17.100 ;
        RECT 130.000 11.050 132.400 99.100 ;
        RECT 132.550 42.150 132.950 58.700 ;
      LAYER met2 ;
        RECT 37.300 101.050 38.600 101.450 ;
        RECT 37.300 100.500 117.050 101.050 ;
        RECT 37.300 100.150 38.600 100.500 ;
        RECT 80.600 100.100 81.000 100.500 ;
        RECT 44.600 99.550 45.100 99.600 ;
        RECT 129.950 99.550 132.400 99.600 ;
        RECT 44.600 99.150 77.100 99.550 ;
        RECT 84.500 99.150 132.400 99.550 ;
        RECT 44.600 99.100 45.100 99.150 ;
        RECT 129.950 99.100 132.400 99.150 ;
        RECT 45.850 97.600 91.350 98.000 ;
        RECT 37.300 96.250 88.250 97.450 ;
        RECT 90.950 95.900 91.350 96.300 ;
        RECT 43.850 92.150 46.250 94.300 ;
        RECT 87.750 92.150 90.150 94.300 ;
        RECT 93.200 92.350 93.700 92.850 ;
        RECT 90.600 88.900 91.000 89.300 ;
        RECT 55.700 85.700 58.250 86.100 ;
        RECT 66.200 85.700 77.100 86.100 ;
        RECT 87.800 85.350 94.400 85.850 ;
        RECT 89.750 81.900 95.350 82.300 ;
        RECT 81.750 78.350 94.400 78.850 ;
        RECT 76.700 75.650 81.600 76.050 ;
        RECT 51.750 75.250 75.100 75.650 ;
        RECT 55.700 73.700 59.900 74.100 ;
        RECT 72.900 73.700 81.150 74.100 ;
        RECT 75.500 73.150 78.950 73.550 ;
        RECT 48.400 72.100 84.300 72.500 ;
        RECT 53.100 71.550 93.650 71.950 ;
        RECT 47.300 70.700 55.800 71.100 ;
        RECT 77.350 70.500 92.900 71.300 ;
        RECT 55.800 70.150 56.200 70.250 ;
        RECT 56.600 70.150 57.000 70.250 ;
        RECT 57.400 70.150 57.800 70.250 ;
        RECT 58.200 70.150 58.600 70.250 ;
        RECT 59.000 70.150 59.400 70.250 ;
        RECT 59.800 70.150 60.200 70.250 ;
        RECT 60.600 70.150 61.000 70.250 ;
        RECT 61.400 70.150 61.800 70.250 ;
        RECT 62.200 70.150 62.600 70.250 ;
        RECT 63.000 70.150 63.400 70.250 ;
        RECT 63.800 70.150 64.200 70.250 ;
        RECT 64.600 70.150 65.000 70.250 ;
        RECT 65.400 70.150 65.800 70.250 ;
        RECT 55.800 69.950 65.800 70.150 ;
        RECT 55.800 69.850 56.200 69.950 ;
        RECT 56.600 69.850 57.000 69.950 ;
        RECT 57.400 69.850 57.800 69.950 ;
        RECT 58.200 69.850 58.600 69.950 ;
        RECT 59.000 69.850 59.400 69.950 ;
        RECT 59.800 69.850 60.200 69.950 ;
        RECT 60.600 69.850 61.000 69.950 ;
        RECT 61.400 69.850 61.800 69.950 ;
        RECT 62.200 69.850 62.600 69.950 ;
        RECT 63.000 69.850 63.400 69.950 ;
        RECT 63.800 69.850 64.200 69.950 ;
        RECT 64.600 69.850 65.000 69.950 ;
        RECT 65.400 69.850 65.800 69.950 ;
        RECT 66.200 70.150 66.600 70.250 ;
        RECT 67.000 70.150 67.400 70.250 ;
        RECT 67.800 70.150 68.200 70.250 ;
        RECT 68.600 70.150 69.000 70.250 ;
        RECT 69.400 70.150 69.800 70.250 ;
        RECT 70.200 70.150 70.600 70.250 ;
        RECT 71.000 70.150 71.400 70.250 ;
        RECT 71.800 70.150 72.200 70.250 ;
        RECT 72.600 70.150 73.000 70.250 ;
        RECT 73.400 70.150 73.800 70.250 ;
        RECT 74.200 70.150 74.600 70.250 ;
        RECT 75.000 70.150 75.400 70.250 ;
        RECT 75.800 70.150 76.200 70.250 ;
        RECT 66.200 69.950 76.200 70.150 ;
        RECT 66.200 69.850 66.600 69.950 ;
        RECT 67.000 69.850 67.400 69.950 ;
        RECT 67.800 69.850 68.200 69.950 ;
        RECT 68.600 69.850 69.000 69.950 ;
        RECT 69.400 69.850 69.800 69.950 ;
        RECT 70.200 69.850 70.600 69.950 ;
        RECT 71.000 69.850 71.400 69.950 ;
        RECT 71.800 69.850 72.200 69.950 ;
        RECT 72.600 69.850 73.000 69.950 ;
        RECT 73.400 69.850 73.800 69.950 ;
        RECT 74.200 69.850 74.600 69.950 ;
        RECT 75.000 69.850 75.400 69.950 ;
        RECT 75.800 69.850 76.200 69.950 ;
        RECT 59.500 68.500 92.900 69.700 ;
        RECT 116.050 69.150 116.550 69.650 ;
        RECT 91.700 67.550 115.450 67.950 ;
        RECT 90.200 66.700 91.400 67.200 ;
        RECT 54.600 64.500 91.400 65.700 ;
        RECT 95.700 65.600 104.000 66.000 ;
        RECT 53.700 63.950 62.650 64.350 ;
        RECT 70.150 63.950 79.100 64.350 ;
        RECT 48.400 63.450 62.245 63.800 ;
        RECT 48.400 63.400 48.800 63.450 ;
        RECT 47.850 62.300 62.750 62.650 ;
        RECT 64.000 62.500 68.800 63.700 ;
        RECT 70.555 63.450 81.150 63.800 ;
        RECT 80.750 63.400 81.150 63.450 ;
        RECT 70.050 62.300 81.600 62.650 ;
        RECT 99.600 62.300 106.000 62.700 ;
        RECT 47.850 62.250 48.250 62.300 ;
        RECT 81.200 62.250 81.600 62.300 ;
        RECT 58.000 61.750 63.200 62.150 ;
        RECT 69.600 61.750 74.800 62.150 ;
        RECT 90.200 62.000 91.400 62.050 ;
        RECT 90.200 61.600 111.000 62.000 ;
        RECT 56.800 61.200 62.000 61.600 ;
        RECT 70.800 61.200 76.000 61.600 ;
        RECT 90.200 61.550 91.400 61.600 ;
        RECT 99.600 61.050 100.000 61.450 ;
        RECT 53.100 59.850 64.100 60.250 ;
        RECT 68.700 59.850 82.950 61.050 ;
        RECT 54.400 59.550 54.800 59.650 ;
        RECT 58.000 59.550 58.400 59.650 ;
        RECT 61.600 59.550 62.000 59.650 ;
        RECT 54.400 59.350 62.000 59.550 ;
        RECT 54.400 59.250 54.800 59.350 ;
        RECT 58.000 59.250 58.400 59.350 ;
        RECT 61.600 59.250 62.000 59.350 ;
        RECT 70.800 59.550 71.200 59.650 ;
        RECT 74.400 59.550 74.800 59.650 ;
        RECT 78.000 59.550 78.400 59.650 ;
        RECT 70.800 59.350 78.400 59.550 ;
        RECT 70.800 59.250 71.200 59.350 ;
        RECT 74.400 59.250 74.800 59.350 ;
        RECT 78.000 59.250 78.400 59.350 ;
        RECT 95.150 59.000 95.550 59.100 ;
        RECT 98.100 59.000 98.500 59.550 ;
        RECT 100.300 59.150 100.700 59.550 ;
        RECT 105.650 59.350 106.050 59.450 ;
        RECT 109.500 59.350 109.900 59.550 ;
        RECT 105.650 59.150 109.900 59.350 ;
        RECT 113.700 59.150 116.500 59.550 ;
        RECT 117.700 59.450 118.250 60.000 ;
        RECT 105.650 59.050 106.050 59.150 ;
        RECT 103.600 59.000 104.000 59.050 ;
        RECT 95.150 58.800 104.000 59.000 ;
        RECT 95.150 58.700 95.550 58.800 ;
        RECT 103.600 58.750 104.000 58.800 ;
        RECT 99.850 58.600 100.250 58.650 ;
        RECT 99.850 58.400 109.900 58.600 ;
        RECT 99.850 58.350 100.250 58.400 ;
        RECT 94.600 58.200 95.000 58.300 ;
        RECT 56.850 57.950 57.150 58.100 ;
        RECT 75.650 57.950 75.950 58.150 ;
        RECT 94.600 58.000 106.400 58.200 ;
        RECT 109.500 58.050 109.900 58.400 ;
        RECT 110.150 58.300 132.950 58.700 ;
        RECT 43.950 57.550 65.700 57.950 ;
        RECT 67.100 57.550 88.250 57.950 ;
        RECT 94.600 57.900 95.000 58.000 ;
        RECT 100.300 57.800 100.700 58.000 ;
        RECT 103.800 57.450 104.200 57.850 ;
        RECT 106.000 57.450 106.400 58.000 ;
        RECT 113.700 57.450 116.500 57.850 ;
        RECT 52.600 56.200 91.400 57.400 ;
        RECT 117.700 56.900 118.250 57.450 ;
        RECT 104.900 56.050 105.300 56.450 ;
        RECT 47.850 55.650 73.800 56.050 ;
        RECT 91.700 55.900 92.900 55.950 ;
        RECT 91.700 55.500 111.000 55.900 ;
        RECT 47.300 55.100 78.950 55.500 ;
        RECT 91.700 55.450 92.900 55.500 ;
        RECT 104.900 54.950 105.300 55.350 ;
        RECT 62.600 54.550 81.600 54.950 ;
        RECT 64.400 54.000 81.150 54.400 ;
        RECT 59.500 53.450 73.300 53.850 ;
        RECT 77.950 52.450 79.550 52.850 ;
        RECT 76.200 51.050 76.600 51.150 ;
        RECT 78.550 51.050 78.950 51.150 ;
        RECT 76.200 50.850 78.950 51.050 ;
        RECT 76.200 50.750 76.600 50.850 ;
        RECT 78.550 50.750 78.950 50.850 ;
        RECT 58.100 48.950 91.400 50.150 ;
        RECT 91.700 49.900 115.450 50.300 ;
        RECT 43.950 48.450 73.770 48.800 ;
        RECT 116.050 47.300 116.550 47.800 ;
        RECT 90.200 47.150 91.400 47.200 ;
        RECT 58.150 46.750 91.400 47.150 ;
        RECT 90.200 46.700 91.400 46.750 ;
        RECT 48.400 46.200 64.600 46.600 ;
        RECT 68.200 45.350 94.450 46.550 ;
        RECT 95.150 42.700 132.400 43.900 ;
        RECT 95.700 42.150 132.950 42.550 ;
        RECT 64.550 41.550 65.050 41.950 ;
        RECT 115.450 41.900 116.000 42.000 ;
        RECT 64.550 41.150 89.650 41.550 ;
        RECT 90.500 41.500 116.000 41.900 ;
        RECT 115.450 41.450 116.000 41.500 ;
        RECT 64.550 40.750 65.050 41.150 ;
        RECT 84.500 40.600 84.900 41.000 ;
        RECT 87.650 40.600 90.900 41.000 ;
        RECT 91.700 40.800 112.300 41.200 ;
        RECT 60.250 38.700 66.050 39.100 ;
        RECT 75.250 38.650 75.650 39.050 ;
        RECT 80.400 38.650 80.800 39.050 ;
        RECT 90.000 38.900 91.300 39.300 ;
        RECT 113.700 37.900 114.250 38.050 ;
        RECT 109.050 37.500 109.450 37.900 ;
        RECT 110.350 37.500 114.250 37.900 ;
        RECT 90.900 37.100 109.450 37.500 ;
        RECT 90.900 36.550 99.300 36.950 ;
        RECT 68.500 36.100 68.900 36.200 ;
        RECT 76.150 36.150 76.550 36.200 ;
        RECT 81.150 36.150 81.550 36.250 ;
        RECT 76.150 36.100 81.550 36.150 ;
        RECT 64.550 35.650 65.050 36.050 ;
        RECT 68.500 35.950 81.550 36.100 ;
        RECT 68.500 35.900 76.550 35.950 ;
        RECT 68.500 35.800 68.900 35.900 ;
        RECT 76.150 35.800 76.550 35.900 ;
        RECT 81.150 35.850 81.550 35.950 ;
        RECT 83.250 36.100 83.650 36.150 ;
        RECT 84.100 36.100 84.500 36.200 ;
        RECT 83.250 35.900 84.500 36.100 ;
        RECT 83.250 35.850 83.650 35.900 ;
        RECT 84.100 35.850 84.500 35.900 ;
        RECT 87.300 35.800 91.300 36.200 ;
        RECT 91.450 36.000 107.250 36.400 ;
        RECT 109.700 36.250 132.400 36.650 ;
        RECT 64.550 35.250 89.650 35.650 ;
        RECT 92.000 35.450 101.400 35.850 ;
        RECT 64.550 34.850 65.050 35.250 ;
        RECT 76.250 34.700 76.650 35.050 ;
        RECT 94.600 34.850 104.700 35.250 ;
        RECT 106.850 35.000 107.250 35.400 ;
        RECT 107.500 34.850 110.100 35.250 ;
        RECT 110.350 35.000 114.250 35.400 ;
        RECT 113.700 34.850 114.250 35.000 ;
        RECT 59.700 31.800 66.050 32.200 ;
        RECT 75.150 31.650 75.550 32.050 ;
        RECT 80.600 31.850 81.000 32.250 ;
        RECT 88.450 32.000 88.850 32.400 ;
        RECT 90.000 31.600 91.850 32.000 ;
        RECT 96.200 31.600 112.300 32.000 ;
        RECT 81.150 30.300 81.550 30.400 ;
        RECT 64.550 29.750 65.050 30.150 ;
        RECT 68.300 30.100 81.550 30.300 ;
        RECT 68.300 29.900 68.700 30.100 ;
        RECT 76.900 29.900 77.300 30.100 ;
        RECT 81.150 30.000 81.550 30.100 ;
        RECT 87.300 29.900 92.400 30.300 ;
        RECT 64.550 29.350 86.250 29.750 ;
        RECT 114.900 29.450 115.450 29.500 ;
        RECT 64.550 28.950 65.050 29.350 ;
        RECT 88.450 29.050 115.450 29.450 ;
        RECT 114.900 28.950 115.450 29.050 ;
        RECT 112.950 28.250 113.450 28.650 ;
        RECT 112.950 27.850 126.100 28.250 ;
        RECT 112.950 27.450 113.450 27.850 ;
        RECT 116.950 24.600 125.100 25.000 ;
        RECT 116.550 23.700 118.300 24.100 ;
        RECT 119.150 23.700 120.900 24.100 ;
        RECT 121.750 23.700 123.500 24.100 ;
        RECT 116.600 20.750 117.450 21.150 ;
        RECT 119.200 20.750 120.050 21.150 ;
        RECT 121.800 20.750 122.650 21.150 ;
        RECT 116.400 20.200 118.000 20.550 ;
        RECT 119.000 20.200 120.600 20.550 ;
        RECT 121.600 20.200 123.200 20.550 ;
        RECT 117.600 20.150 118.000 20.200 ;
        RECT 120.200 20.150 120.600 20.200 ;
        RECT 122.800 20.150 123.200 20.200 ;
        RECT 60.800 18.750 61.300 19.150 ;
        RECT 60.800 18.350 113.100 18.750 ;
        RECT 60.800 17.950 61.300 18.350 ;
        RECT 60.250 16.350 61.600 16.750 ;
        RECT 114.050 16.700 116.550 17.100 ;
        RECT 113.760 16.300 116.550 16.700 ;
        RECT 114.050 15.900 116.550 16.300 ;
        RECT 116.700 15.900 119.150 17.100 ;
        RECT 119.300 15.900 121.750 17.100 ;
        RECT 121.900 15.900 133.350 17.100 ;
        RECT 60.800 14.850 61.300 15.250 ;
        RECT 60.800 14.450 113.100 14.850 ;
        RECT 60.800 14.050 61.300 14.450 ;
        RECT 117.050 13.800 117.450 13.850 ;
        RECT 119.650 13.800 120.050 13.850 ;
        RECT 122.250 13.800 122.650 13.850 ;
        RECT 116.400 13.450 117.450 13.800 ;
        RECT 119.000 13.450 120.050 13.800 ;
        RECT 121.600 13.450 122.650 13.800 ;
        RECT 116.600 12.850 118.000 13.250 ;
        RECT 119.200 12.850 120.600 13.250 ;
        RECT 121.800 12.850 123.200 13.250 ;
        RECT 116.325 11.050 132.400 11.400 ;
        RECT 112.950 7.850 113.450 8.250 ;
        RECT 114.050 8.000 127.050 9.200 ;
        RECT 112.950 7.450 124.600 7.850 ;
        RECT 112.950 7.050 113.450 7.450 ;
        RECT 151.850 6.700 152.650 6.900 ;
        RECT 59.700 6.300 152.650 6.700 ;
        RECT 151.850 6.100 152.650 6.300 ;
      LAYER met3 ;
        RECT 44.600 102.250 114.700 162.550 ;
        RECT 116.350 102.250 130.450 162.550 ;
        RECT 4.000 100.150 38.600 101.450 ;
        RECT 44.600 99.100 45.100 102.250 ;
        RECT 114.000 100.500 114.550 101.050 ;
        RECT 116.500 100.500 117.050 101.050 ;
        RECT 129.950 99.100 130.450 102.250 ;
        RECT 4.000 96.250 38.600 97.450 ;
        RECT 95.600 96.350 97.900 97.200 ;
        RECT 99.100 96.350 101.400 97.200 ;
        RECT 102.600 96.350 104.900 97.200 ;
        RECT 106.100 96.350 108.400 97.200 ;
        RECT 109.600 96.350 111.900 97.200 ;
        RECT 113.100 96.350 115.400 97.200 ;
        RECT 116.600 96.350 118.900 97.200 ;
        RECT 120.100 96.350 122.400 97.200 ;
        RECT 123.600 96.350 125.900 97.200 ;
        RECT 127.100 96.350 129.400 97.200 ;
        RECT 95.600 96.300 129.400 96.350 ;
        RECT 90.950 95.900 129.400 96.300 ;
        RECT 95.600 95.850 129.400 95.900 ;
        RECT 95.600 94.900 97.900 95.850 ;
        RECT 99.100 94.900 101.400 95.850 ;
        RECT 102.600 94.900 104.900 95.850 ;
        RECT 106.100 94.900 108.400 95.850 ;
        RECT 109.600 94.900 111.900 95.850 ;
        RECT 113.100 94.900 115.400 95.850 ;
        RECT 116.600 94.900 118.900 95.850 ;
        RECT 120.100 94.900 122.400 95.850 ;
        RECT 123.600 94.900 125.900 95.850 ;
        RECT 127.100 94.900 129.400 95.850 ;
        RECT 128.000 93.700 128.500 94.900 ;
        RECT 95.600 92.850 97.900 93.700 ;
        RECT 99.100 92.850 101.400 93.700 ;
        RECT 102.600 92.850 104.900 93.700 ;
        RECT 106.100 92.850 108.400 93.700 ;
        RECT 109.600 92.850 111.900 93.700 ;
        RECT 113.100 92.850 115.400 93.700 ;
        RECT 116.600 92.850 118.900 93.700 ;
        RECT 120.100 92.850 122.400 93.700 ;
        RECT 123.600 92.850 125.900 93.700 ;
        RECT 127.100 92.850 129.400 93.700 ;
        RECT 93.200 92.350 93.700 92.850 ;
        RECT 95.600 92.350 129.400 92.850 ;
        RECT 95.600 91.400 97.900 92.350 ;
        RECT 99.100 91.400 101.400 92.350 ;
        RECT 102.600 91.400 104.900 92.350 ;
        RECT 106.100 91.400 108.400 92.350 ;
        RECT 109.600 91.400 111.900 92.350 ;
        RECT 113.100 91.400 115.400 92.350 ;
        RECT 116.600 91.400 118.900 92.350 ;
        RECT 120.100 91.400 122.400 92.350 ;
        RECT 123.600 91.400 125.900 92.350 ;
        RECT 127.100 91.400 129.400 92.350 ;
        RECT 95.600 89.350 97.900 90.200 ;
        RECT 99.100 89.350 101.400 90.200 ;
        RECT 102.600 89.350 104.900 90.200 ;
        RECT 106.100 89.350 108.400 90.200 ;
        RECT 109.600 89.350 111.900 90.200 ;
        RECT 113.100 89.350 115.400 90.200 ;
        RECT 116.600 89.350 118.900 90.200 ;
        RECT 120.100 89.350 122.400 90.200 ;
        RECT 123.600 89.350 125.900 90.200 ;
        RECT 127.100 89.350 129.400 90.200 ;
        RECT 95.600 89.300 129.400 89.350 ;
        RECT 90.600 88.900 129.400 89.300 ;
        RECT 95.600 88.850 129.400 88.900 ;
        RECT 95.600 87.900 97.900 88.850 ;
        RECT 99.100 87.900 101.400 88.850 ;
        RECT 102.600 87.900 104.900 88.850 ;
        RECT 106.100 87.900 108.400 88.850 ;
        RECT 109.600 87.900 111.900 88.850 ;
        RECT 113.100 87.900 115.400 88.850 ;
        RECT 116.600 87.900 118.900 88.850 ;
        RECT 120.100 87.900 122.400 88.850 ;
        RECT 123.600 87.900 125.900 88.850 ;
        RECT 127.100 87.900 129.400 88.850 ;
        RECT 128.000 86.700 128.500 87.900 ;
        RECT 95.600 85.850 97.900 86.700 ;
        RECT 99.100 85.850 101.400 86.700 ;
        RECT 102.600 85.850 104.900 86.700 ;
        RECT 106.100 85.850 108.400 86.700 ;
        RECT 109.600 85.850 111.900 86.700 ;
        RECT 113.100 85.850 115.400 86.700 ;
        RECT 116.600 85.850 118.900 86.700 ;
        RECT 120.100 85.850 122.400 86.700 ;
        RECT 123.600 85.850 125.900 86.700 ;
        RECT 127.100 85.850 129.400 86.700 ;
        RECT 93.900 85.350 94.400 85.850 ;
        RECT 95.600 85.350 129.400 85.850 ;
        RECT 95.600 84.400 97.900 85.350 ;
        RECT 99.100 84.400 101.400 85.350 ;
        RECT 102.600 84.400 104.900 85.350 ;
        RECT 106.100 84.400 108.400 85.350 ;
        RECT 109.600 84.400 111.900 85.350 ;
        RECT 113.100 84.400 115.400 85.350 ;
        RECT 116.600 84.400 118.900 85.350 ;
        RECT 120.100 84.400 122.400 85.350 ;
        RECT 123.600 84.400 125.900 85.350 ;
        RECT 127.100 84.400 129.400 85.350 ;
        RECT 95.600 82.350 97.900 83.200 ;
        RECT 99.100 82.350 101.400 83.200 ;
        RECT 102.600 82.350 104.900 83.200 ;
        RECT 106.100 82.350 108.400 83.200 ;
        RECT 109.600 82.350 111.900 83.200 ;
        RECT 113.100 82.350 115.400 83.200 ;
        RECT 116.600 82.350 118.900 83.200 ;
        RECT 120.100 82.350 122.400 83.200 ;
        RECT 123.600 82.350 125.900 83.200 ;
        RECT 127.100 82.350 129.400 83.200 ;
        RECT 95.600 82.300 129.400 82.350 ;
        RECT 94.950 81.900 129.400 82.300 ;
        RECT 95.600 81.850 129.400 81.900 ;
        RECT 95.600 80.900 97.900 81.850 ;
        RECT 99.100 80.900 101.400 81.850 ;
        RECT 102.600 80.900 104.900 81.850 ;
        RECT 106.100 80.900 108.400 81.850 ;
        RECT 109.600 80.900 111.900 81.850 ;
        RECT 113.100 80.900 115.400 81.850 ;
        RECT 116.600 80.900 118.900 81.850 ;
        RECT 120.100 80.900 122.400 81.850 ;
        RECT 123.600 80.900 125.900 81.850 ;
        RECT 127.100 80.900 129.400 81.850 ;
        RECT 128.000 79.700 128.500 80.900 ;
        RECT 95.600 78.850 97.900 79.700 ;
        RECT 99.100 78.850 101.400 79.700 ;
        RECT 102.600 78.850 104.900 79.700 ;
        RECT 106.100 78.850 108.400 79.700 ;
        RECT 109.600 78.850 111.900 79.700 ;
        RECT 113.100 78.850 115.400 79.700 ;
        RECT 116.600 78.850 118.900 79.700 ;
        RECT 120.100 78.850 122.400 79.700 ;
        RECT 123.600 78.850 125.900 79.700 ;
        RECT 127.100 78.850 129.400 79.700 ;
        RECT 93.900 78.350 94.400 78.850 ;
        RECT 95.600 78.350 129.400 78.850 ;
        RECT 95.600 77.400 97.900 78.350 ;
        RECT 99.100 77.400 101.400 78.350 ;
        RECT 102.600 77.400 104.900 78.350 ;
        RECT 106.100 77.400 108.400 78.350 ;
        RECT 109.600 77.400 111.900 78.350 ;
        RECT 113.100 77.400 115.400 78.350 ;
        RECT 116.600 77.400 118.900 78.350 ;
        RECT 120.100 77.400 122.400 78.350 ;
        RECT 123.600 77.400 125.900 78.350 ;
        RECT 127.100 77.400 129.400 78.350 ;
        RECT 90.200 45.200 91.400 67.200 ;
        RECT 1.000 44.000 91.400 45.200 ;
        RECT 91.700 43.700 92.900 71.300 ;
        RECT 116.050 69.600 116.550 69.650 ;
        RECT 116.050 69.150 129.750 69.600 ;
        RECT 117.700 59.450 118.250 60.000 ;
        RECT 119.450 59.300 129.750 69.150 ;
        RECT 117.700 56.900 118.250 57.450 ;
        RECT 116.050 47.750 116.550 47.800 ;
        RECT 119.450 47.750 129.750 57.600 ;
        RECT 116.050 47.300 129.750 47.750 ;
        RECT 4.000 42.500 92.900 43.700 ;
        RECT 4.000 40.750 65.050 41.950 ;
        RECT 91.700 40.800 92.900 42.500 ;
        RECT 115.450 41.450 116.000 42.000 ;
        RECT 113.700 37.500 114.250 38.050 ;
        RECT 115.450 37.350 118.450 41.450 ;
        RECT 1.000 34.850 65.050 36.050 ;
        RECT 113.700 34.850 114.250 35.400 ;
        RECT 4.000 28.950 65.050 30.150 ;
        RECT 96.200 28.650 97.400 32.000 ;
        RECT 115.450 29.500 120.950 35.550 ;
        RECT 114.900 28.950 120.950 29.500 ;
        RECT 1.000 27.450 113.450 28.650 ;
        RECT 1.000 17.950 61.300 19.150 ;
        RECT 132.550 15.900 133.350 17.100 ;
        RECT 4.000 14.050 61.300 15.250 ;
        RECT 4.000 7.050 113.450 8.250 ;
        RECT 151.850 6.100 152.650 6.900 ;
      LAYER met4 ;
        RECT 114.000 100.500 114.550 102.900 ;
        RECT 116.500 100.500 117.050 102.900 ;
        RECT 96.550 95.850 128.500 96.350 ;
        RECT 128.000 92.850 128.500 95.850 ;
        RECT 93.200 92.350 128.500 92.850 ;
        RECT 96.550 88.850 128.500 89.350 ;
        RECT 128.000 85.850 128.500 88.850 ;
        RECT 93.900 85.350 128.500 85.850 ;
        RECT 96.550 81.850 128.500 82.350 ;
        RECT 128.000 78.850 128.500 81.850 ;
        RECT 93.900 78.350 128.500 78.850 ;
        RECT 117.700 59.450 120.100 60.000 ;
        RECT 117.700 56.900 120.100 57.450 ;
        RECT 113.700 37.500 116.150 38.050 ;
        RECT 113.700 34.850 116.150 35.400 ;
        RECT 132.550 1.000 133.350 17.100 ;
        RECT 151.850 1.000 152.650 6.900 ;
  END
END tt_um_jyblue1001_pll
END LIBRARY

