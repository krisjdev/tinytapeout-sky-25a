module tt_um_regfield (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \thechain[0].chain1.dout ;
 wire \thechain[0].chain1.ff[0] ;
 wire \thechain[0].chain1.ff[10] ;
 wire \thechain[0].chain1.ff[11] ;
 wire \thechain[0].chain1.ff[12] ;
 wire \thechain[0].chain1.ff[13] ;
 wire \thechain[0].chain1.ff[14] ;
 wire \thechain[0].chain1.ff[15] ;
 wire \thechain[0].chain1.ff[16] ;
 wire \thechain[0].chain1.ff[17] ;
 wire \thechain[0].chain1.ff[18] ;
 wire \thechain[0].chain1.ff[19] ;
 wire \thechain[0].chain1.ff[1] ;
 wire \thechain[0].chain1.ff[20] ;
 wire \thechain[0].chain1.ff[21] ;
 wire \thechain[0].chain1.ff[22] ;
 wire \thechain[0].chain1.ff[23] ;
 wire \thechain[0].chain1.ff[24] ;
 wire \thechain[0].chain1.ff[25] ;
 wire \thechain[0].chain1.ff[26] ;
 wire \thechain[0].chain1.ff[27] ;
 wire \thechain[0].chain1.ff[28] ;
 wire \thechain[0].chain1.ff[29] ;
 wire \thechain[0].chain1.ff[2] ;
 wire \thechain[0].chain1.ff[30] ;
 wire \thechain[0].chain1.ff[31] ;
 wire \thechain[0].chain1.ff[32] ;
 wire \thechain[0].chain1.ff[33] ;
 wire \thechain[0].chain1.ff[34] ;
 wire \thechain[0].chain1.ff[35] ;
 wire \thechain[0].chain1.ff[36] ;
 wire \thechain[0].chain1.ff[37] ;
 wire \thechain[0].chain1.ff[38] ;
 wire \thechain[0].chain1.ff[39] ;
 wire \thechain[0].chain1.ff[3] ;
 wire \thechain[0].chain1.ff[40] ;
 wire \thechain[0].chain1.ff[41] ;
 wire \thechain[0].chain1.ff[42] ;
 wire \thechain[0].chain1.ff[43] ;
 wire \thechain[0].chain1.ff[44] ;
 wire \thechain[0].chain1.ff[45] ;
 wire \thechain[0].chain1.ff[46] ;
 wire \thechain[0].chain1.ff[47] ;
 wire \thechain[0].chain1.ff[48] ;
 wire \thechain[0].chain1.ff[49] ;
 wire \thechain[0].chain1.ff[4] ;
 wire \thechain[0].chain1.ff[50] ;
 wire \thechain[0].chain1.ff[51] ;
 wire \thechain[0].chain1.ff[52] ;
 wire \thechain[0].chain1.ff[53] ;
 wire \thechain[0].chain1.ff[54] ;
 wire \thechain[0].chain1.ff[55] ;
 wire \thechain[0].chain1.ff[56] ;
 wire \thechain[0].chain1.ff[57] ;
 wire \thechain[0].chain1.ff[58] ;
 wire \thechain[0].chain1.ff[59] ;
 wire \thechain[0].chain1.ff[5] ;
 wire \thechain[0].chain1.ff[60] ;
 wire \thechain[0].chain1.ff[61] ;
 wire \thechain[0].chain1.ff[62] ;
 wire \thechain[0].chain1.ff[63] ;
 wire \thechain[0].chain1.ff[64] ;
 wire \thechain[0].chain1.ff[65] ;
 wire \thechain[0].chain1.ff[66] ;
 wire \thechain[0].chain1.ff[67] ;
 wire \thechain[0].chain1.ff[68] ;
 wire \thechain[0].chain1.ff[69] ;
 wire \thechain[0].chain1.ff[6] ;
 wire \thechain[0].chain1.ff[70] ;
 wire \thechain[0].chain1.ff[71] ;
 wire \thechain[0].chain1.ff[72] ;
 wire \thechain[0].chain1.ff[73] ;
 wire \thechain[0].chain1.ff[74] ;
 wire \thechain[0].chain1.ff[75] ;
 wire \thechain[0].chain1.ff[76] ;
 wire \thechain[0].chain1.ff[77] ;
 wire \thechain[0].chain1.ff[78] ;
 wire \thechain[0].chain1.ff[7] ;
 wire \thechain[0].chain1.ff[8] ;
 wire \thechain[0].chain1.ff[9] ;
 wire \thechain[0].chain1.flip1[0] ;
 wire \thechain[0].chain1.flip1[10] ;
 wire \thechain[0].chain1.flip1[11] ;
 wire \thechain[0].chain1.flip1[12] ;
 wire \thechain[0].chain1.flip1[13] ;
 wire \thechain[0].chain1.flip1[14] ;
 wire \thechain[0].chain1.flip1[15] ;
 wire \thechain[0].chain1.flip1[16] ;
 wire \thechain[0].chain1.flip1[17] ;
 wire \thechain[0].chain1.flip1[18] ;
 wire \thechain[0].chain1.flip1[19] ;
 wire \thechain[0].chain1.flip1[1] ;
 wire \thechain[0].chain1.flip1[20] ;
 wire \thechain[0].chain1.flip1[21] ;
 wire \thechain[0].chain1.flip1[22] ;
 wire \thechain[0].chain1.flip1[23] ;
 wire \thechain[0].chain1.flip1[24] ;
 wire \thechain[0].chain1.flip1[25] ;
 wire \thechain[0].chain1.flip1[26] ;
 wire \thechain[0].chain1.flip1[27] ;
 wire \thechain[0].chain1.flip1[28] ;
 wire \thechain[0].chain1.flip1[29] ;
 wire \thechain[0].chain1.flip1[2] ;
 wire \thechain[0].chain1.flip1[30] ;
 wire \thechain[0].chain1.flip1[31] ;
 wire \thechain[0].chain1.flip1[32] ;
 wire \thechain[0].chain1.flip1[33] ;
 wire \thechain[0].chain1.flip1[34] ;
 wire \thechain[0].chain1.flip1[35] ;
 wire \thechain[0].chain1.flip1[36] ;
 wire \thechain[0].chain1.flip1[37] ;
 wire \thechain[0].chain1.flip1[38] ;
 wire \thechain[0].chain1.flip1[39] ;
 wire \thechain[0].chain1.flip1[3] ;
 wire \thechain[0].chain1.flip1[40] ;
 wire \thechain[0].chain1.flip1[41] ;
 wire \thechain[0].chain1.flip1[42] ;
 wire \thechain[0].chain1.flip1[43] ;
 wire \thechain[0].chain1.flip1[44] ;
 wire \thechain[0].chain1.flip1[45] ;
 wire \thechain[0].chain1.flip1[46] ;
 wire \thechain[0].chain1.flip1[47] ;
 wire \thechain[0].chain1.flip1[48] ;
 wire \thechain[0].chain1.flip1[49] ;
 wire \thechain[0].chain1.flip1[4] ;
 wire \thechain[0].chain1.flip1[50] ;
 wire \thechain[0].chain1.flip1[51] ;
 wire \thechain[0].chain1.flip1[52] ;
 wire \thechain[0].chain1.flip1[53] ;
 wire \thechain[0].chain1.flip1[54] ;
 wire \thechain[0].chain1.flip1[55] ;
 wire \thechain[0].chain1.flip1[56] ;
 wire \thechain[0].chain1.flip1[57] ;
 wire \thechain[0].chain1.flip1[58] ;
 wire \thechain[0].chain1.flip1[59] ;
 wire \thechain[0].chain1.flip1[5] ;
 wire \thechain[0].chain1.flip1[60] ;
 wire \thechain[0].chain1.flip1[61] ;
 wire \thechain[0].chain1.flip1[62] ;
 wire \thechain[0].chain1.flip1[63] ;
 wire \thechain[0].chain1.flip1[64] ;
 wire \thechain[0].chain1.flip1[65] ;
 wire \thechain[0].chain1.flip1[66] ;
 wire \thechain[0].chain1.flip1[67] ;
 wire \thechain[0].chain1.flip1[68] ;
 wire \thechain[0].chain1.flip1[69] ;
 wire \thechain[0].chain1.flip1[6] ;
 wire \thechain[0].chain1.flip1[70] ;
 wire \thechain[0].chain1.flip1[71] ;
 wire \thechain[0].chain1.flip1[72] ;
 wire \thechain[0].chain1.flip1[73] ;
 wire \thechain[0].chain1.flip1[74] ;
 wire \thechain[0].chain1.flip1[75] ;
 wire \thechain[0].chain1.flip1[76] ;
 wire \thechain[0].chain1.flip1[77] ;
 wire \thechain[0].chain1.flip1[78] ;
 wire \thechain[0].chain1.flip1[79] ;
 wire \thechain[0].chain1.flip1[7] ;
 wire \thechain[0].chain1.flip1[8] ;
 wire \thechain[0].chain1.flip1[9] ;
 wire \thechain[0].chain1.flip2[0] ;
 wire \thechain[0].chain1.flip2[10] ;
 wire \thechain[0].chain1.flip2[11] ;
 wire \thechain[0].chain1.flip2[12] ;
 wire \thechain[0].chain1.flip2[13] ;
 wire \thechain[0].chain1.flip2[14] ;
 wire \thechain[0].chain1.flip2[15] ;
 wire \thechain[0].chain1.flip2[16] ;
 wire \thechain[0].chain1.flip2[17] ;
 wire \thechain[0].chain1.flip2[18] ;
 wire \thechain[0].chain1.flip2[19] ;
 wire \thechain[0].chain1.flip2[1] ;
 wire \thechain[0].chain1.flip2[20] ;
 wire \thechain[0].chain1.flip2[21] ;
 wire \thechain[0].chain1.flip2[22] ;
 wire \thechain[0].chain1.flip2[23] ;
 wire \thechain[0].chain1.flip2[24] ;
 wire \thechain[0].chain1.flip2[25] ;
 wire \thechain[0].chain1.flip2[26] ;
 wire \thechain[0].chain1.flip2[27] ;
 wire \thechain[0].chain1.flip2[28] ;
 wire \thechain[0].chain1.flip2[29] ;
 wire \thechain[0].chain1.flip2[2] ;
 wire \thechain[0].chain1.flip2[30] ;
 wire \thechain[0].chain1.flip2[31] ;
 wire \thechain[0].chain1.flip2[32] ;
 wire \thechain[0].chain1.flip2[33] ;
 wire \thechain[0].chain1.flip2[34] ;
 wire \thechain[0].chain1.flip2[35] ;
 wire \thechain[0].chain1.flip2[36] ;
 wire \thechain[0].chain1.flip2[37] ;
 wire \thechain[0].chain1.flip2[38] ;
 wire \thechain[0].chain1.flip2[39] ;
 wire \thechain[0].chain1.flip2[3] ;
 wire \thechain[0].chain1.flip2[40] ;
 wire \thechain[0].chain1.flip2[41] ;
 wire \thechain[0].chain1.flip2[42] ;
 wire \thechain[0].chain1.flip2[43] ;
 wire \thechain[0].chain1.flip2[44] ;
 wire \thechain[0].chain1.flip2[45] ;
 wire \thechain[0].chain1.flip2[46] ;
 wire \thechain[0].chain1.flip2[47] ;
 wire \thechain[0].chain1.flip2[48] ;
 wire \thechain[0].chain1.flip2[49] ;
 wire \thechain[0].chain1.flip2[4] ;
 wire \thechain[0].chain1.flip2[50] ;
 wire \thechain[0].chain1.flip2[51] ;
 wire \thechain[0].chain1.flip2[52] ;
 wire \thechain[0].chain1.flip2[53] ;
 wire \thechain[0].chain1.flip2[54] ;
 wire \thechain[0].chain1.flip2[55] ;
 wire \thechain[0].chain1.flip2[56] ;
 wire \thechain[0].chain1.flip2[57] ;
 wire \thechain[0].chain1.flip2[58] ;
 wire \thechain[0].chain1.flip2[59] ;
 wire \thechain[0].chain1.flip2[5] ;
 wire \thechain[0].chain1.flip2[60] ;
 wire \thechain[0].chain1.flip2[61] ;
 wire \thechain[0].chain1.flip2[62] ;
 wire \thechain[0].chain1.flip2[63] ;
 wire \thechain[0].chain1.flip2[64] ;
 wire \thechain[0].chain1.flip2[65] ;
 wire \thechain[0].chain1.flip2[66] ;
 wire \thechain[0].chain1.flip2[67] ;
 wire \thechain[0].chain1.flip2[68] ;
 wire \thechain[0].chain1.flip2[69] ;
 wire \thechain[0].chain1.flip2[6] ;
 wire \thechain[0].chain1.flip2[70] ;
 wire \thechain[0].chain1.flip2[71] ;
 wire \thechain[0].chain1.flip2[72] ;
 wire \thechain[0].chain1.flip2[73] ;
 wire \thechain[0].chain1.flip2[74] ;
 wire \thechain[0].chain1.flip2[75] ;
 wire \thechain[0].chain1.flip2[76] ;
 wire \thechain[0].chain1.flip2[77] ;
 wire \thechain[0].chain1.flip2[78] ;
 wire \thechain[0].chain1.flip2[79] ;
 wire \thechain[0].chain1.flip2[7] ;
 wire \thechain[0].chain1.flip2[8] ;
 wire \thechain[0].chain1.flip2[9] ;
 wire \thechain[1].chain1.dout ;
 wire \thechain[1].chain1.ff[0] ;
 wire \thechain[1].chain1.ff[10] ;
 wire \thechain[1].chain1.ff[11] ;
 wire \thechain[1].chain1.ff[12] ;
 wire \thechain[1].chain1.ff[13] ;
 wire \thechain[1].chain1.ff[14] ;
 wire \thechain[1].chain1.ff[15] ;
 wire \thechain[1].chain1.ff[16] ;
 wire \thechain[1].chain1.ff[17] ;
 wire \thechain[1].chain1.ff[18] ;
 wire \thechain[1].chain1.ff[19] ;
 wire \thechain[1].chain1.ff[1] ;
 wire \thechain[1].chain1.ff[20] ;
 wire \thechain[1].chain1.ff[21] ;
 wire \thechain[1].chain1.ff[22] ;
 wire \thechain[1].chain1.ff[23] ;
 wire \thechain[1].chain1.ff[24] ;
 wire \thechain[1].chain1.ff[25] ;
 wire \thechain[1].chain1.ff[26] ;
 wire \thechain[1].chain1.ff[27] ;
 wire \thechain[1].chain1.ff[28] ;
 wire \thechain[1].chain1.ff[29] ;
 wire \thechain[1].chain1.ff[2] ;
 wire \thechain[1].chain1.ff[30] ;
 wire \thechain[1].chain1.ff[31] ;
 wire \thechain[1].chain1.ff[32] ;
 wire \thechain[1].chain1.ff[33] ;
 wire \thechain[1].chain1.ff[34] ;
 wire \thechain[1].chain1.ff[35] ;
 wire \thechain[1].chain1.ff[36] ;
 wire \thechain[1].chain1.ff[37] ;
 wire \thechain[1].chain1.ff[38] ;
 wire \thechain[1].chain1.ff[39] ;
 wire \thechain[1].chain1.ff[3] ;
 wire \thechain[1].chain1.ff[40] ;
 wire \thechain[1].chain1.ff[41] ;
 wire \thechain[1].chain1.ff[42] ;
 wire \thechain[1].chain1.ff[43] ;
 wire \thechain[1].chain1.ff[44] ;
 wire \thechain[1].chain1.ff[45] ;
 wire \thechain[1].chain1.ff[46] ;
 wire \thechain[1].chain1.ff[47] ;
 wire \thechain[1].chain1.ff[48] ;
 wire \thechain[1].chain1.ff[49] ;
 wire \thechain[1].chain1.ff[4] ;
 wire \thechain[1].chain1.ff[50] ;
 wire \thechain[1].chain1.ff[51] ;
 wire \thechain[1].chain1.ff[52] ;
 wire \thechain[1].chain1.ff[53] ;
 wire \thechain[1].chain1.ff[54] ;
 wire \thechain[1].chain1.ff[55] ;
 wire \thechain[1].chain1.ff[56] ;
 wire \thechain[1].chain1.ff[57] ;
 wire \thechain[1].chain1.ff[58] ;
 wire \thechain[1].chain1.ff[59] ;
 wire \thechain[1].chain1.ff[5] ;
 wire \thechain[1].chain1.ff[60] ;
 wire \thechain[1].chain1.ff[61] ;
 wire \thechain[1].chain1.ff[62] ;
 wire \thechain[1].chain1.ff[63] ;
 wire \thechain[1].chain1.ff[64] ;
 wire \thechain[1].chain1.ff[65] ;
 wire \thechain[1].chain1.ff[66] ;
 wire \thechain[1].chain1.ff[67] ;
 wire \thechain[1].chain1.ff[68] ;
 wire \thechain[1].chain1.ff[69] ;
 wire \thechain[1].chain1.ff[6] ;
 wire \thechain[1].chain1.ff[70] ;
 wire \thechain[1].chain1.ff[71] ;
 wire \thechain[1].chain1.ff[72] ;
 wire \thechain[1].chain1.ff[73] ;
 wire \thechain[1].chain1.ff[74] ;
 wire \thechain[1].chain1.ff[75] ;
 wire \thechain[1].chain1.ff[76] ;
 wire \thechain[1].chain1.ff[77] ;
 wire \thechain[1].chain1.ff[78] ;
 wire \thechain[1].chain1.ff[7] ;
 wire \thechain[1].chain1.ff[8] ;
 wire \thechain[1].chain1.ff[9] ;
 wire \thechain[1].chain1.flip1[0] ;
 wire \thechain[1].chain1.flip1[10] ;
 wire \thechain[1].chain1.flip1[11] ;
 wire \thechain[1].chain1.flip1[12] ;
 wire \thechain[1].chain1.flip1[13] ;
 wire \thechain[1].chain1.flip1[14] ;
 wire \thechain[1].chain1.flip1[15] ;
 wire \thechain[1].chain1.flip1[16] ;
 wire \thechain[1].chain1.flip1[17] ;
 wire \thechain[1].chain1.flip1[18] ;
 wire \thechain[1].chain1.flip1[19] ;
 wire \thechain[1].chain1.flip1[1] ;
 wire \thechain[1].chain1.flip1[20] ;
 wire \thechain[1].chain1.flip1[21] ;
 wire \thechain[1].chain1.flip1[22] ;
 wire \thechain[1].chain1.flip1[23] ;
 wire \thechain[1].chain1.flip1[24] ;
 wire \thechain[1].chain1.flip1[25] ;
 wire \thechain[1].chain1.flip1[26] ;
 wire \thechain[1].chain1.flip1[27] ;
 wire \thechain[1].chain1.flip1[28] ;
 wire \thechain[1].chain1.flip1[29] ;
 wire \thechain[1].chain1.flip1[2] ;
 wire \thechain[1].chain1.flip1[30] ;
 wire \thechain[1].chain1.flip1[31] ;
 wire \thechain[1].chain1.flip1[32] ;
 wire \thechain[1].chain1.flip1[33] ;
 wire \thechain[1].chain1.flip1[34] ;
 wire \thechain[1].chain1.flip1[35] ;
 wire \thechain[1].chain1.flip1[36] ;
 wire \thechain[1].chain1.flip1[37] ;
 wire \thechain[1].chain1.flip1[38] ;
 wire \thechain[1].chain1.flip1[39] ;
 wire \thechain[1].chain1.flip1[3] ;
 wire \thechain[1].chain1.flip1[40] ;
 wire \thechain[1].chain1.flip1[41] ;
 wire \thechain[1].chain1.flip1[42] ;
 wire \thechain[1].chain1.flip1[43] ;
 wire \thechain[1].chain1.flip1[44] ;
 wire \thechain[1].chain1.flip1[45] ;
 wire \thechain[1].chain1.flip1[46] ;
 wire \thechain[1].chain1.flip1[47] ;
 wire \thechain[1].chain1.flip1[48] ;
 wire \thechain[1].chain1.flip1[49] ;
 wire \thechain[1].chain1.flip1[4] ;
 wire \thechain[1].chain1.flip1[50] ;
 wire \thechain[1].chain1.flip1[51] ;
 wire \thechain[1].chain1.flip1[52] ;
 wire \thechain[1].chain1.flip1[53] ;
 wire \thechain[1].chain1.flip1[54] ;
 wire \thechain[1].chain1.flip1[55] ;
 wire \thechain[1].chain1.flip1[56] ;
 wire \thechain[1].chain1.flip1[57] ;
 wire \thechain[1].chain1.flip1[58] ;
 wire \thechain[1].chain1.flip1[59] ;
 wire \thechain[1].chain1.flip1[5] ;
 wire \thechain[1].chain1.flip1[60] ;
 wire \thechain[1].chain1.flip1[61] ;
 wire \thechain[1].chain1.flip1[62] ;
 wire \thechain[1].chain1.flip1[63] ;
 wire \thechain[1].chain1.flip1[64] ;
 wire \thechain[1].chain1.flip1[65] ;
 wire \thechain[1].chain1.flip1[66] ;
 wire \thechain[1].chain1.flip1[67] ;
 wire \thechain[1].chain1.flip1[68] ;
 wire \thechain[1].chain1.flip1[69] ;
 wire \thechain[1].chain1.flip1[6] ;
 wire \thechain[1].chain1.flip1[70] ;
 wire \thechain[1].chain1.flip1[71] ;
 wire \thechain[1].chain1.flip1[72] ;
 wire \thechain[1].chain1.flip1[73] ;
 wire \thechain[1].chain1.flip1[74] ;
 wire \thechain[1].chain1.flip1[75] ;
 wire \thechain[1].chain1.flip1[76] ;
 wire \thechain[1].chain1.flip1[77] ;
 wire \thechain[1].chain1.flip1[78] ;
 wire \thechain[1].chain1.flip1[79] ;
 wire \thechain[1].chain1.flip1[7] ;
 wire \thechain[1].chain1.flip1[8] ;
 wire \thechain[1].chain1.flip1[9] ;
 wire \thechain[1].chain1.flip2[0] ;
 wire \thechain[1].chain1.flip2[10] ;
 wire \thechain[1].chain1.flip2[11] ;
 wire \thechain[1].chain1.flip2[12] ;
 wire \thechain[1].chain1.flip2[13] ;
 wire \thechain[1].chain1.flip2[14] ;
 wire \thechain[1].chain1.flip2[15] ;
 wire \thechain[1].chain1.flip2[16] ;
 wire \thechain[1].chain1.flip2[17] ;
 wire \thechain[1].chain1.flip2[18] ;
 wire \thechain[1].chain1.flip2[19] ;
 wire \thechain[1].chain1.flip2[1] ;
 wire \thechain[1].chain1.flip2[20] ;
 wire \thechain[1].chain1.flip2[21] ;
 wire \thechain[1].chain1.flip2[22] ;
 wire \thechain[1].chain1.flip2[23] ;
 wire \thechain[1].chain1.flip2[24] ;
 wire \thechain[1].chain1.flip2[25] ;
 wire \thechain[1].chain1.flip2[26] ;
 wire \thechain[1].chain1.flip2[27] ;
 wire \thechain[1].chain1.flip2[28] ;
 wire \thechain[1].chain1.flip2[29] ;
 wire \thechain[1].chain1.flip2[2] ;
 wire \thechain[1].chain1.flip2[30] ;
 wire \thechain[1].chain1.flip2[31] ;
 wire \thechain[1].chain1.flip2[32] ;
 wire \thechain[1].chain1.flip2[33] ;
 wire \thechain[1].chain1.flip2[34] ;
 wire \thechain[1].chain1.flip2[35] ;
 wire \thechain[1].chain1.flip2[36] ;
 wire \thechain[1].chain1.flip2[37] ;
 wire \thechain[1].chain1.flip2[38] ;
 wire \thechain[1].chain1.flip2[39] ;
 wire \thechain[1].chain1.flip2[3] ;
 wire \thechain[1].chain1.flip2[40] ;
 wire \thechain[1].chain1.flip2[41] ;
 wire \thechain[1].chain1.flip2[42] ;
 wire \thechain[1].chain1.flip2[43] ;
 wire \thechain[1].chain1.flip2[44] ;
 wire \thechain[1].chain1.flip2[45] ;
 wire \thechain[1].chain1.flip2[46] ;
 wire \thechain[1].chain1.flip2[47] ;
 wire \thechain[1].chain1.flip2[48] ;
 wire \thechain[1].chain1.flip2[49] ;
 wire \thechain[1].chain1.flip2[4] ;
 wire \thechain[1].chain1.flip2[50] ;
 wire \thechain[1].chain1.flip2[51] ;
 wire \thechain[1].chain1.flip2[52] ;
 wire \thechain[1].chain1.flip2[53] ;
 wire \thechain[1].chain1.flip2[54] ;
 wire \thechain[1].chain1.flip2[55] ;
 wire \thechain[1].chain1.flip2[56] ;
 wire \thechain[1].chain1.flip2[57] ;
 wire \thechain[1].chain1.flip2[58] ;
 wire \thechain[1].chain1.flip2[59] ;
 wire \thechain[1].chain1.flip2[5] ;
 wire \thechain[1].chain1.flip2[60] ;
 wire \thechain[1].chain1.flip2[61] ;
 wire \thechain[1].chain1.flip2[62] ;
 wire \thechain[1].chain1.flip2[63] ;
 wire \thechain[1].chain1.flip2[64] ;
 wire \thechain[1].chain1.flip2[65] ;
 wire \thechain[1].chain1.flip2[66] ;
 wire \thechain[1].chain1.flip2[67] ;
 wire \thechain[1].chain1.flip2[68] ;
 wire \thechain[1].chain1.flip2[69] ;
 wire \thechain[1].chain1.flip2[6] ;
 wire \thechain[1].chain1.flip2[70] ;
 wire \thechain[1].chain1.flip2[71] ;
 wire \thechain[1].chain1.flip2[72] ;
 wire \thechain[1].chain1.flip2[73] ;
 wire \thechain[1].chain1.flip2[74] ;
 wire \thechain[1].chain1.flip2[75] ;
 wire \thechain[1].chain1.flip2[76] ;
 wire \thechain[1].chain1.flip2[77] ;
 wire \thechain[1].chain1.flip2[78] ;
 wire \thechain[1].chain1.flip2[79] ;
 wire \thechain[1].chain1.flip2[7] ;
 wire \thechain[1].chain1.flip2[8] ;
 wire \thechain[1].chain1.flip2[9] ;
 wire \thechain[2].chain1.dout ;
 wire \thechain[2].chain1.ff[0] ;
 wire \thechain[2].chain1.ff[10] ;
 wire \thechain[2].chain1.ff[11] ;
 wire \thechain[2].chain1.ff[12] ;
 wire \thechain[2].chain1.ff[13] ;
 wire \thechain[2].chain1.ff[14] ;
 wire \thechain[2].chain1.ff[15] ;
 wire \thechain[2].chain1.ff[16] ;
 wire \thechain[2].chain1.ff[17] ;
 wire \thechain[2].chain1.ff[18] ;
 wire \thechain[2].chain1.ff[19] ;
 wire \thechain[2].chain1.ff[1] ;
 wire \thechain[2].chain1.ff[20] ;
 wire \thechain[2].chain1.ff[21] ;
 wire \thechain[2].chain1.ff[22] ;
 wire \thechain[2].chain1.ff[23] ;
 wire \thechain[2].chain1.ff[24] ;
 wire \thechain[2].chain1.ff[25] ;
 wire \thechain[2].chain1.ff[26] ;
 wire \thechain[2].chain1.ff[27] ;
 wire \thechain[2].chain1.ff[28] ;
 wire \thechain[2].chain1.ff[29] ;
 wire \thechain[2].chain1.ff[2] ;
 wire \thechain[2].chain1.ff[30] ;
 wire \thechain[2].chain1.ff[31] ;
 wire \thechain[2].chain1.ff[32] ;
 wire \thechain[2].chain1.ff[33] ;
 wire \thechain[2].chain1.ff[34] ;
 wire \thechain[2].chain1.ff[35] ;
 wire \thechain[2].chain1.ff[36] ;
 wire \thechain[2].chain1.ff[37] ;
 wire \thechain[2].chain1.ff[38] ;
 wire \thechain[2].chain1.ff[39] ;
 wire \thechain[2].chain1.ff[3] ;
 wire \thechain[2].chain1.ff[40] ;
 wire \thechain[2].chain1.ff[41] ;
 wire \thechain[2].chain1.ff[42] ;
 wire \thechain[2].chain1.ff[43] ;
 wire \thechain[2].chain1.ff[44] ;
 wire \thechain[2].chain1.ff[45] ;
 wire \thechain[2].chain1.ff[46] ;
 wire \thechain[2].chain1.ff[47] ;
 wire \thechain[2].chain1.ff[48] ;
 wire \thechain[2].chain1.ff[49] ;
 wire \thechain[2].chain1.ff[4] ;
 wire \thechain[2].chain1.ff[50] ;
 wire \thechain[2].chain1.ff[51] ;
 wire \thechain[2].chain1.ff[52] ;
 wire \thechain[2].chain1.ff[53] ;
 wire \thechain[2].chain1.ff[54] ;
 wire \thechain[2].chain1.ff[55] ;
 wire \thechain[2].chain1.ff[56] ;
 wire \thechain[2].chain1.ff[57] ;
 wire \thechain[2].chain1.ff[58] ;
 wire \thechain[2].chain1.ff[59] ;
 wire \thechain[2].chain1.ff[5] ;
 wire \thechain[2].chain1.ff[60] ;
 wire \thechain[2].chain1.ff[61] ;
 wire \thechain[2].chain1.ff[62] ;
 wire \thechain[2].chain1.ff[63] ;
 wire \thechain[2].chain1.ff[64] ;
 wire \thechain[2].chain1.ff[65] ;
 wire \thechain[2].chain1.ff[66] ;
 wire \thechain[2].chain1.ff[67] ;
 wire \thechain[2].chain1.ff[68] ;
 wire \thechain[2].chain1.ff[69] ;
 wire \thechain[2].chain1.ff[6] ;
 wire \thechain[2].chain1.ff[70] ;
 wire \thechain[2].chain1.ff[71] ;
 wire \thechain[2].chain1.ff[72] ;
 wire \thechain[2].chain1.ff[73] ;
 wire \thechain[2].chain1.ff[74] ;
 wire \thechain[2].chain1.ff[75] ;
 wire \thechain[2].chain1.ff[76] ;
 wire \thechain[2].chain1.ff[77] ;
 wire \thechain[2].chain1.ff[78] ;
 wire \thechain[2].chain1.ff[7] ;
 wire \thechain[2].chain1.ff[8] ;
 wire \thechain[2].chain1.ff[9] ;
 wire \thechain[2].chain1.flip1[0] ;
 wire \thechain[2].chain1.flip1[10] ;
 wire \thechain[2].chain1.flip1[11] ;
 wire \thechain[2].chain1.flip1[12] ;
 wire \thechain[2].chain1.flip1[13] ;
 wire \thechain[2].chain1.flip1[14] ;
 wire \thechain[2].chain1.flip1[15] ;
 wire \thechain[2].chain1.flip1[16] ;
 wire \thechain[2].chain1.flip1[17] ;
 wire \thechain[2].chain1.flip1[18] ;
 wire \thechain[2].chain1.flip1[19] ;
 wire \thechain[2].chain1.flip1[1] ;
 wire \thechain[2].chain1.flip1[20] ;
 wire \thechain[2].chain1.flip1[21] ;
 wire \thechain[2].chain1.flip1[22] ;
 wire \thechain[2].chain1.flip1[23] ;
 wire \thechain[2].chain1.flip1[24] ;
 wire \thechain[2].chain1.flip1[25] ;
 wire \thechain[2].chain1.flip1[26] ;
 wire \thechain[2].chain1.flip1[27] ;
 wire \thechain[2].chain1.flip1[28] ;
 wire \thechain[2].chain1.flip1[29] ;
 wire \thechain[2].chain1.flip1[2] ;
 wire \thechain[2].chain1.flip1[30] ;
 wire \thechain[2].chain1.flip1[31] ;
 wire \thechain[2].chain1.flip1[32] ;
 wire \thechain[2].chain1.flip1[33] ;
 wire \thechain[2].chain1.flip1[34] ;
 wire \thechain[2].chain1.flip1[35] ;
 wire \thechain[2].chain1.flip1[36] ;
 wire \thechain[2].chain1.flip1[37] ;
 wire \thechain[2].chain1.flip1[38] ;
 wire \thechain[2].chain1.flip1[39] ;
 wire \thechain[2].chain1.flip1[3] ;
 wire \thechain[2].chain1.flip1[40] ;
 wire \thechain[2].chain1.flip1[41] ;
 wire \thechain[2].chain1.flip1[42] ;
 wire \thechain[2].chain1.flip1[43] ;
 wire \thechain[2].chain1.flip1[44] ;
 wire \thechain[2].chain1.flip1[45] ;
 wire \thechain[2].chain1.flip1[46] ;
 wire \thechain[2].chain1.flip1[47] ;
 wire \thechain[2].chain1.flip1[48] ;
 wire \thechain[2].chain1.flip1[49] ;
 wire \thechain[2].chain1.flip1[4] ;
 wire \thechain[2].chain1.flip1[50] ;
 wire \thechain[2].chain1.flip1[51] ;
 wire \thechain[2].chain1.flip1[52] ;
 wire \thechain[2].chain1.flip1[53] ;
 wire \thechain[2].chain1.flip1[54] ;
 wire \thechain[2].chain1.flip1[55] ;
 wire \thechain[2].chain1.flip1[56] ;
 wire \thechain[2].chain1.flip1[57] ;
 wire \thechain[2].chain1.flip1[58] ;
 wire \thechain[2].chain1.flip1[59] ;
 wire \thechain[2].chain1.flip1[5] ;
 wire \thechain[2].chain1.flip1[60] ;
 wire \thechain[2].chain1.flip1[61] ;
 wire \thechain[2].chain1.flip1[62] ;
 wire \thechain[2].chain1.flip1[63] ;
 wire \thechain[2].chain1.flip1[64] ;
 wire \thechain[2].chain1.flip1[65] ;
 wire \thechain[2].chain1.flip1[66] ;
 wire \thechain[2].chain1.flip1[67] ;
 wire \thechain[2].chain1.flip1[68] ;
 wire \thechain[2].chain1.flip1[69] ;
 wire \thechain[2].chain1.flip1[6] ;
 wire \thechain[2].chain1.flip1[70] ;
 wire \thechain[2].chain1.flip1[71] ;
 wire \thechain[2].chain1.flip1[72] ;
 wire \thechain[2].chain1.flip1[73] ;
 wire \thechain[2].chain1.flip1[74] ;
 wire \thechain[2].chain1.flip1[75] ;
 wire \thechain[2].chain1.flip1[76] ;
 wire \thechain[2].chain1.flip1[77] ;
 wire \thechain[2].chain1.flip1[78] ;
 wire \thechain[2].chain1.flip1[79] ;
 wire \thechain[2].chain1.flip1[7] ;
 wire \thechain[2].chain1.flip1[8] ;
 wire \thechain[2].chain1.flip1[9] ;
 wire \thechain[2].chain1.flip2[0] ;
 wire \thechain[2].chain1.flip2[10] ;
 wire \thechain[2].chain1.flip2[11] ;
 wire \thechain[2].chain1.flip2[12] ;
 wire \thechain[2].chain1.flip2[13] ;
 wire \thechain[2].chain1.flip2[14] ;
 wire \thechain[2].chain1.flip2[15] ;
 wire \thechain[2].chain1.flip2[16] ;
 wire \thechain[2].chain1.flip2[17] ;
 wire \thechain[2].chain1.flip2[18] ;
 wire \thechain[2].chain1.flip2[19] ;
 wire \thechain[2].chain1.flip2[1] ;
 wire \thechain[2].chain1.flip2[20] ;
 wire \thechain[2].chain1.flip2[21] ;
 wire \thechain[2].chain1.flip2[22] ;
 wire \thechain[2].chain1.flip2[23] ;
 wire \thechain[2].chain1.flip2[24] ;
 wire \thechain[2].chain1.flip2[25] ;
 wire \thechain[2].chain1.flip2[26] ;
 wire \thechain[2].chain1.flip2[27] ;
 wire \thechain[2].chain1.flip2[28] ;
 wire \thechain[2].chain1.flip2[29] ;
 wire \thechain[2].chain1.flip2[2] ;
 wire \thechain[2].chain1.flip2[30] ;
 wire \thechain[2].chain1.flip2[31] ;
 wire \thechain[2].chain1.flip2[32] ;
 wire \thechain[2].chain1.flip2[33] ;
 wire \thechain[2].chain1.flip2[34] ;
 wire \thechain[2].chain1.flip2[35] ;
 wire \thechain[2].chain1.flip2[36] ;
 wire \thechain[2].chain1.flip2[37] ;
 wire \thechain[2].chain1.flip2[38] ;
 wire \thechain[2].chain1.flip2[39] ;
 wire \thechain[2].chain1.flip2[3] ;
 wire \thechain[2].chain1.flip2[40] ;
 wire \thechain[2].chain1.flip2[41] ;
 wire \thechain[2].chain1.flip2[42] ;
 wire \thechain[2].chain1.flip2[43] ;
 wire \thechain[2].chain1.flip2[44] ;
 wire \thechain[2].chain1.flip2[45] ;
 wire \thechain[2].chain1.flip2[46] ;
 wire \thechain[2].chain1.flip2[47] ;
 wire \thechain[2].chain1.flip2[48] ;
 wire \thechain[2].chain1.flip2[49] ;
 wire \thechain[2].chain1.flip2[4] ;
 wire \thechain[2].chain1.flip2[50] ;
 wire \thechain[2].chain1.flip2[51] ;
 wire \thechain[2].chain1.flip2[52] ;
 wire \thechain[2].chain1.flip2[53] ;
 wire \thechain[2].chain1.flip2[54] ;
 wire \thechain[2].chain1.flip2[55] ;
 wire \thechain[2].chain1.flip2[56] ;
 wire \thechain[2].chain1.flip2[57] ;
 wire \thechain[2].chain1.flip2[58] ;
 wire \thechain[2].chain1.flip2[59] ;
 wire \thechain[2].chain1.flip2[5] ;
 wire \thechain[2].chain1.flip2[60] ;
 wire \thechain[2].chain1.flip2[61] ;
 wire \thechain[2].chain1.flip2[62] ;
 wire \thechain[2].chain1.flip2[63] ;
 wire \thechain[2].chain1.flip2[64] ;
 wire \thechain[2].chain1.flip2[65] ;
 wire \thechain[2].chain1.flip2[66] ;
 wire \thechain[2].chain1.flip2[67] ;
 wire \thechain[2].chain1.flip2[68] ;
 wire \thechain[2].chain1.flip2[69] ;
 wire \thechain[2].chain1.flip2[6] ;
 wire \thechain[2].chain1.flip2[70] ;
 wire \thechain[2].chain1.flip2[71] ;
 wire \thechain[2].chain1.flip2[72] ;
 wire \thechain[2].chain1.flip2[73] ;
 wire \thechain[2].chain1.flip2[74] ;
 wire \thechain[2].chain1.flip2[75] ;
 wire \thechain[2].chain1.flip2[76] ;
 wire \thechain[2].chain1.flip2[77] ;
 wire \thechain[2].chain1.flip2[78] ;
 wire \thechain[2].chain1.flip2[79] ;
 wire \thechain[2].chain1.flip2[7] ;
 wire \thechain[2].chain1.flip2[8] ;
 wire \thechain[2].chain1.flip2[9] ;
 wire \thechain[3].chain1.dout ;
 wire \thechain[3].chain1.ff[0] ;
 wire \thechain[3].chain1.ff[10] ;
 wire \thechain[3].chain1.ff[11] ;
 wire \thechain[3].chain1.ff[12] ;
 wire \thechain[3].chain1.ff[13] ;
 wire \thechain[3].chain1.ff[14] ;
 wire \thechain[3].chain1.ff[15] ;
 wire \thechain[3].chain1.ff[16] ;
 wire \thechain[3].chain1.ff[17] ;
 wire \thechain[3].chain1.ff[18] ;
 wire \thechain[3].chain1.ff[19] ;
 wire \thechain[3].chain1.ff[1] ;
 wire \thechain[3].chain1.ff[20] ;
 wire \thechain[3].chain1.ff[21] ;
 wire \thechain[3].chain1.ff[22] ;
 wire \thechain[3].chain1.ff[23] ;
 wire \thechain[3].chain1.ff[24] ;
 wire \thechain[3].chain1.ff[25] ;
 wire \thechain[3].chain1.ff[26] ;
 wire \thechain[3].chain1.ff[27] ;
 wire \thechain[3].chain1.ff[28] ;
 wire \thechain[3].chain1.ff[29] ;
 wire \thechain[3].chain1.ff[2] ;
 wire \thechain[3].chain1.ff[30] ;
 wire \thechain[3].chain1.ff[31] ;
 wire \thechain[3].chain1.ff[32] ;
 wire \thechain[3].chain1.ff[33] ;
 wire \thechain[3].chain1.ff[34] ;
 wire \thechain[3].chain1.ff[35] ;
 wire \thechain[3].chain1.ff[36] ;
 wire \thechain[3].chain1.ff[37] ;
 wire \thechain[3].chain1.ff[38] ;
 wire \thechain[3].chain1.ff[39] ;
 wire \thechain[3].chain1.ff[3] ;
 wire \thechain[3].chain1.ff[40] ;
 wire \thechain[3].chain1.ff[41] ;
 wire \thechain[3].chain1.ff[42] ;
 wire \thechain[3].chain1.ff[43] ;
 wire \thechain[3].chain1.ff[44] ;
 wire \thechain[3].chain1.ff[45] ;
 wire \thechain[3].chain1.ff[46] ;
 wire \thechain[3].chain1.ff[47] ;
 wire \thechain[3].chain1.ff[48] ;
 wire \thechain[3].chain1.ff[49] ;
 wire \thechain[3].chain1.ff[4] ;
 wire \thechain[3].chain1.ff[50] ;
 wire \thechain[3].chain1.ff[51] ;
 wire \thechain[3].chain1.ff[52] ;
 wire \thechain[3].chain1.ff[53] ;
 wire \thechain[3].chain1.ff[54] ;
 wire \thechain[3].chain1.ff[55] ;
 wire \thechain[3].chain1.ff[56] ;
 wire \thechain[3].chain1.ff[57] ;
 wire \thechain[3].chain1.ff[58] ;
 wire \thechain[3].chain1.ff[59] ;
 wire \thechain[3].chain1.ff[5] ;
 wire \thechain[3].chain1.ff[60] ;
 wire \thechain[3].chain1.ff[61] ;
 wire \thechain[3].chain1.ff[62] ;
 wire \thechain[3].chain1.ff[63] ;
 wire \thechain[3].chain1.ff[64] ;
 wire \thechain[3].chain1.ff[65] ;
 wire \thechain[3].chain1.ff[66] ;
 wire \thechain[3].chain1.ff[67] ;
 wire \thechain[3].chain1.ff[68] ;
 wire \thechain[3].chain1.ff[69] ;
 wire \thechain[3].chain1.ff[6] ;
 wire \thechain[3].chain1.ff[70] ;
 wire \thechain[3].chain1.ff[71] ;
 wire \thechain[3].chain1.ff[72] ;
 wire \thechain[3].chain1.ff[73] ;
 wire \thechain[3].chain1.ff[74] ;
 wire \thechain[3].chain1.ff[75] ;
 wire \thechain[3].chain1.ff[76] ;
 wire \thechain[3].chain1.ff[77] ;
 wire \thechain[3].chain1.ff[78] ;
 wire \thechain[3].chain1.ff[7] ;
 wire \thechain[3].chain1.ff[8] ;
 wire \thechain[3].chain1.ff[9] ;
 wire \thechain[3].chain1.flip1[0] ;
 wire \thechain[3].chain1.flip1[10] ;
 wire \thechain[3].chain1.flip1[11] ;
 wire \thechain[3].chain1.flip1[12] ;
 wire \thechain[3].chain1.flip1[13] ;
 wire \thechain[3].chain1.flip1[14] ;
 wire \thechain[3].chain1.flip1[15] ;
 wire \thechain[3].chain1.flip1[16] ;
 wire \thechain[3].chain1.flip1[17] ;
 wire \thechain[3].chain1.flip1[18] ;
 wire \thechain[3].chain1.flip1[19] ;
 wire \thechain[3].chain1.flip1[1] ;
 wire \thechain[3].chain1.flip1[20] ;
 wire \thechain[3].chain1.flip1[21] ;
 wire \thechain[3].chain1.flip1[22] ;
 wire \thechain[3].chain1.flip1[23] ;
 wire \thechain[3].chain1.flip1[24] ;
 wire \thechain[3].chain1.flip1[25] ;
 wire \thechain[3].chain1.flip1[26] ;
 wire \thechain[3].chain1.flip1[27] ;
 wire \thechain[3].chain1.flip1[28] ;
 wire \thechain[3].chain1.flip1[29] ;
 wire \thechain[3].chain1.flip1[2] ;
 wire \thechain[3].chain1.flip1[30] ;
 wire \thechain[3].chain1.flip1[31] ;
 wire \thechain[3].chain1.flip1[32] ;
 wire \thechain[3].chain1.flip1[33] ;
 wire \thechain[3].chain1.flip1[34] ;
 wire \thechain[3].chain1.flip1[35] ;
 wire \thechain[3].chain1.flip1[36] ;
 wire \thechain[3].chain1.flip1[37] ;
 wire \thechain[3].chain1.flip1[38] ;
 wire \thechain[3].chain1.flip1[39] ;
 wire \thechain[3].chain1.flip1[3] ;
 wire \thechain[3].chain1.flip1[40] ;
 wire \thechain[3].chain1.flip1[41] ;
 wire \thechain[3].chain1.flip1[42] ;
 wire \thechain[3].chain1.flip1[43] ;
 wire \thechain[3].chain1.flip1[44] ;
 wire \thechain[3].chain1.flip1[45] ;
 wire \thechain[3].chain1.flip1[46] ;
 wire \thechain[3].chain1.flip1[47] ;
 wire \thechain[3].chain1.flip1[48] ;
 wire \thechain[3].chain1.flip1[49] ;
 wire \thechain[3].chain1.flip1[4] ;
 wire \thechain[3].chain1.flip1[50] ;
 wire \thechain[3].chain1.flip1[51] ;
 wire \thechain[3].chain1.flip1[52] ;
 wire \thechain[3].chain1.flip1[53] ;
 wire \thechain[3].chain1.flip1[54] ;
 wire \thechain[3].chain1.flip1[55] ;
 wire \thechain[3].chain1.flip1[56] ;
 wire \thechain[3].chain1.flip1[57] ;
 wire \thechain[3].chain1.flip1[58] ;
 wire \thechain[3].chain1.flip1[59] ;
 wire \thechain[3].chain1.flip1[5] ;
 wire \thechain[3].chain1.flip1[60] ;
 wire \thechain[3].chain1.flip1[61] ;
 wire \thechain[3].chain1.flip1[62] ;
 wire \thechain[3].chain1.flip1[63] ;
 wire \thechain[3].chain1.flip1[64] ;
 wire \thechain[3].chain1.flip1[65] ;
 wire \thechain[3].chain1.flip1[66] ;
 wire \thechain[3].chain1.flip1[67] ;
 wire \thechain[3].chain1.flip1[68] ;
 wire \thechain[3].chain1.flip1[69] ;
 wire \thechain[3].chain1.flip1[6] ;
 wire \thechain[3].chain1.flip1[70] ;
 wire \thechain[3].chain1.flip1[71] ;
 wire \thechain[3].chain1.flip1[72] ;
 wire \thechain[3].chain1.flip1[73] ;
 wire \thechain[3].chain1.flip1[74] ;
 wire \thechain[3].chain1.flip1[75] ;
 wire \thechain[3].chain1.flip1[76] ;
 wire \thechain[3].chain1.flip1[77] ;
 wire \thechain[3].chain1.flip1[78] ;
 wire \thechain[3].chain1.flip1[79] ;
 wire \thechain[3].chain1.flip1[7] ;
 wire \thechain[3].chain1.flip1[8] ;
 wire \thechain[3].chain1.flip1[9] ;
 wire \thechain[3].chain1.flip2[0] ;
 wire \thechain[3].chain1.flip2[10] ;
 wire \thechain[3].chain1.flip2[11] ;
 wire \thechain[3].chain1.flip2[12] ;
 wire \thechain[3].chain1.flip2[13] ;
 wire \thechain[3].chain1.flip2[14] ;
 wire \thechain[3].chain1.flip2[15] ;
 wire \thechain[3].chain1.flip2[16] ;
 wire \thechain[3].chain1.flip2[17] ;
 wire \thechain[3].chain1.flip2[18] ;
 wire \thechain[3].chain1.flip2[19] ;
 wire \thechain[3].chain1.flip2[1] ;
 wire \thechain[3].chain1.flip2[20] ;
 wire \thechain[3].chain1.flip2[21] ;
 wire \thechain[3].chain1.flip2[22] ;
 wire \thechain[3].chain1.flip2[23] ;
 wire \thechain[3].chain1.flip2[24] ;
 wire \thechain[3].chain1.flip2[25] ;
 wire \thechain[3].chain1.flip2[26] ;
 wire \thechain[3].chain1.flip2[27] ;
 wire \thechain[3].chain1.flip2[28] ;
 wire \thechain[3].chain1.flip2[29] ;
 wire \thechain[3].chain1.flip2[2] ;
 wire \thechain[3].chain1.flip2[30] ;
 wire \thechain[3].chain1.flip2[31] ;
 wire \thechain[3].chain1.flip2[32] ;
 wire \thechain[3].chain1.flip2[33] ;
 wire \thechain[3].chain1.flip2[34] ;
 wire \thechain[3].chain1.flip2[35] ;
 wire \thechain[3].chain1.flip2[36] ;
 wire \thechain[3].chain1.flip2[37] ;
 wire \thechain[3].chain1.flip2[38] ;
 wire \thechain[3].chain1.flip2[39] ;
 wire \thechain[3].chain1.flip2[3] ;
 wire \thechain[3].chain1.flip2[40] ;
 wire \thechain[3].chain1.flip2[41] ;
 wire \thechain[3].chain1.flip2[42] ;
 wire \thechain[3].chain1.flip2[43] ;
 wire \thechain[3].chain1.flip2[44] ;
 wire \thechain[3].chain1.flip2[45] ;
 wire \thechain[3].chain1.flip2[46] ;
 wire \thechain[3].chain1.flip2[47] ;
 wire \thechain[3].chain1.flip2[48] ;
 wire \thechain[3].chain1.flip2[49] ;
 wire \thechain[3].chain1.flip2[4] ;
 wire \thechain[3].chain1.flip2[50] ;
 wire \thechain[3].chain1.flip2[51] ;
 wire \thechain[3].chain1.flip2[52] ;
 wire \thechain[3].chain1.flip2[53] ;
 wire \thechain[3].chain1.flip2[54] ;
 wire \thechain[3].chain1.flip2[55] ;
 wire \thechain[3].chain1.flip2[56] ;
 wire \thechain[3].chain1.flip2[57] ;
 wire \thechain[3].chain1.flip2[58] ;
 wire \thechain[3].chain1.flip2[59] ;
 wire \thechain[3].chain1.flip2[5] ;
 wire \thechain[3].chain1.flip2[60] ;
 wire \thechain[3].chain1.flip2[61] ;
 wire \thechain[3].chain1.flip2[62] ;
 wire \thechain[3].chain1.flip2[63] ;
 wire \thechain[3].chain1.flip2[64] ;
 wire \thechain[3].chain1.flip2[65] ;
 wire \thechain[3].chain1.flip2[66] ;
 wire \thechain[3].chain1.flip2[67] ;
 wire \thechain[3].chain1.flip2[68] ;
 wire \thechain[3].chain1.flip2[69] ;
 wire \thechain[3].chain1.flip2[6] ;
 wire \thechain[3].chain1.flip2[70] ;
 wire \thechain[3].chain1.flip2[71] ;
 wire \thechain[3].chain1.flip2[72] ;
 wire \thechain[3].chain1.flip2[73] ;
 wire \thechain[3].chain1.flip2[74] ;
 wire \thechain[3].chain1.flip2[75] ;
 wire \thechain[3].chain1.flip2[76] ;
 wire \thechain[3].chain1.flip2[77] ;
 wire \thechain[3].chain1.flip2[78] ;
 wire \thechain[3].chain1.flip2[79] ;
 wire \thechain[3].chain1.flip2[7] ;
 wire \thechain[3].chain1.flip2[8] ;
 wire \thechain[3].chain1.flip2[9] ;
 wire \thechain[4].chain1.dout ;
 wire \thechain[4].chain1.ff[0] ;
 wire \thechain[4].chain1.ff[10] ;
 wire \thechain[4].chain1.ff[11] ;
 wire \thechain[4].chain1.ff[12] ;
 wire \thechain[4].chain1.ff[13] ;
 wire \thechain[4].chain1.ff[14] ;
 wire \thechain[4].chain1.ff[15] ;
 wire \thechain[4].chain1.ff[16] ;
 wire \thechain[4].chain1.ff[17] ;
 wire \thechain[4].chain1.ff[18] ;
 wire \thechain[4].chain1.ff[19] ;
 wire \thechain[4].chain1.ff[1] ;
 wire \thechain[4].chain1.ff[20] ;
 wire \thechain[4].chain1.ff[21] ;
 wire \thechain[4].chain1.ff[22] ;
 wire \thechain[4].chain1.ff[23] ;
 wire \thechain[4].chain1.ff[24] ;
 wire \thechain[4].chain1.ff[25] ;
 wire \thechain[4].chain1.ff[26] ;
 wire \thechain[4].chain1.ff[27] ;
 wire \thechain[4].chain1.ff[28] ;
 wire \thechain[4].chain1.ff[29] ;
 wire \thechain[4].chain1.ff[2] ;
 wire \thechain[4].chain1.ff[30] ;
 wire \thechain[4].chain1.ff[31] ;
 wire \thechain[4].chain1.ff[32] ;
 wire \thechain[4].chain1.ff[33] ;
 wire \thechain[4].chain1.ff[34] ;
 wire \thechain[4].chain1.ff[35] ;
 wire \thechain[4].chain1.ff[36] ;
 wire \thechain[4].chain1.ff[37] ;
 wire \thechain[4].chain1.ff[38] ;
 wire \thechain[4].chain1.ff[39] ;
 wire \thechain[4].chain1.ff[3] ;
 wire \thechain[4].chain1.ff[40] ;
 wire \thechain[4].chain1.ff[41] ;
 wire \thechain[4].chain1.ff[42] ;
 wire \thechain[4].chain1.ff[43] ;
 wire \thechain[4].chain1.ff[44] ;
 wire \thechain[4].chain1.ff[45] ;
 wire \thechain[4].chain1.ff[46] ;
 wire \thechain[4].chain1.ff[47] ;
 wire \thechain[4].chain1.ff[48] ;
 wire \thechain[4].chain1.ff[49] ;
 wire \thechain[4].chain1.ff[4] ;
 wire \thechain[4].chain1.ff[50] ;
 wire \thechain[4].chain1.ff[51] ;
 wire \thechain[4].chain1.ff[52] ;
 wire \thechain[4].chain1.ff[53] ;
 wire \thechain[4].chain1.ff[54] ;
 wire \thechain[4].chain1.ff[55] ;
 wire \thechain[4].chain1.ff[56] ;
 wire \thechain[4].chain1.ff[57] ;
 wire \thechain[4].chain1.ff[58] ;
 wire \thechain[4].chain1.ff[59] ;
 wire \thechain[4].chain1.ff[5] ;
 wire \thechain[4].chain1.ff[60] ;
 wire \thechain[4].chain1.ff[61] ;
 wire \thechain[4].chain1.ff[62] ;
 wire \thechain[4].chain1.ff[63] ;
 wire \thechain[4].chain1.ff[64] ;
 wire \thechain[4].chain1.ff[65] ;
 wire \thechain[4].chain1.ff[66] ;
 wire \thechain[4].chain1.ff[67] ;
 wire \thechain[4].chain1.ff[68] ;
 wire \thechain[4].chain1.ff[69] ;
 wire \thechain[4].chain1.ff[6] ;
 wire \thechain[4].chain1.ff[70] ;
 wire \thechain[4].chain1.ff[71] ;
 wire \thechain[4].chain1.ff[72] ;
 wire \thechain[4].chain1.ff[73] ;
 wire \thechain[4].chain1.ff[74] ;
 wire \thechain[4].chain1.ff[75] ;
 wire \thechain[4].chain1.ff[76] ;
 wire \thechain[4].chain1.ff[77] ;
 wire \thechain[4].chain1.ff[78] ;
 wire \thechain[4].chain1.ff[7] ;
 wire \thechain[4].chain1.ff[8] ;
 wire \thechain[4].chain1.ff[9] ;
 wire \thechain[4].chain1.flip1[0] ;
 wire \thechain[4].chain1.flip1[10] ;
 wire \thechain[4].chain1.flip1[11] ;
 wire \thechain[4].chain1.flip1[12] ;
 wire \thechain[4].chain1.flip1[13] ;
 wire \thechain[4].chain1.flip1[14] ;
 wire \thechain[4].chain1.flip1[15] ;
 wire \thechain[4].chain1.flip1[16] ;
 wire \thechain[4].chain1.flip1[17] ;
 wire \thechain[4].chain1.flip1[18] ;
 wire \thechain[4].chain1.flip1[19] ;
 wire \thechain[4].chain1.flip1[1] ;
 wire \thechain[4].chain1.flip1[20] ;
 wire \thechain[4].chain1.flip1[21] ;
 wire \thechain[4].chain1.flip1[22] ;
 wire \thechain[4].chain1.flip1[23] ;
 wire \thechain[4].chain1.flip1[24] ;
 wire \thechain[4].chain1.flip1[25] ;
 wire \thechain[4].chain1.flip1[26] ;
 wire \thechain[4].chain1.flip1[27] ;
 wire \thechain[4].chain1.flip1[28] ;
 wire \thechain[4].chain1.flip1[29] ;
 wire \thechain[4].chain1.flip1[2] ;
 wire \thechain[4].chain1.flip1[30] ;
 wire \thechain[4].chain1.flip1[31] ;
 wire \thechain[4].chain1.flip1[32] ;
 wire \thechain[4].chain1.flip1[33] ;
 wire \thechain[4].chain1.flip1[34] ;
 wire \thechain[4].chain1.flip1[35] ;
 wire \thechain[4].chain1.flip1[36] ;
 wire \thechain[4].chain1.flip1[37] ;
 wire \thechain[4].chain1.flip1[38] ;
 wire \thechain[4].chain1.flip1[39] ;
 wire \thechain[4].chain1.flip1[3] ;
 wire \thechain[4].chain1.flip1[40] ;
 wire \thechain[4].chain1.flip1[41] ;
 wire \thechain[4].chain1.flip1[42] ;
 wire \thechain[4].chain1.flip1[43] ;
 wire \thechain[4].chain1.flip1[44] ;
 wire \thechain[4].chain1.flip1[45] ;
 wire \thechain[4].chain1.flip1[46] ;
 wire \thechain[4].chain1.flip1[47] ;
 wire \thechain[4].chain1.flip1[48] ;
 wire \thechain[4].chain1.flip1[49] ;
 wire \thechain[4].chain1.flip1[4] ;
 wire \thechain[4].chain1.flip1[50] ;
 wire \thechain[4].chain1.flip1[51] ;
 wire \thechain[4].chain1.flip1[52] ;
 wire \thechain[4].chain1.flip1[53] ;
 wire \thechain[4].chain1.flip1[54] ;
 wire \thechain[4].chain1.flip1[55] ;
 wire \thechain[4].chain1.flip1[56] ;
 wire \thechain[4].chain1.flip1[57] ;
 wire \thechain[4].chain1.flip1[58] ;
 wire \thechain[4].chain1.flip1[59] ;
 wire \thechain[4].chain1.flip1[5] ;
 wire \thechain[4].chain1.flip1[60] ;
 wire \thechain[4].chain1.flip1[61] ;
 wire \thechain[4].chain1.flip1[62] ;
 wire \thechain[4].chain1.flip1[63] ;
 wire \thechain[4].chain1.flip1[64] ;
 wire \thechain[4].chain1.flip1[65] ;
 wire \thechain[4].chain1.flip1[66] ;
 wire \thechain[4].chain1.flip1[67] ;
 wire \thechain[4].chain1.flip1[68] ;
 wire \thechain[4].chain1.flip1[69] ;
 wire \thechain[4].chain1.flip1[6] ;
 wire \thechain[4].chain1.flip1[70] ;
 wire \thechain[4].chain1.flip1[71] ;
 wire \thechain[4].chain1.flip1[72] ;
 wire \thechain[4].chain1.flip1[73] ;
 wire \thechain[4].chain1.flip1[74] ;
 wire \thechain[4].chain1.flip1[75] ;
 wire \thechain[4].chain1.flip1[76] ;
 wire \thechain[4].chain1.flip1[77] ;
 wire \thechain[4].chain1.flip1[78] ;
 wire \thechain[4].chain1.flip1[79] ;
 wire \thechain[4].chain1.flip1[7] ;
 wire \thechain[4].chain1.flip1[8] ;
 wire \thechain[4].chain1.flip1[9] ;
 wire \thechain[4].chain1.flip2[0] ;
 wire \thechain[4].chain1.flip2[10] ;
 wire \thechain[4].chain1.flip2[11] ;
 wire \thechain[4].chain1.flip2[12] ;
 wire \thechain[4].chain1.flip2[13] ;
 wire \thechain[4].chain1.flip2[14] ;
 wire \thechain[4].chain1.flip2[15] ;
 wire \thechain[4].chain1.flip2[16] ;
 wire \thechain[4].chain1.flip2[17] ;
 wire \thechain[4].chain1.flip2[18] ;
 wire \thechain[4].chain1.flip2[19] ;
 wire \thechain[4].chain1.flip2[1] ;
 wire \thechain[4].chain1.flip2[20] ;
 wire \thechain[4].chain1.flip2[21] ;
 wire \thechain[4].chain1.flip2[22] ;
 wire \thechain[4].chain1.flip2[23] ;
 wire \thechain[4].chain1.flip2[24] ;
 wire \thechain[4].chain1.flip2[25] ;
 wire \thechain[4].chain1.flip2[26] ;
 wire \thechain[4].chain1.flip2[27] ;
 wire \thechain[4].chain1.flip2[28] ;
 wire \thechain[4].chain1.flip2[29] ;
 wire \thechain[4].chain1.flip2[2] ;
 wire \thechain[4].chain1.flip2[30] ;
 wire \thechain[4].chain1.flip2[31] ;
 wire \thechain[4].chain1.flip2[32] ;
 wire \thechain[4].chain1.flip2[33] ;
 wire \thechain[4].chain1.flip2[34] ;
 wire \thechain[4].chain1.flip2[35] ;
 wire \thechain[4].chain1.flip2[36] ;
 wire \thechain[4].chain1.flip2[37] ;
 wire \thechain[4].chain1.flip2[38] ;
 wire \thechain[4].chain1.flip2[39] ;
 wire \thechain[4].chain1.flip2[3] ;
 wire \thechain[4].chain1.flip2[40] ;
 wire \thechain[4].chain1.flip2[41] ;
 wire \thechain[4].chain1.flip2[42] ;
 wire \thechain[4].chain1.flip2[43] ;
 wire \thechain[4].chain1.flip2[44] ;
 wire \thechain[4].chain1.flip2[45] ;
 wire \thechain[4].chain1.flip2[46] ;
 wire \thechain[4].chain1.flip2[47] ;
 wire \thechain[4].chain1.flip2[48] ;
 wire \thechain[4].chain1.flip2[49] ;
 wire \thechain[4].chain1.flip2[4] ;
 wire \thechain[4].chain1.flip2[50] ;
 wire \thechain[4].chain1.flip2[51] ;
 wire \thechain[4].chain1.flip2[52] ;
 wire \thechain[4].chain1.flip2[53] ;
 wire \thechain[4].chain1.flip2[54] ;
 wire \thechain[4].chain1.flip2[55] ;
 wire \thechain[4].chain1.flip2[56] ;
 wire \thechain[4].chain1.flip2[57] ;
 wire \thechain[4].chain1.flip2[58] ;
 wire \thechain[4].chain1.flip2[59] ;
 wire \thechain[4].chain1.flip2[5] ;
 wire \thechain[4].chain1.flip2[60] ;
 wire \thechain[4].chain1.flip2[61] ;
 wire \thechain[4].chain1.flip2[62] ;
 wire \thechain[4].chain1.flip2[63] ;
 wire \thechain[4].chain1.flip2[64] ;
 wire \thechain[4].chain1.flip2[65] ;
 wire \thechain[4].chain1.flip2[66] ;
 wire \thechain[4].chain1.flip2[67] ;
 wire \thechain[4].chain1.flip2[68] ;
 wire \thechain[4].chain1.flip2[69] ;
 wire \thechain[4].chain1.flip2[6] ;
 wire \thechain[4].chain1.flip2[70] ;
 wire \thechain[4].chain1.flip2[71] ;
 wire \thechain[4].chain1.flip2[72] ;
 wire \thechain[4].chain1.flip2[73] ;
 wire \thechain[4].chain1.flip2[74] ;
 wire \thechain[4].chain1.flip2[75] ;
 wire \thechain[4].chain1.flip2[76] ;
 wire \thechain[4].chain1.flip2[77] ;
 wire \thechain[4].chain1.flip2[78] ;
 wire \thechain[4].chain1.flip2[79] ;
 wire \thechain[4].chain1.flip2[7] ;
 wire \thechain[4].chain1.flip2[8] ;
 wire \thechain[4].chain1.flip2[9] ;
 wire \thechain[5].chain1.dout ;
 wire \thechain[5].chain1.ff[0] ;
 wire \thechain[5].chain1.ff[10] ;
 wire \thechain[5].chain1.ff[11] ;
 wire \thechain[5].chain1.ff[12] ;
 wire \thechain[5].chain1.ff[13] ;
 wire \thechain[5].chain1.ff[14] ;
 wire \thechain[5].chain1.ff[15] ;
 wire \thechain[5].chain1.ff[16] ;
 wire \thechain[5].chain1.ff[17] ;
 wire \thechain[5].chain1.ff[18] ;
 wire \thechain[5].chain1.ff[19] ;
 wire \thechain[5].chain1.ff[1] ;
 wire \thechain[5].chain1.ff[20] ;
 wire \thechain[5].chain1.ff[21] ;
 wire \thechain[5].chain1.ff[22] ;
 wire \thechain[5].chain1.ff[23] ;
 wire \thechain[5].chain1.ff[24] ;
 wire \thechain[5].chain1.ff[25] ;
 wire \thechain[5].chain1.ff[26] ;
 wire \thechain[5].chain1.ff[27] ;
 wire \thechain[5].chain1.ff[28] ;
 wire \thechain[5].chain1.ff[29] ;
 wire \thechain[5].chain1.ff[2] ;
 wire \thechain[5].chain1.ff[30] ;
 wire \thechain[5].chain1.ff[31] ;
 wire \thechain[5].chain1.ff[32] ;
 wire \thechain[5].chain1.ff[33] ;
 wire \thechain[5].chain1.ff[34] ;
 wire \thechain[5].chain1.ff[35] ;
 wire \thechain[5].chain1.ff[36] ;
 wire \thechain[5].chain1.ff[37] ;
 wire \thechain[5].chain1.ff[38] ;
 wire \thechain[5].chain1.ff[39] ;
 wire \thechain[5].chain1.ff[3] ;
 wire \thechain[5].chain1.ff[40] ;
 wire \thechain[5].chain1.ff[41] ;
 wire \thechain[5].chain1.ff[42] ;
 wire \thechain[5].chain1.ff[43] ;
 wire \thechain[5].chain1.ff[44] ;
 wire \thechain[5].chain1.ff[45] ;
 wire \thechain[5].chain1.ff[46] ;
 wire \thechain[5].chain1.ff[47] ;
 wire \thechain[5].chain1.ff[48] ;
 wire \thechain[5].chain1.ff[49] ;
 wire \thechain[5].chain1.ff[4] ;
 wire \thechain[5].chain1.ff[50] ;
 wire \thechain[5].chain1.ff[51] ;
 wire \thechain[5].chain1.ff[52] ;
 wire \thechain[5].chain1.ff[53] ;
 wire \thechain[5].chain1.ff[54] ;
 wire \thechain[5].chain1.ff[55] ;
 wire \thechain[5].chain1.ff[56] ;
 wire \thechain[5].chain1.ff[57] ;
 wire \thechain[5].chain1.ff[58] ;
 wire \thechain[5].chain1.ff[59] ;
 wire \thechain[5].chain1.ff[5] ;
 wire \thechain[5].chain1.ff[60] ;
 wire \thechain[5].chain1.ff[61] ;
 wire \thechain[5].chain1.ff[62] ;
 wire \thechain[5].chain1.ff[63] ;
 wire \thechain[5].chain1.ff[64] ;
 wire \thechain[5].chain1.ff[65] ;
 wire \thechain[5].chain1.ff[66] ;
 wire \thechain[5].chain1.ff[67] ;
 wire \thechain[5].chain1.ff[68] ;
 wire \thechain[5].chain1.ff[69] ;
 wire \thechain[5].chain1.ff[6] ;
 wire \thechain[5].chain1.ff[70] ;
 wire \thechain[5].chain1.ff[71] ;
 wire \thechain[5].chain1.ff[72] ;
 wire \thechain[5].chain1.ff[73] ;
 wire \thechain[5].chain1.ff[74] ;
 wire \thechain[5].chain1.ff[75] ;
 wire \thechain[5].chain1.ff[76] ;
 wire \thechain[5].chain1.ff[77] ;
 wire \thechain[5].chain1.ff[78] ;
 wire \thechain[5].chain1.ff[7] ;
 wire \thechain[5].chain1.ff[8] ;
 wire \thechain[5].chain1.ff[9] ;
 wire \thechain[5].chain1.flip1[0] ;
 wire \thechain[5].chain1.flip1[10] ;
 wire \thechain[5].chain1.flip1[11] ;
 wire \thechain[5].chain1.flip1[12] ;
 wire \thechain[5].chain1.flip1[13] ;
 wire \thechain[5].chain1.flip1[14] ;
 wire \thechain[5].chain1.flip1[15] ;
 wire \thechain[5].chain1.flip1[16] ;
 wire \thechain[5].chain1.flip1[17] ;
 wire \thechain[5].chain1.flip1[18] ;
 wire \thechain[5].chain1.flip1[19] ;
 wire \thechain[5].chain1.flip1[1] ;
 wire \thechain[5].chain1.flip1[20] ;
 wire \thechain[5].chain1.flip1[21] ;
 wire \thechain[5].chain1.flip1[22] ;
 wire \thechain[5].chain1.flip1[23] ;
 wire \thechain[5].chain1.flip1[24] ;
 wire \thechain[5].chain1.flip1[25] ;
 wire \thechain[5].chain1.flip1[26] ;
 wire \thechain[5].chain1.flip1[27] ;
 wire \thechain[5].chain1.flip1[28] ;
 wire \thechain[5].chain1.flip1[29] ;
 wire \thechain[5].chain1.flip1[2] ;
 wire \thechain[5].chain1.flip1[30] ;
 wire \thechain[5].chain1.flip1[31] ;
 wire \thechain[5].chain1.flip1[32] ;
 wire \thechain[5].chain1.flip1[33] ;
 wire \thechain[5].chain1.flip1[34] ;
 wire \thechain[5].chain1.flip1[35] ;
 wire \thechain[5].chain1.flip1[36] ;
 wire \thechain[5].chain1.flip1[37] ;
 wire \thechain[5].chain1.flip1[38] ;
 wire \thechain[5].chain1.flip1[39] ;
 wire \thechain[5].chain1.flip1[3] ;
 wire \thechain[5].chain1.flip1[40] ;
 wire \thechain[5].chain1.flip1[41] ;
 wire \thechain[5].chain1.flip1[42] ;
 wire \thechain[5].chain1.flip1[43] ;
 wire \thechain[5].chain1.flip1[44] ;
 wire \thechain[5].chain1.flip1[45] ;
 wire \thechain[5].chain1.flip1[46] ;
 wire \thechain[5].chain1.flip1[47] ;
 wire \thechain[5].chain1.flip1[48] ;
 wire \thechain[5].chain1.flip1[49] ;
 wire \thechain[5].chain1.flip1[4] ;
 wire \thechain[5].chain1.flip1[50] ;
 wire \thechain[5].chain1.flip1[51] ;
 wire \thechain[5].chain1.flip1[52] ;
 wire \thechain[5].chain1.flip1[53] ;
 wire \thechain[5].chain1.flip1[54] ;
 wire \thechain[5].chain1.flip1[55] ;
 wire \thechain[5].chain1.flip1[56] ;
 wire \thechain[5].chain1.flip1[57] ;
 wire \thechain[5].chain1.flip1[58] ;
 wire \thechain[5].chain1.flip1[59] ;
 wire \thechain[5].chain1.flip1[5] ;
 wire \thechain[5].chain1.flip1[60] ;
 wire \thechain[5].chain1.flip1[61] ;
 wire \thechain[5].chain1.flip1[62] ;
 wire \thechain[5].chain1.flip1[63] ;
 wire \thechain[5].chain1.flip1[64] ;
 wire \thechain[5].chain1.flip1[65] ;
 wire \thechain[5].chain1.flip1[66] ;
 wire \thechain[5].chain1.flip1[67] ;
 wire \thechain[5].chain1.flip1[68] ;
 wire \thechain[5].chain1.flip1[69] ;
 wire \thechain[5].chain1.flip1[6] ;
 wire \thechain[5].chain1.flip1[70] ;
 wire \thechain[5].chain1.flip1[71] ;
 wire \thechain[5].chain1.flip1[72] ;
 wire \thechain[5].chain1.flip1[73] ;
 wire \thechain[5].chain1.flip1[74] ;
 wire \thechain[5].chain1.flip1[75] ;
 wire \thechain[5].chain1.flip1[76] ;
 wire \thechain[5].chain1.flip1[77] ;
 wire \thechain[5].chain1.flip1[78] ;
 wire \thechain[5].chain1.flip1[79] ;
 wire \thechain[5].chain1.flip1[7] ;
 wire \thechain[5].chain1.flip1[8] ;
 wire \thechain[5].chain1.flip1[9] ;
 wire \thechain[5].chain1.flip2[0] ;
 wire \thechain[5].chain1.flip2[10] ;
 wire \thechain[5].chain1.flip2[11] ;
 wire \thechain[5].chain1.flip2[12] ;
 wire \thechain[5].chain1.flip2[13] ;
 wire \thechain[5].chain1.flip2[14] ;
 wire \thechain[5].chain1.flip2[15] ;
 wire \thechain[5].chain1.flip2[16] ;
 wire \thechain[5].chain1.flip2[17] ;
 wire \thechain[5].chain1.flip2[18] ;
 wire \thechain[5].chain1.flip2[19] ;
 wire \thechain[5].chain1.flip2[1] ;
 wire \thechain[5].chain1.flip2[20] ;
 wire \thechain[5].chain1.flip2[21] ;
 wire \thechain[5].chain1.flip2[22] ;
 wire \thechain[5].chain1.flip2[23] ;
 wire \thechain[5].chain1.flip2[24] ;
 wire \thechain[5].chain1.flip2[25] ;
 wire \thechain[5].chain1.flip2[26] ;
 wire \thechain[5].chain1.flip2[27] ;
 wire \thechain[5].chain1.flip2[28] ;
 wire \thechain[5].chain1.flip2[29] ;
 wire \thechain[5].chain1.flip2[2] ;
 wire \thechain[5].chain1.flip2[30] ;
 wire \thechain[5].chain1.flip2[31] ;
 wire \thechain[5].chain1.flip2[32] ;
 wire \thechain[5].chain1.flip2[33] ;
 wire \thechain[5].chain1.flip2[34] ;
 wire \thechain[5].chain1.flip2[35] ;
 wire \thechain[5].chain1.flip2[36] ;
 wire \thechain[5].chain1.flip2[37] ;
 wire \thechain[5].chain1.flip2[38] ;
 wire \thechain[5].chain1.flip2[39] ;
 wire \thechain[5].chain1.flip2[3] ;
 wire \thechain[5].chain1.flip2[40] ;
 wire \thechain[5].chain1.flip2[41] ;
 wire \thechain[5].chain1.flip2[42] ;
 wire \thechain[5].chain1.flip2[43] ;
 wire \thechain[5].chain1.flip2[44] ;
 wire \thechain[5].chain1.flip2[45] ;
 wire \thechain[5].chain1.flip2[46] ;
 wire \thechain[5].chain1.flip2[47] ;
 wire \thechain[5].chain1.flip2[48] ;
 wire \thechain[5].chain1.flip2[49] ;
 wire \thechain[5].chain1.flip2[4] ;
 wire \thechain[5].chain1.flip2[50] ;
 wire \thechain[5].chain1.flip2[51] ;
 wire \thechain[5].chain1.flip2[52] ;
 wire \thechain[5].chain1.flip2[53] ;
 wire \thechain[5].chain1.flip2[54] ;
 wire \thechain[5].chain1.flip2[55] ;
 wire \thechain[5].chain1.flip2[56] ;
 wire \thechain[5].chain1.flip2[57] ;
 wire \thechain[5].chain1.flip2[58] ;
 wire \thechain[5].chain1.flip2[59] ;
 wire \thechain[5].chain1.flip2[5] ;
 wire \thechain[5].chain1.flip2[60] ;
 wire \thechain[5].chain1.flip2[61] ;
 wire \thechain[5].chain1.flip2[62] ;
 wire \thechain[5].chain1.flip2[63] ;
 wire \thechain[5].chain1.flip2[64] ;
 wire \thechain[5].chain1.flip2[65] ;
 wire \thechain[5].chain1.flip2[66] ;
 wire \thechain[5].chain1.flip2[67] ;
 wire \thechain[5].chain1.flip2[68] ;
 wire \thechain[5].chain1.flip2[69] ;
 wire \thechain[5].chain1.flip2[6] ;
 wire \thechain[5].chain1.flip2[70] ;
 wire \thechain[5].chain1.flip2[71] ;
 wire \thechain[5].chain1.flip2[72] ;
 wire \thechain[5].chain1.flip2[73] ;
 wire \thechain[5].chain1.flip2[74] ;
 wire \thechain[5].chain1.flip2[75] ;
 wire \thechain[5].chain1.flip2[76] ;
 wire \thechain[5].chain1.flip2[77] ;
 wire \thechain[5].chain1.flip2[78] ;
 wire \thechain[5].chain1.flip2[79] ;
 wire \thechain[5].chain1.flip2[7] ;
 wire \thechain[5].chain1.flip2[8] ;
 wire \thechain[5].chain1.flip2[9] ;
 wire \thechain[6].chain1.dout ;
 wire \thechain[6].chain1.ff[0] ;
 wire \thechain[6].chain1.ff[10] ;
 wire \thechain[6].chain1.ff[11] ;
 wire \thechain[6].chain1.ff[12] ;
 wire \thechain[6].chain1.ff[13] ;
 wire \thechain[6].chain1.ff[14] ;
 wire \thechain[6].chain1.ff[15] ;
 wire \thechain[6].chain1.ff[16] ;
 wire \thechain[6].chain1.ff[17] ;
 wire \thechain[6].chain1.ff[18] ;
 wire \thechain[6].chain1.ff[19] ;
 wire \thechain[6].chain1.ff[1] ;
 wire \thechain[6].chain1.ff[20] ;
 wire \thechain[6].chain1.ff[21] ;
 wire \thechain[6].chain1.ff[22] ;
 wire \thechain[6].chain1.ff[23] ;
 wire \thechain[6].chain1.ff[24] ;
 wire \thechain[6].chain1.ff[25] ;
 wire \thechain[6].chain1.ff[26] ;
 wire \thechain[6].chain1.ff[27] ;
 wire \thechain[6].chain1.ff[28] ;
 wire \thechain[6].chain1.ff[29] ;
 wire \thechain[6].chain1.ff[2] ;
 wire \thechain[6].chain1.ff[30] ;
 wire \thechain[6].chain1.ff[31] ;
 wire \thechain[6].chain1.ff[32] ;
 wire \thechain[6].chain1.ff[33] ;
 wire \thechain[6].chain1.ff[34] ;
 wire \thechain[6].chain1.ff[35] ;
 wire \thechain[6].chain1.ff[36] ;
 wire \thechain[6].chain1.ff[37] ;
 wire \thechain[6].chain1.ff[38] ;
 wire \thechain[6].chain1.ff[39] ;
 wire \thechain[6].chain1.ff[3] ;
 wire \thechain[6].chain1.ff[40] ;
 wire \thechain[6].chain1.ff[41] ;
 wire \thechain[6].chain1.ff[42] ;
 wire \thechain[6].chain1.ff[43] ;
 wire \thechain[6].chain1.ff[44] ;
 wire \thechain[6].chain1.ff[45] ;
 wire \thechain[6].chain1.ff[46] ;
 wire \thechain[6].chain1.ff[47] ;
 wire \thechain[6].chain1.ff[48] ;
 wire \thechain[6].chain1.ff[49] ;
 wire \thechain[6].chain1.ff[4] ;
 wire \thechain[6].chain1.ff[50] ;
 wire \thechain[6].chain1.ff[51] ;
 wire \thechain[6].chain1.ff[52] ;
 wire \thechain[6].chain1.ff[53] ;
 wire \thechain[6].chain1.ff[54] ;
 wire \thechain[6].chain1.ff[55] ;
 wire \thechain[6].chain1.ff[56] ;
 wire \thechain[6].chain1.ff[57] ;
 wire \thechain[6].chain1.ff[58] ;
 wire \thechain[6].chain1.ff[59] ;
 wire \thechain[6].chain1.ff[5] ;
 wire \thechain[6].chain1.ff[60] ;
 wire \thechain[6].chain1.ff[61] ;
 wire \thechain[6].chain1.ff[62] ;
 wire \thechain[6].chain1.ff[63] ;
 wire \thechain[6].chain1.ff[64] ;
 wire \thechain[6].chain1.ff[65] ;
 wire \thechain[6].chain1.ff[66] ;
 wire \thechain[6].chain1.ff[67] ;
 wire \thechain[6].chain1.ff[68] ;
 wire \thechain[6].chain1.ff[69] ;
 wire \thechain[6].chain1.ff[6] ;
 wire \thechain[6].chain1.ff[70] ;
 wire \thechain[6].chain1.ff[71] ;
 wire \thechain[6].chain1.ff[72] ;
 wire \thechain[6].chain1.ff[73] ;
 wire \thechain[6].chain1.ff[74] ;
 wire \thechain[6].chain1.ff[75] ;
 wire \thechain[6].chain1.ff[76] ;
 wire \thechain[6].chain1.ff[77] ;
 wire \thechain[6].chain1.ff[78] ;
 wire \thechain[6].chain1.ff[7] ;
 wire \thechain[6].chain1.ff[8] ;
 wire \thechain[6].chain1.ff[9] ;
 wire \thechain[6].chain1.flip1[0] ;
 wire \thechain[6].chain1.flip1[10] ;
 wire \thechain[6].chain1.flip1[11] ;
 wire \thechain[6].chain1.flip1[12] ;
 wire \thechain[6].chain1.flip1[13] ;
 wire \thechain[6].chain1.flip1[14] ;
 wire \thechain[6].chain1.flip1[15] ;
 wire \thechain[6].chain1.flip1[16] ;
 wire \thechain[6].chain1.flip1[17] ;
 wire \thechain[6].chain1.flip1[18] ;
 wire \thechain[6].chain1.flip1[19] ;
 wire \thechain[6].chain1.flip1[1] ;
 wire \thechain[6].chain1.flip1[20] ;
 wire \thechain[6].chain1.flip1[21] ;
 wire \thechain[6].chain1.flip1[22] ;
 wire \thechain[6].chain1.flip1[23] ;
 wire \thechain[6].chain1.flip1[24] ;
 wire \thechain[6].chain1.flip1[25] ;
 wire \thechain[6].chain1.flip1[26] ;
 wire \thechain[6].chain1.flip1[27] ;
 wire \thechain[6].chain1.flip1[28] ;
 wire \thechain[6].chain1.flip1[29] ;
 wire \thechain[6].chain1.flip1[2] ;
 wire \thechain[6].chain1.flip1[30] ;
 wire \thechain[6].chain1.flip1[31] ;
 wire \thechain[6].chain1.flip1[32] ;
 wire \thechain[6].chain1.flip1[33] ;
 wire \thechain[6].chain1.flip1[34] ;
 wire \thechain[6].chain1.flip1[35] ;
 wire \thechain[6].chain1.flip1[36] ;
 wire \thechain[6].chain1.flip1[37] ;
 wire \thechain[6].chain1.flip1[38] ;
 wire \thechain[6].chain1.flip1[39] ;
 wire \thechain[6].chain1.flip1[3] ;
 wire \thechain[6].chain1.flip1[40] ;
 wire \thechain[6].chain1.flip1[41] ;
 wire \thechain[6].chain1.flip1[42] ;
 wire \thechain[6].chain1.flip1[43] ;
 wire \thechain[6].chain1.flip1[44] ;
 wire \thechain[6].chain1.flip1[45] ;
 wire \thechain[6].chain1.flip1[46] ;
 wire \thechain[6].chain1.flip1[47] ;
 wire \thechain[6].chain1.flip1[48] ;
 wire \thechain[6].chain1.flip1[49] ;
 wire \thechain[6].chain1.flip1[4] ;
 wire \thechain[6].chain1.flip1[50] ;
 wire \thechain[6].chain1.flip1[51] ;
 wire \thechain[6].chain1.flip1[52] ;
 wire \thechain[6].chain1.flip1[53] ;
 wire \thechain[6].chain1.flip1[54] ;
 wire \thechain[6].chain1.flip1[55] ;
 wire \thechain[6].chain1.flip1[56] ;
 wire \thechain[6].chain1.flip1[57] ;
 wire \thechain[6].chain1.flip1[58] ;
 wire \thechain[6].chain1.flip1[59] ;
 wire \thechain[6].chain1.flip1[5] ;
 wire \thechain[6].chain1.flip1[60] ;
 wire \thechain[6].chain1.flip1[61] ;
 wire \thechain[6].chain1.flip1[62] ;
 wire \thechain[6].chain1.flip1[63] ;
 wire \thechain[6].chain1.flip1[64] ;
 wire \thechain[6].chain1.flip1[65] ;
 wire \thechain[6].chain1.flip1[66] ;
 wire \thechain[6].chain1.flip1[67] ;
 wire \thechain[6].chain1.flip1[68] ;
 wire \thechain[6].chain1.flip1[69] ;
 wire \thechain[6].chain1.flip1[6] ;
 wire \thechain[6].chain1.flip1[70] ;
 wire \thechain[6].chain1.flip1[71] ;
 wire \thechain[6].chain1.flip1[72] ;
 wire \thechain[6].chain1.flip1[73] ;
 wire \thechain[6].chain1.flip1[74] ;
 wire \thechain[6].chain1.flip1[75] ;
 wire \thechain[6].chain1.flip1[76] ;
 wire \thechain[6].chain1.flip1[77] ;
 wire \thechain[6].chain1.flip1[78] ;
 wire \thechain[6].chain1.flip1[79] ;
 wire \thechain[6].chain1.flip1[7] ;
 wire \thechain[6].chain1.flip1[8] ;
 wire \thechain[6].chain1.flip1[9] ;
 wire \thechain[6].chain1.flip2[0] ;
 wire \thechain[6].chain1.flip2[10] ;
 wire \thechain[6].chain1.flip2[11] ;
 wire \thechain[6].chain1.flip2[12] ;
 wire \thechain[6].chain1.flip2[13] ;
 wire \thechain[6].chain1.flip2[14] ;
 wire \thechain[6].chain1.flip2[15] ;
 wire \thechain[6].chain1.flip2[16] ;
 wire \thechain[6].chain1.flip2[17] ;
 wire \thechain[6].chain1.flip2[18] ;
 wire \thechain[6].chain1.flip2[19] ;
 wire \thechain[6].chain1.flip2[1] ;
 wire \thechain[6].chain1.flip2[20] ;
 wire \thechain[6].chain1.flip2[21] ;
 wire \thechain[6].chain1.flip2[22] ;
 wire \thechain[6].chain1.flip2[23] ;
 wire \thechain[6].chain1.flip2[24] ;
 wire \thechain[6].chain1.flip2[25] ;
 wire \thechain[6].chain1.flip2[26] ;
 wire \thechain[6].chain1.flip2[27] ;
 wire \thechain[6].chain1.flip2[28] ;
 wire \thechain[6].chain1.flip2[29] ;
 wire \thechain[6].chain1.flip2[2] ;
 wire \thechain[6].chain1.flip2[30] ;
 wire \thechain[6].chain1.flip2[31] ;
 wire \thechain[6].chain1.flip2[32] ;
 wire \thechain[6].chain1.flip2[33] ;
 wire \thechain[6].chain1.flip2[34] ;
 wire \thechain[6].chain1.flip2[35] ;
 wire \thechain[6].chain1.flip2[36] ;
 wire \thechain[6].chain1.flip2[37] ;
 wire \thechain[6].chain1.flip2[38] ;
 wire \thechain[6].chain1.flip2[39] ;
 wire \thechain[6].chain1.flip2[3] ;
 wire \thechain[6].chain1.flip2[40] ;
 wire \thechain[6].chain1.flip2[41] ;
 wire \thechain[6].chain1.flip2[42] ;
 wire \thechain[6].chain1.flip2[43] ;
 wire \thechain[6].chain1.flip2[44] ;
 wire \thechain[6].chain1.flip2[45] ;
 wire \thechain[6].chain1.flip2[46] ;
 wire \thechain[6].chain1.flip2[47] ;
 wire \thechain[6].chain1.flip2[48] ;
 wire \thechain[6].chain1.flip2[49] ;
 wire \thechain[6].chain1.flip2[4] ;
 wire \thechain[6].chain1.flip2[50] ;
 wire \thechain[6].chain1.flip2[51] ;
 wire \thechain[6].chain1.flip2[52] ;
 wire \thechain[6].chain1.flip2[53] ;
 wire \thechain[6].chain1.flip2[54] ;
 wire \thechain[6].chain1.flip2[55] ;
 wire \thechain[6].chain1.flip2[56] ;
 wire \thechain[6].chain1.flip2[57] ;
 wire \thechain[6].chain1.flip2[58] ;
 wire \thechain[6].chain1.flip2[59] ;
 wire \thechain[6].chain1.flip2[5] ;
 wire \thechain[6].chain1.flip2[60] ;
 wire \thechain[6].chain1.flip2[61] ;
 wire \thechain[6].chain1.flip2[62] ;
 wire \thechain[6].chain1.flip2[63] ;
 wire \thechain[6].chain1.flip2[64] ;
 wire \thechain[6].chain1.flip2[65] ;
 wire \thechain[6].chain1.flip2[66] ;
 wire \thechain[6].chain1.flip2[67] ;
 wire \thechain[6].chain1.flip2[68] ;
 wire \thechain[6].chain1.flip2[69] ;
 wire \thechain[6].chain1.flip2[6] ;
 wire \thechain[6].chain1.flip2[70] ;
 wire \thechain[6].chain1.flip2[71] ;
 wire \thechain[6].chain1.flip2[72] ;
 wire \thechain[6].chain1.flip2[73] ;
 wire \thechain[6].chain1.flip2[74] ;
 wire \thechain[6].chain1.flip2[75] ;
 wire \thechain[6].chain1.flip2[76] ;
 wire \thechain[6].chain1.flip2[77] ;
 wire \thechain[6].chain1.flip2[78] ;
 wire \thechain[6].chain1.flip2[79] ;
 wire \thechain[6].chain1.flip2[7] ;
 wire \thechain[6].chain1.flip2[8] ;
 wire \thechain[6].chain1.flip2[9] ;
 wire \thechain[7].chain1.dout ;
 wire \thechain[7].chain1.ff[0] ;
 wire \thechain[7].chain1.ff[10] ;
 wire \thechain[7].chain1.ff[11] ;
 wire \thechain[7].chain1.ff[12] ;
 wire \thechain[7].chain1.ff[13] ;
 wire \thechain[7].chain1.ff[14] ;
 wire \thechain[7].chain1.ff[15] ;
 wire \thechain[7].chain1.ff[16] ;
 wire \thechain[7].chain1.ff[17] ;
 wire \thechain[7].chain1.ff[18] ;
 wire \thechain[7].chain1.ff[19] ;
 wire \thechain[7].chain1.ff[1] ;
 wire \thechain[7].chain1.ff[20] ;
 wire \thechain[7].chain1.ff[21] ;
 wire \thechain[7].chain1.ff[22] ;
 wire \thechain[7].chain1.ff[23] ;
 wire \thechain[7].chain1.ff[24] ;
 wire \thechain[7].chain1.ff[25] ;
 wire \thechain[7].chain1.ff[26] ;
 wire \thechain[7].chain1.ff[27] ;
 wire \thechain[7].chain1.ff[28] ;
 wire \thechain[7].chain1.ff[29] ;
 wire \thechain[7].chain1.ff[2] ;
 wire \thechain[7].chain1.ff[30] ;
 wire \thechain[7].chain1.ff[31] ;
 wire \thechain[7].chain1.ff[32] ;
 wire \thechain[7].chain1.ff[33] ;
 wire \thechain[7].chain1.ff[34] ;
 wire \thechain[7].chain1.ff[35] ;
 wire \thechain[7].chain1.ff[36] ;
 wire \thechain[7].chain1.ff[37] ;
 wire \thechain[7].chain1.ff[38] ;
 wire \thechain[7].chain1.ff[39] ;
 wire \thechain[7].chain1.ff[3] ;
 wire \thechain[7].chain1.ff[40] ;
 wire \thechain[7].chain1.ff[41] ;
 wire \thechain[7].chain1.ff[42] ;
 wire \thechain[7].chain1.ff[43] ;
 wire \thechain[7].chain1.ff[44] ;
 wire \thechain[7].chain1.ff[45] ;
 wire \thechain[7].chain1.ff[46] ;
 wire \thechain[7].chain1.ff[47] ;
 wire \thechain[7].chain1.ff[48] ;
 wire \thechain[7].chain1.ff[49] ;
 wire \thechain[7].chain1.ff[4] ;
 wire \thechain[7].chain1.ff[50] ;
 wire \thechain[7].chain1.ff[51] ;
 wire \thechain[7].chain1.ff[52] ;
 wire \thechain[7].chain1.ff[53] ;
 wire \thechain[7].chain1.ff[54] ;
 wire \thechain[7].chain1.ff[55] ;
 wire \thechain[7].chain1.ff[56] ;
 wire \thechain[7].chain1.ff[57] ;
 wire \thechain[7].chain1.ff[58] ;
 wire \thechain[7].chain1.ff[59] ;
 wire \thechain[7].chain1.ff[5] ;
 wire \thechain[7].chain1.ff[60] ;
 wire \thechain[7].chain1.ff[61] ;
 wire \thechain[7].chain1.ff[62] ;
 wire \thechain[7].chain1.ff[63] ;
 wire \thechain[7].chain1.ff[64] ;
 wire \thechain[7].chain1.ff[65] ;
 wire \thechain[7].chain1.ff[66] ;
 wire \thechain[7].chain1.ff[67] ;
 wire \thechain[7].chain1.ff[68] ;
 wire \thechain[7].chain1.ff[69] ;
 wire \thechain[7].chain1.ff[6] ;
 wire \thechain[7].chain1.ff[70] ;
 wire \thechain[7].chain1.ff[71] ;
 wire \thechain[7].chain1.ff[72] ;
 wire \thechain[7].chain1.ff[73] ;
 wire \thechain[7].chain1.ff[74] ;
 wire \thechain[7].chain1.ff[75] ;
 wire \thechain[7].chain1.ff[76] ;
 wire \thechain[7].chain1.ff[77] ;
 wire \thechain[7].chain1.ff[78] ;
 wire \thechain[7].chain1.ff[7] ;
 wire \thechain[7].chain1.ff[8] ;
 wire \thechain[7].chain1.ff[9] ;
 wire \thechain[7].chain1.flip1[0] ;
 wire \thechain[7].chain1.flip1[10] ;
 wire \thechain[7].chain1.flip1[11] ;
 wire \thechain[7].chain1.flip1[12] ;
 wire \thechain[7].chain1.flip1[13] ;
 wire \thechain[7].chain1.flip1[14] ;
 wire \thechain[7].chain1.flip1[15] ;
 wire \thechain[7].chain1.flip1[16] ;
 wire \thechain[7].chain1.flip1[17] ;
 wire \thechain[7].chain1.flip1[18] ;
 wire \thechain[7].chain1.flip1[19] ;
 wire \thechain[7].chain1.flip1[1] ;
 wire \thechain[7].chain1.flip1[20] ;
 wire \thechain[7].chain1.flip1[21] ;
 wire \thechain[7].chain1.flip1[22] ;
 wire \thechain[7].chain1.flip1[23] ;
 wire \thechain[7].chain1.flip1[24] ;
 wire \thechain[7].chain1.flip1[25] ;
 wire \thechain[7].chain1.flip1[26] ;
 wire \thechain[7].chain1.flip1[27] ;
 wire \thechain[7].chain1.flip1[28] ;
 wire \thechain[7].chain1.flip1[29] ;
 wire \thechain[7].chain1.flip1[2] ;
 wire \thechain[7].chain1.flip1[30] ;
 wire \thechain[7].chain1.flip1[31] ;
 wire \thechain[7].chain1.flip1[32] ;
 wire \thechain[7].chain1.flip1[33] ;
 wire \thechain[7].chain1.flip1[34] ;
 wire \thechain[7].chain1.flip1[35] ;
 wire \thechain[7].chain1.flip1[36] ;
 wire \thechain[7].chain1.flip1[37] ;
 wire \thechain[7].chain1.flip1[38] ;
 wire \thechain[7].chain1.flip1[39] ;
 wire \thechain[7].chain1.flip1[3] ;
 wire \thechain[7].chain1.flip1[40] ;
 wire \thechain[7].chain1.flip1[41] ;
 wire \thechain[7].chain1.flip1[42] ;
 wire \thechain[7].chain1.flip1[43] ;
 wire \thechain[7].chain1.flip1[44] ;
 wire \thechain[7].chain1.flip1[45] ;
 wire \thechain[7].chain1.flip1[46] ;
 wire \thechain[7].chain1.flip1[47] ;
 wire \thechain[7].chain1.flip1[48] ;
 wire \thechain[7].chain1.flip1[49] ;
 wire \thechain[7].chain1.flip1[4] ;
 wire \thechain[7].chain1.flip1[50] ;
 wire \thechain[7].chain1.flip1[51] ;
 wire \thechain[7].chain1.flip1[52] ;
 wire \thechain[7].chain1.flip1[53] ;
 wire \thechain[7].chain1.flip1[54] ;
 wire \thechain[7].chain1.flip1[55] ;
 wire \thechain[7].chain1.flip1[56] ;
 wire \thechain[7].chain1.flip1[57] ;
 wire \thechain[7].chain1.flip1[58] ;
 wire \thechain[7].chain1.flip1[59] ;
 wire \thechain[7].chain1.flip1[5] ;
 wire \thechain[7].chain1.flip1[60] ;
 wire \thechain[7].chain1.flip1[61] ;
 wire \thechain[7].chain1.flip1[62] ;
 wire \thechain[7].chain1.flip1[63] ;
 wire \thechain[7].chain1.flip1[64] ;
 wire \thechain[7].chain1.flip1[65] ;
 wire \thechain[7].chain1.flip1[66] ;
 wire \thechain[7].chain1.flip1[67] ;
 wire \thechain[7].chain1.flip1[68] ;
 wire \thechain[7].chain1.flip1[69] ;
 wire \thechain[7].chain1.flip1[6] ;
 wire \thechain[7].chain1.flip1[70] ;
 wire \thechain[7].chain1.flip1[71] ;
 wire \thechain[7].chain1.flip1[72] ;
 wire \thechain[7].chain1.flip1[73] ;
 wire \thechain[7].chain1.flip1[74] ;
 wire \thechain[7].chain1.flip1[75] ;
 wire \thechain[7].chain1.flip1[76] ;
 wire \thechain[7].chain1.flip1[77] ;
 wire \thechain[7].chain1.flip1[78] ;
 wire \thechain[7].chain1.flip1[79] ;
 wire \thechain[7].chain1.flip1[7] ;
 wire \thechain[7].chain1.flip1[8] ;
 wire \thechain[7].chain1.flip1[9] ;
 wire \thechain[7].chain1.flip2[0] ;
 wire \thechain[7].chain1.flip2[10] ;
 wire \thechain[7].chain1.flip2[11] ;
 wire \thechain[7].chain1.flip2[12] ;
 wire \thechain[7].chain1.flip2[13] ;
 wire \thechain[7].chain1.flip2[14] ;
 wire \thechain[7].chain1.flip2[15] ;
 wire \thechain[7].chain1.flip2[16] ;
 wire \thechain[7].chain1.flip2[17] ;
 wire \thechain[7].chain1.flip2[18] ;
 wire \thechain[7].chain1.flip2[19] ;
 wire \thechain[7].chain1.flip2[1] ;
 wire \thechain[7].chain1.flip2[20] ;
 wire \thechain[7].chain1.flip2[21] ;
 wire \thechain[7].chain1.flip2[22] ;
 wire \thechain[7].chain1.flip2[23] ;
 wire \thechain[7].chain1.flip2[24] ;
 wire \thechain[7].chain1.flip2[25] ;
 wire \thechain[7].chain1.flip2[26] ;
 wire \thechain[7].chain1.flip2[27] ;
 wire \thechain[7].chain1.flip2[28] ;
 wire \thechain[7].chain1.flip2[29] ;
 wire \thechain[7].chain1.flip2[2] ;
 wire \thechain[7].chain1.flip2[30] ;
 wire \thechain[7].chain1.flip2[31] ;
 wire \thechain[7].chain1.flip2[32] ;
 wire \thechain[7].chain1.flip2[33] ;
 wire \thechain[7].chain1.flip2[34] ;
 wire \thechain[7].chain1.flip2[35] ;
 wire \thechain[7].chain1.flip2[36] ;
 wire \thechain[7].chain1.flip2[37] ;
 wire \thechain[7].chain1.flip2[38] ;
 wire \thechain[7].chain1.flip2[39] ;
 wire \thechain[7].chain1.flip2[3] ;
 wire \thechain[7].chain1.flip2[40] ;
 wire \thechain[7].chain1.flip2[41] ;
 wire \thechain[7].chain1.flip2[42] ;
 wire \thechain[7].chain1.flip2[43] ;
 wire \thechain[7].chain1.flip2[44] ;
 wire \thechain[7].chain1.flip2[45] ;
 wire \thechain[7].chain1.flip2[46] ;
 wire \thechain[7].chain1.flip2[47] ;
 wire \thechain[7].chain1.flip2[48] ;
 wire \thechain[7].chain1.flip2[49] ;
 wire \thechain[7].chain1.flip2[4] ;
 wire \thechain[7].chain1.flip2[50] ;
 wire \thechain[7].chain1.flip2[51] ;
 wire \thechain[7].chain1.flip2[52] ;
 wire \thechain[7].chain1.flip2[53] ;
 wire \thechain[7].chain1.flip2[54] ;
 wire \thechain[7].chain1.flip2[55] ;
 wire \thechain[7].chain1.flip2[56] ;
 wire \thechain[7].chain1.flip2[57] ;
 wire \thechain[7].chain1.flip2[58] ;
 wire \thechain[7].chain1.flip2[59] ;
 wire \thechain[7].chain1.flip2[5] ;
 wire \thechain[7].chain1.flip2[60] ;
 wire \thechain[7].chain1.flip2[61] ;
 wire \thechain[7].chain1.flip2[62] ;
 wire \thechain[7].chain1.flip2[63] ;
 wire \thechain[7].chain1.flip2[64] ;
 wire \thechain[7].chain1.flip2[65] ;
 wire \thechain[7].chain1.flip2[66] ;
 wire \thechain[7].chain1.flip2[67] ;
 wire \thechain[7].chain1.flip2[68] ;
 wire \thechain[7].chain1.flip2[69] ;
 wire \thechain[7].chain1.flip2[6] ;
 wire \thechain[7].chain1.flip2[70] ;
 wire \thechain[7].chain1.flip2[71] ;
 wire \thechain[7].chain1.flip2[72] ;
 wire \thechain[7].chain1.flip2[73] ;
 wire \thechain[7].chain1.flip2[74] ;
 wire \thechain[7].chain1.flip2[75] ;
 wire \thechain[7].chain1.flip2[76] ;
 wire \thechain[7].chain1.flip2[77] ;
 wire \thechain[7].chain1.flip2[78] ;
 wire \thechain[7].chain1.flip2[79] ;
 wire \thechain[7].chain1.flip2[7] ;
 wire \thechain[7].chain1.flip2[8] ;
 wire \thechain[7].chain1.flip2[9] ;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;

 sky130_fd_sc_hd__dfrtp_1 _000_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[3].chain1.flip1[48] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _001_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[3].chain1.flip1[23] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _002_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[3].chain1.flip1[49] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _003_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[3].chain1.flip1[10] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _004_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[3].chain1.flip1[50] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _005_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[51] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _006_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[52] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _007_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[3].chain1.flip1[9] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _008_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[53] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _009_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[54] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _010_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[55] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _011_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[3].chain1.flip1[8] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _012_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[56] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _013_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[3].chain1.flip1[57] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _014_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[3].chain1.flip1[24] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _015_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[3].chain1.flip1[58] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _016_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[3].chain1.flip1[7] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _017_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[3].chain1.flip1[59] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _018_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[3].chain1.flip1[60] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _019_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[3].chain1.flip1[61] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _020_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[3].chain1.flip1[6] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _021_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[3].chain1.flip1[62] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _022_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[3].chain1.flip1[63] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _023_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[3].chain1.flip1[64] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _024_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[3].chain1.flip1[5] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _025_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[3].chain1.flip1[65] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _026_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[3].chain1.flip1[66] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _027_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[3].chain1.flip1[25] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _028_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[3].chain1.flip1[67] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _029_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[3].chain1.flip1[4] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _030_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[3].chain1.flip1[68] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _031_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[3].chain1.flip1[69] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _032_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[18] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _033_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[3].chain1.flip1[70] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _034_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[3].chain1.flip1[3] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _035_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[3].chain1.flip1[71] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _036_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[3].chain1.flip1[72] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _037_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[3].chain1.flip1[73] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _038_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[3].chain1.flip1[2] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _039_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[3].chain1.flip1[74] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _040_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[3].chain1.flip1[75] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _041_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[3].chain1.flip1[26] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _042_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[3].chain1.flip1[76] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _043_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[3].chain1.flip1[1] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _044_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[3].chain1.flip1[77] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _045_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[3].chain1.flip1[78] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _046_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[3].chain1.flip1[79] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _047_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[3].chain1.flip1[0] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _048_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[4].chain1.flip1[27] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _049_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[4].chain1.flip1[28] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _050_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[17] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _051_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[4].chain1.flip1[29] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _052_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[4].chain1.flip1[30] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _053_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[21] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _054_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[4].chain1.flip1[31] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _055_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[16] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _056_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[4].chain1.flip1[32] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _057_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[4].chain1.flip1[33] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _058_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[20] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _059_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[4].chain1.flip1[34] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _060_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[15] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _061_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[4].chain1.flip1[35] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _062_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[4].chain1.flip1[36] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _063_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[4].chain1.flip1[37] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _064_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[14] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _065_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[4].chain1.flip1[38] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _066_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[39] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _067_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[22] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _068_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[40] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _069_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[13] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _070_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[41] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _071_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[42] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _072_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[19] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _073_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[43] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _074_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[12] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _075_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[44] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _076_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[4].chain1.flip1[45] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _077_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[4].chain1.flip1[46] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _078_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[11] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _079_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[4].chain1.flip1[47] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _080_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[4].chain1.flip1[48] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _081_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[4].chain1.flip1[23] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _082_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[4].chain1.flip1[49] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _083_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[10] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _084_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[4].chain1.flip1[50] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _085_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[4].chain1.flip1[51] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _086_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[52] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _087_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[9] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _088_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[53] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _089_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[54] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _090_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[55] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _091_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[8] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _092_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[56] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _093_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[57] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _094_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[4].chain1.flip1[24] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _095_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[58] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _096_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[4].chain1.flip1[7] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _097_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[59] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _098_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[60] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _099_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[4].chain1.flip1[61] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _100_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[4].chain1.flip1[6] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _101_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[4].chain1.flip1[62] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _102_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[4].chain1.flip1[63] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _103_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[4].chain1.flip1[64] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _104_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[4].chain1.flip1[5] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _105_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[65] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _106_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[66] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _107_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[4].chain1.flip1[25] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _108_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[67] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _109_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[4].chain1.flip1[4] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _110_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[68] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _111_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[69] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _112_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[4].chain1.flip1[18] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _113_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[70] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _114_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[4].chain1.flip1[3] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _115_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[4].chain1.flip1[71] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _116_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[4].chain1.flip1[72] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _117_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[4].chain1.flip1[73] ),
    .RESET_B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _118_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[4].chain1.flip1[2] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _119_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[4].chain1.flip1[74] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _120_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[4].chain1.flip1[75] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _121_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[4].chain1.flip1[26] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _122_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[4].chain1.flip1[76] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _123_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[4].chain1.flip1[1] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _124_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[4].chain1.flip1[77] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _125_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[4].chain1.flip1[78] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _126_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[4].chain1.flip1[79] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _127_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[4].chain1.flip1[0] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _128_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[5].chain1.flip1[27] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _129_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[5].chain1.flip1[28] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _130_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[5].chain1.flip1[17] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _131_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[5].chain1.flip1[29] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _132_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[5].chain1.flip1[30] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _133_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[5].chain1.flip1[21] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _134_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[5].chain1.flip1[31] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _135_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[16] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _136_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[5].chain1.flip1[32] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _137_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[5].chain1.flip1[33] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _138_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[5].chain1.flip1[20] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _139_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[5].chain1.flip1[34] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _140_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[15] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _141_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[5].chain1.flip1[35] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _142_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[5].chain1.flip1[36] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[5].chain1.flip1[37] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[14] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _145_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[5].chain1.flip1[38] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _146_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[5].chain1.flip1[39] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _147_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[5].chain1.flip1[22] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _148_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[40] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _149_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[13] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _150_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[41] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _151_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[42] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _152_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[5].chain1.flip1[19] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _153_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[43] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _154_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[12] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _155_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[44] ),
    .RESET_B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _156_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[45] ),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _157_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[46] ),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _158_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[11] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _159_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[47] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _160_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[48] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _161_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[5].chain1.flip1[23] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _162_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[49] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _163_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[10] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _164_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[50] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _165_ (.CLK(clknet_leaf_31_clk),
    .D(\thechain[5].chain1.flip1[51] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _166_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[5].chain1.flip1[52] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _167_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[9] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _168_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[5].chain1.flip1[53] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _169_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[5].chain1.flip1[54] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _170_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[5].chain1.flip1[55] ),
    .RESET_B(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _171_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[8] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _172_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[5].chain1.flip1[56] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _173_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[5].chain1.flip1[57] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _174_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[5].chain1.flip1[24] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _175_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[5].chain1.flip1[58] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _176_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[7] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _177_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[5].chain1.flip1[59] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _178_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[5].chain1.flip1[60] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _179_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[5].chain1.flip1[61] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _180_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[5].chain1.flip1[6] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _181_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[62] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _182_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[63] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _183_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[64] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _184_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[5].chain1.flip1[5] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _185_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[65] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _186_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[66] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _187_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[5].chain1.flip1[25] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _188_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[67] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _189_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[5].chain1.flip1[4] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _190_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[5].chain1.flip1[68] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _191_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[5].chain1.flip1[69] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _192_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[5].chain1.flip1[18] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _193_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[5].chain1.flip1[70] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _194_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[5].chain1.flip1[3] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _195_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[5].chain1.flip1[71] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _196_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[5].chain1.flip1[72] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _197_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[5].chain1.flip1[73] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _198_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[5].chain1.flip1[2] ),
    .RESET_B(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _199_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[5].chain1.flip1[74] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _200_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[5].chain1.flip1[75] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _201_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[5].chain1.flip1[26] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _202_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[5].chain1.flip1[76] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _203_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[5].chain1.flip1[1] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _204_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[5].chain1.flip1[77] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _205_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[5].chain1.flip1[78] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _206_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[5].chain1.flip1[79] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _207_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[5].chain1.flip1[0] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _208_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[27] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _209_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[28] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _210_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[17] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _211_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[29] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _212_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[30] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _213_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[21] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _214_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[31] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _215_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[16] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _216_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[32] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _217_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[33] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _218_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[20] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _219_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[6].chain1.flip1[34] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _220_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[6].chain1.flip1[15] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _221_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[6].chain1.flip1[35] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _222_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[6].chain1.flip1[36] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _223_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[6].chain1.flip1[37] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _224_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[14] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _225_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[6].chain1.flip1[38] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _226_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[6].chain1.flip1[39] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _227_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[22] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _228_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[6].chain1.flip1[40] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _229_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[13] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _230_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[6].chain1.flip1[41] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _231_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[6].chain1.flip1[42] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _232_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[19] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _233_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[6].chain1.flip1[43] ),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _234_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[12] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _235_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[6].chain1.flip1[44] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _236_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[6].chain1.flip1[45] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _237_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[6].chain1.flip1[46] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _238_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[11] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _239_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[6].chain1.flip1[47] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _240_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[48] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _241_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[23] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _242_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[6].chain1.flip1[49] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _243_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[10] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _244_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[50] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _245_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[51] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _246_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[52] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _247_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[9] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _248_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[53] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _249_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[54] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _250_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[6].chain1.flip1[55] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _251_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[8] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _252_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[6].chain1.flip1[56] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _253_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[6].chain1.flip1[57] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _254_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[24] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _255_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[6].chain1.flip1[58] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _256_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[7] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _257_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[6].chain1.flip1[59] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _258_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[6].chain1.flip1[60] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _259_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[6].chain1.flip1[61] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _260_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[6].chain1.flip1[6] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _261_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[6].chain1.flip1[62] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _262_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[6].chain1.flip1[63] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _263_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[6].chain1.flip1[64] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _264_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[6].chain1.flip1[5] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _265_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[65] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _266_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[66] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _267_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[25] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _268_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[67] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _269_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[6].chain1.flip1[4] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _270_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[68] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _271_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[69] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _272_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[6].chain1.flip1[18] ),
    .RESET_B(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _273_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[70] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _274_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[6].chain1.flip1[3] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _275_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[71] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _276_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[72] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _277_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[73] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _278_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[6].chain1.flip1[2] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _279_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[74] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _280_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[6].chain1.flip1[75] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _281_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[6].chain1.flip1[26] ),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _282_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[6].chain1.flip1[76] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _283_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[6].chain1.flip1[1] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _284_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[6].chain1.flip1[77] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _285_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[6].chain1.flip1[78] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _286_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[6].chain1.flip1[79] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _287_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[6].chain1.flip1[0] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _288_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[27] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _289_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[28] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _290_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[7].chain1.flip1[17] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _291_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[29] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _292_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[30] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _293_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[7].chain1.flip1[21] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _294_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[31] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _295_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[16] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _296_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[32] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _297_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[33] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _298_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[7].chain1.flip1[20] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _299_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[7].chain1.flip1[34] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _300_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[15] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _301_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[7].chain1.flip1[35] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _302_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[7].chain1.flip1[36] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _303_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[7].chain1.flip1[37] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _304_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[14] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _305_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[7].chain1.flip1[38] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _306_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[7].chain1.flip1[39] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _307_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[7].chain1.flip1[22] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _308_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[7].chain1.flip1[40] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _309_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[13] ),
    .RESET_B(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _310_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[7].chain1.flip1[41] ),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _311_ (.CLK(clknet_leaf_1_clk),
    .D(\thechain[7].chain1.flip1[42] ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _312_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[7].chain1.flip1[19] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _313_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[43] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _314_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[12] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _315_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[44] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _316_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[45] ),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _317_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[46] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _318_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[11] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _319_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[47] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _320_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[48] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _321_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[7].chain1.flip1[23] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _322_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[49] ),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _323_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[10] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _324_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[50] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _325_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[7].chain1.flip1[51] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _326_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[7].chain1.flip1[52] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _327_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[7].chain1.flip1[9] ),
    .RESET_B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _328_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[7].chain1.flip1[53] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _329_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[7].chain1.flip1[54] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _330_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[7].chain1.flip1[55] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _331_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[8] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _332_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[7].chain1.flip1[56] ),
    .RESET_B(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _333_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[57] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _334_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[7].chain1.flip1[24] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _335_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[58] ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _336_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[7].chain1.flip1[7] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _337_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[59] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _338_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[60] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _339_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[61] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _340_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[6] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _341_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[62] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _342_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[63] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _343_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[64] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _344_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[5] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _345_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[65] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _346_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[66] ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _347_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[25] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _348_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[67] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _349_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[4] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _350_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[68] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _351_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[69] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _352_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[7].chain1.flip1[18] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _353_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[70] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _354_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[3] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _355_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[71] ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _356_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[72] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _357_ (.CLK(clknet_leaf_7_clk),
    .D(\thechain[7].chain1.flip1[73] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _358_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[2] ),
    .RESET_B(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _359_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[7].chain1.flip1[74] ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _360_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[7].chain1.flip1[75] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _361_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[7].chain1.flip1[26] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _362_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[7].chain1.flip1[76] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _363_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[7].chain1.flip1[1] ),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _364_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[7].chain1.flip1[77] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _365_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[7].chain1.flip1[78] ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _366_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[7].chain1.flip1[79] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _367_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[7].chain1.flip1[0] ),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _368_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[27] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _369_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[28] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _370_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[17] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _371_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[29] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _372_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[30] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _373_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[21] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _374_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[31] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _375_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[16] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _376_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[32] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _377_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[33] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _378_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[20] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _379_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[34] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _380_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[15] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _381_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[35] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _382_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[36] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _383_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[37] ),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _384_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[14] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _385_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[0].chain1.flip1[38] ),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _386_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[39] ),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _387_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[22] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _388_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[40] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _389_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[0].chain1.flip1[13] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _390_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[41] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _391_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[42] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _392_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[19] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _393_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[43] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _394_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[0].chain1.flip1[12] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _395_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[44] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _396_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[45] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _397_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[46] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _398_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[0].chain1.flip1[11] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _399_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[0].chain1.flip1[47] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _400_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[0].chain1.flip1[48] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _401_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[23] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _402_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[0].chain1.flip1[49] ),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _403_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[0].chain1.flip1[10] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _404_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[0].chain1.flip1[50] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _405_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[0].chain1.flip1[51] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _406_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[0].chain1.flip1[52] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _407_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[0].chain1.flip1[9] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _408_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[0].chain1.flip1[53] ),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _409_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[0].chain1.flip1[54] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _410_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[0].chain1.flip1[55] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _411_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[0].chain1.flip1[8] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _412_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[0].chain1.flip1[56] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _413_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[0].chain1.flip1[57] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _414_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[24] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _415_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[0].chain1.flip1[58] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _416_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[7] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _417_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[0].chain1.flip1[59] ),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _418_ (.CLK(clknet_leaf_19_clk),
    .D(\thechain[0].chain1.flip1[60] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _419_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[61] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _420_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[6] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _421_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[62] ),
    .RESET_B(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _422_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[63] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _423_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[64] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _424_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[5] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _425_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[65] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _426_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[0].chain1.flip1[66] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _427_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[25] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _428_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[0].chain1.flip1[67] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _429_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[4] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _430_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[0].chain1.flip1[68] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _431_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[0].chain1.flip1[69] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _432_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[0].chain1.flip1[18] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _433_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[70] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _434_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[3] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _435_ (.CLK(clknet_leaf_11_clk),
    .D(\thechain[0].chain1.flip1[71] ),
    .RESET_B(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _436_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[0].chain1.flip1[72] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _437_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[0].chain1.flip1[73] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _438_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[2] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _439_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[0].chain1.flip1[74] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _440_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[0].chain1.flip1[75] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _441_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[0].chain1.flip1[26] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _442_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[0].chain1.flip1[76] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _443_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[1] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _444_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[0].chain1.flip1[77] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _445_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[0].chain1.flip1[78] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _446_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[0].chain1.flip1[79] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _447_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[0].chain1.flip1[0] ),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _448_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[27] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _449_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[28] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _450_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[17] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _451_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[29] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _452_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[30] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _453_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[21] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _454_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[31] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _455_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[16] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _456_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[32] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _457_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[33] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _458_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[20] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _459_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[34] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _460_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[15] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _461_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[35] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _462_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[36] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _463_ (.CLK(clknet_leaf_23_clk),
    .D(\thechain[1].chain1.flip1[37] ),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[1].chain1.flip1[14] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[1].chain1.flip1[38] ),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _466_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[1].chain1.flip1[39] ),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _467_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[22] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _468_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[1].chain1.flip1[40] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _469_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[1].chain1.flip1[13] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _470_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[1].chain1.flip1[41] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _471_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[1].chain1.flip1[42] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _472_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[19] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _473_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[1].chain1.flip1[43] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _474_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[1].chain1.flip1[12] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _475_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[1].chain1.flip1[44] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _476_ (.CLK(clknet_leaf_26_clk),
    .D(\thechain[1].chain1.flip1[45] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _477_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[1].chain1.flip1[46] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _478_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[1].chain1.flip1[11] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _479_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[1].chain1.flip1[47] ),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _480_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[1].chain1.flip1[48] ),
    .RESET_B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _481_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[23] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _482_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[1].chain1.flip1[49] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _483_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[1].chain1.flip1[10] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _484_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[1].chain1.flip1[50] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _485_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[1].chain1.flip1[51] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _486_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[1].chain1.flip1[52] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _487_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[1].chain1.flip1[9] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _488_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[1].chain1.flip1[53] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _489_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[1].chain1.flip1[54] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _490_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[1].chain1.flip1[55] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _491_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[1].chain1.flip1[8] ),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _492_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[1].chain1.flip1[56] ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _493_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[1].chain1.flip1[57] ),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _494_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[1].chain1.flip1[24] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _495_ (.CLK(clknet_leaf_27_clk),
    .D(\thechain[1].chain1.flip1[58] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _496_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[7] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _497_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[1].chain1.flip1[59] ),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _498_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[1].chain1.flip1[60] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _499_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[1].chain1.flip1[61] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[6] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _501_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[1].chain1.flip1[62] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[1].chain1.flip1[63] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _503_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[1].chain1.flip1[64] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _504_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[5] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _505_ (.CLK(clknet_leaf_3_clk),
    .D(\thechain[1].chain1.flip1[65] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[1].chain1.flip1[66] ),
    .RESET_B(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _507_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[1].chain1.flip1[25] ),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _508_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[1].chain1.flip1[67] ),
    .RESET_B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _509_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[4] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _510_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[68] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _511_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[69] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[1].chain1.flip1[18] ),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _513_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[70] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _514_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[3] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _515_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[71] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _516_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[72] ),
    .RESET_B(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _517_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[73] ),
    .RESET_B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _518_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[2] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _519_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[1].chain1.flip1[74] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(clknet_leaf_12_clk),
    .D(\thechain[1].chain1.flip1[75] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _521_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[1].chain1.flip1[26] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _522_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[1].chain1.flip1[76] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _523_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[1].chain1.flip1[1] ),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[1].chain1.flip1[77] ),
    .RESET_B(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _525_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[1].chain1.flip1[78] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _526_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[1].chain1.flip1[79] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _527_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[1].chain1.flip1[0] ),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _528_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[27] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _529_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[28] ),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _530_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[2].chain1.flip1[17] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _531_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[29] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _532_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[30] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _533_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[2].chain1.flip1[21] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _534_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[31] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _535_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[2].chain1.flip1[16] ),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _536_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[32] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _537_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[33] ),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _538_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[2].chain1.flip1[20] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _539_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[34] ),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _540_ (.CLK(clknet_leaf_21_clk),
    .D(\thechain[2].chain1.flip1[15] ),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _541_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[35] ),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _542_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[36] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _543_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[37] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _544_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[2].chain1.flip1[14] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _545_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[38] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _546_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[2].chain1.flip1[39] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _547_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[2].chain1.flip1[22] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _548_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[2].chain1.flip1[40] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _549_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[2].chain1.flip1[13] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _550_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[2].chain1.flip1[41] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _551_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[2].chain1.flip1[42] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _552_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[2].chain1.flip1[19] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _553_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[2].chain1.flip1[43] ),
    .RESET_B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _554_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[2].chain1.flip1[12] ),
    .RESET_B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _555_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[2].chain1.flip1[44] ),
    .RESET_B(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _556_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[2].chain1.flip1[45] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _557_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[2].chain1.flip1[46] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _558_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[2].chain1.flip1[11] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _559_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[2].chain1.flip1[47] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[47] ));
 sky130_fd_sc_hd__dfrtp_1 _560_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[2].chain1.flip1[48] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[48] ));
 sky130_fd_sc_hd__dfrtp_1 _561_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[2].chain1.flip1[23] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[23] ));
 sky130_fd_sc_hd__dfrtp_1 _562_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[2].chain1.flip1[49] ),
    .RESET_B(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[49] ));
 sky130_fd_sc_hd__dfrtp_1 _563_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[2].chain1.flip1[10] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[10] ));
 sky130_fd_sc_hd__dfrtp_1 _564_ (.CLK(clknet_leaf_28_clk),
    .D(\thechain[2].chain1.flip1[50] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[50] ));
 sky130_fd_sc_hd__dfrtp_1 _565_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[2].chain1.flip1[51] ),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[51] ));
 sky130_fd_sc_hd__dfrtp_1 _566_ (.CLK(clknet_leaf_0_clk),
    .D(\thechain[2].chain1.flip1[52] ),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[52] ));
 sky130_fd_sc_hd__dfrtp_1 _567_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[2].chain1.flip1[9] ),
    .RESET_B(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[9] ));
 sky130_fd_sc_hd__dfrtp_1 _568_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[2].chain1.flip1[53] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[53] ));
 sky130_fd_sc_hd__dfrtp_1 _569_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[2].chain1.flip1[54] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[54] ));
 sky130_fd_sc_hd__dfrtp_1 _570_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[2].chain1.flip1[55] ),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[55] ));
 sky130_fd_sc_hd__dfrtp_1 _571_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[2].chain1.flip1[8] ),
    .RESET_B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[8] ));
 sky130_fd_sc_hd__dfrtp_1 _572_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[2].chain1.flip1[56] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[56] ));
 sky130_fd_sc_hd__dfrtp_1 _573_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[2].chain1.flip1[57] ),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[57] ));
 sky130_fd_sc_hd__dfrtp_1 _574_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[2].chain1.flip1[24] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[24] ));
 sky130_fd_sc_hd__dfrtp_1 _575_ (.CLK(clknet_leaf_2_clk),
    .D(\thechain[2].chain1.flip1[58] ),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[58] ));
 sky130_fd_sc_hd__dfrtp_1 _576_ (.CLK(clknet_leaf_16_clk),
    .D(\thechain[2].chain1.flip1[7] ),
    .RESET_B(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[7] ));
 sky130_fd_sc_hd__dfrtp_1 _577_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[2].chain1.flip1[59] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[59] ));
 sky130_fd_sc_hd__dfrtp_1 _578_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[2].chain1.flip1[60] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[60] ));
 sky130_fd_sc_hd__dfrtp_1 _579_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[2].chain1.flip1[61] ),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[61] ));
 sky130_fd_sc_hd__dfrtp_1 _580_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[2].chain1.flip1[6] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _581_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[2].chain1.flip1[62] ),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[62] ));
 sky130_fd_sc_hd__dfrtp_1 _582_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[2].chain1.flip1[63] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[63] ));
 sky130_fd_sc_hd__dfrtp_1 _583_ (.CLK(clknet_leaf_4_clk),
    .D(\thechain[2].chain1.flip1[64] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[64] ));
 sky130_fd_sc_hd__dfrtp_1 _584_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[2].chain1.flip1[5] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _585_ (.CLK(clknet_leaf_5_clk),
    .D(\thechain[2].chain1.flip1[65] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[65] ));
 sky130_fd_sc_hd__dfrtp_1 _586_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[2].chain1.flip1[66] ),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[66] ));
 sky130_fd_sc_hd__dfrtp_1 _587_ (.CLK(clknet_leaf_22_clk),
    .D(\thechain[2].chain1.flip1[25] ),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[25] ));
 sky130_fd_sc_hd__dfrtp_1 _588_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[2].chain1.flip1[67] ),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[67] ));
 sky130_fd_sc_hd__dfrtp_1 _589_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[2].chain1.flip1[4] ),
    .RESET_B(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[4] ));
 sky130_fd_sc_hd__dfrtp_1 _590_ (.CLK(clknet_leaf_6_clk),
    .D(\thechain[2].chain1.flip1[68] ),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[68] ));
 sky130_fd_sc_hd__dfrtp_1 _591_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[2].chain1.flip1[69] ),
    .RESET_B(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[69] ));
 sky130_fd_sc_hd__dfrtp_1 _592_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[2].chain1.flip1[18] ),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _593_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[2].chain1.flip1[70] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[70] ));
 sky130_fd_sc_hd__dfrtp_1 _594_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[2].chain1.flip1[3] ),
    .RESET_B(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[3] ));
 sky130_fd_sc_hd__dfrtp_1 _595_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[2].chain1.flip1[71] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[71] ));
 sky130_fd_sc_hd__dfrtp_1 _596_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[2].chain1.flip1[72] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[72] ));
 sky130_fd_sc_hd__dfrtp_1 _597_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[2].chain1.flip1[73] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[73] ));
 sky130_fd_sc_hd__dfrtp_1 _598_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[2].chain1.flip1[2] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[2] ));
 sky130_fd_sc_hd__dfrtp_1 _599_ (.CLK(clknet_leaf_8_clk),
    .D(\thechain[2].chain1.flip1[74] ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[74] ));
 sky130_fd_sc_hd__dfrtp_1 _600_ (.CLK(clknet_leaf_10_clk),
    .D(\thechain[2].chain1.flip1[75] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[75] ));
 sky130_fd_sc_hd__dfrtp_1 _601_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[2].chain1.flip1[26] ),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[26] ));
 sky130_fd_sc_hd__dfrtp_1 _602_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[2].chain1.flip1[76] ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[76] ));
 sky130_fd_sc_hd__dfrtp_1 _603_ (.CLK(clknet_leaf_15_clk),
    .D(\thechain[2].chain1.flip1[1] ),
    .RESET_B(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[1] ));
 sky130_fd_sc_hd__dfrtp_1 _604_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[2].chain1.flip1[77] ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[77] ));
 sky130_fd_sc_hd__dfrtp_1 _605_ (.CLK(clknet_leaf_9_clk),
    .D(\thechain[2].chain1.flip1[78] ),
    .RESET_B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[78] ));
 sky130_fd_sc_hd__dfrtp_1 _606_ (.CLK(clknet_leaf_13_clk),
    .D(\thechain[2].chain1.flip1[79] ),
    .RESET_B(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _607_ (.CLK(clknet_leaf_14_clk),
    .D(\thechain[2].chain1.flip1[0] ),
    .RESET_B(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.ff[0] ));
 sky130_fd_sc_hd__dfrtp_1 _608_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[27] ),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[27] ));
 sky130_fd_sc_hd__dfrtp_1 _609_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[28] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[28] ));
 sky130_fd_sc_hd__dfrtp_1 _610_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[17] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _611_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[29] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[29] ));
 sky130_fd_sc_hd__dfrtp_1 _612_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[30] ),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[30] ));
 sky130_fd_sc_hd__dfrtp_1 _613_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[21] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _614_ (.CLK(clknet_leaf_24_clk),
    .D(\thechain[3].chain1.flip1[31] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[31] ));
 sky130_fd_sc_hd__dfrtp_1 _615_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[16] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _616_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[32] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[32] ));
 sky130_fd_sc_hd__dfrtp_1 _617_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[33] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[33] ));
 sky130_fd_sc_hd__dfrtp_1 _618_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[20] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _619_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[34] ),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[34] ));
 sky130_fd_sc_hd__dfrtp_1 _620_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[15] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _621_ (.CLK(clknet_leaf_25_clk),
    .D(\thechain[3].chain1.flip1[35] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[35] ));
 sky130_fd_sc_hd__dfrtp_1 _622_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[36] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[36] ));
 sky130_fd_sc_hd__dfrtp_1 _623_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[37] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[37] ));
 sky130_fd_sc_hd__dfrtp_1 _624_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[3].chain1.flip1[14] ),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _625_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[38] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[38] ));
 sky130_fd_sc_hd__dfrtp_1 _626_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[39] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[39] ));
 sky130_fd_sc_hd__dfrtp_1 _627_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[22] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _628_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[40] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[40] ));
 sky130_fd_sc_hd__dfrtp_1 _629_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[3].chain1.flip1[13] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _630_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[41] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[41] ));
 sky130_fd_sc_hd__dfrtp_1 _631_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[42] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[42] ));
 sky130_fd_sc_hd__dfrtp_1 _632_ (.CLK(clknet_leaf_20_clk),
    .D(\thechain[3].chain1.flip1[19] ),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _633_ (.CLK(clknet_leaf_29_clk),
    .D(\thechain[3].chain1.flip1[43] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[43] ));
 sky130_fd_sc_hd__dfrtp_1 _634_ (.CLK(clknet_leaf_17_clk),
    .D(\thechain[3].chain1.flip1[12] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _635_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[3].chain1.flip1[44] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[44] ));
 sky130_fd_sc_hd__dfrtp_1 _636_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[3].chain1.flip1[45] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[45] ));
 sky130_fd_sc_hd__dfrtp_1 _637_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[3].chain1.flip1[46] ),
    .RESET_B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[46] ));
 sky130_fd_sc_hd__dfrtp_1 _638_ (.CLK(clknet_leaf_18_clk),
    .D(\thechain[3].chain1.flip1[11] ),
    .RESET_B(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[11] ));
 sky130_fd_sc_hd__dfrtp_1 _639_ (.CLK(clknet_leaf_30_clk),
    .D(\thechain[3].chain1.flip1[47] ),
    .RESET_B(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.ff[47] ));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net92));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net93));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net94));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net95));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net96));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net97));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net98));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net99));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net100));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net101));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net102));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net103));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net104));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net105));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net106));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__buf_2 _656_ (.A(\thechain[0].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _657_ (.A(\thechain[1].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _658_ (.A(\thechain[2].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _659_ (.A(\thechain[3].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _660_ (.A(\thechain[4].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _661_ (.A(\thechain[5].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _662_ (.A(\thechain[6].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _663_ (.A(\thechain[7].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_gate_0/_0_  (.A(\thechain[0].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_gate_1/_0_  (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net408),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net455),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net376),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net670),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net605),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net290),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net296),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net372),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net332),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net632),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net477),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net669),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net445),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net709),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net517),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net400),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net617),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net304),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net335),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net636),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net406),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net580),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net610),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net572),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net421),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net685),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net469),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net329),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net303),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net552),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net506),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net597),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net403),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net489),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net728),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net394),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net665),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net533),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net375),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net647),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net737),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net285),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net522),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net591),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net305),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net492),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net725),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[0].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_gate_0/_0_  (.A(\thechain[1].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_gate_1/_0_  (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net255),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net271),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net463),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net430),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net565),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net384),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net590),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net401),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net405),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net486),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net697),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net396),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net562),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net461),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net568),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net409),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net541),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net619),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net246),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net213),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net444),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net452),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net681),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net614),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net392),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net661),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net482),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net721),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net393),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net443),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net624),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net548),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net578),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net466),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net267),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net410),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net637),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net557),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net716),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net646),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net553),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net511),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net490),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net586),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net675),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net436),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net712),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net479),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net736),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net654),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net343),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net500),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net706),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[1].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_gate_0/_0_  (.A(\thechain[2].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_gate_1/_0_  (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net334),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net440),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net423),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net711),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net473),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net317),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net448),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net485),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net583),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net628),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net538),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net603),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net501),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net641),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net383),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net488),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net678),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net453),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net698),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net600),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net644),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net680),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net404),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net598),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net505),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net664),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net286),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net551),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net496),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net663),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net693),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net281),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net402),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net579),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net640),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net355),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net713),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net260),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net581),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net340),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net615),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net560),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net717),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net537),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net707),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net702),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net569),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[2].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_gate_0/_0_  (.A(\thechain[3].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_gate_1/_0_  (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net438),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net729),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net734),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net655),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net341),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net575),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net660),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net634),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net516),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net164),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net662),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net602),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net478),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net631),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net556),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net398),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net535),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net468),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net692),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net566),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net499),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net518),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net431),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net554),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net673),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net351),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net428),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net306),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net497),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net435),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net630),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net513),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net691),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net611),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net454),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net649),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net442),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net314),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net354),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net386),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net544),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net481),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net416),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net714),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net720),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net390),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net531),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[3].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_gate_0/_0_  (.A(\thechain[4].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_gate_1/_0_  (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net356),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net574),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net621),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net459),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net456),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net524),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net399),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net599),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net526),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net652),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net606),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net613),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net677),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net639),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net699),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net648),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net472),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net498),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net389),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net558),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net674),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net415),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net595),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net688),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net391),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net266),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net427),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net411),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net534),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net687),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net520),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net679),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net385),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net507),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net588),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net559),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net484),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net620),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net464),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net577),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net302),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net726),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net457),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net724),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net268),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net642),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net433),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net297),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net635),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net495),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net504),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net672),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net491),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net567),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net434),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net412),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[4].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net414),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_gate_0/_0_  (.A(\thechain[5].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_gate_1/_0_  (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net487),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net483),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net371),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net585),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net458),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net493),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net555),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net467),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net494),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net683),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net625),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net666),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net352),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net576),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net539),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net564),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net570),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net668),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net608),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net604),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net561),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net449),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net422),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net503),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net540),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net701),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net659),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net607),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net584),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net563),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net381),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net319),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net502),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net379),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net547),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net387),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net474),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net710),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net732),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net465),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net510),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net417),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net470),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net397),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net475),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net718),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net612),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net347),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net284),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net362),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net629),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net480),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net627),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net658),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[5].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net527),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_gate_0/_0_  (.A(\thechain[6].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_gate_1/_0_  (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net407),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net339),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net447),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net545),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net638),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net462),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net622),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net723),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net364),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net509),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net420),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net519),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net288),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net686),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net684),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net532),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net413),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net353),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net300),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net571),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net594),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net616),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net593),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net596),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net425),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net437),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net682),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net429),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net738),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net546),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net643),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net450),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net550),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net382),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net727),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net514),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net298),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net536),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net671),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net301),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net719),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net676),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net378),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net476),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net694),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net282),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net689),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net441),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net525),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net528),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net346),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[6].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net235),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.flip2[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_gate_0/_0_  (.A(\thechain[7].chain1.flip2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_gate_1/_0_  (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[0] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[10].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[10].inv_gate_3/_0_  (.A(net292),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[11].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[11].inv_gate_3/_0_  (.A(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[12].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[12].inv_gate_3/_0_  (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[13].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[13].inv_gate_3/_0_  (.A(net418),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[14].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[14].inv_gate_3/_0_  (.A(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[15].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[15].inv_gate_3/_0_  (.A(net633),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[16].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[16].inv_gate_3/_0_  (.A(net366),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[17].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[17].inv_gate_3/_0_  (.A(net609),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[18].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[18].inv_gate_3/_0_  (.A(net360),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[19].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[19].inv_gate_3/_0_  (.A(net373),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[1].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[1].inv_gate_3/_0_  (.A(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[20].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[20].inv_gate_3/_0_  (.A(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[21].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[21].inv_gate_3/_0_  (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[22].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[22].inv_gate_3/_0_  (.A(net735),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[23].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[23].inv_gate_3/_0_  (.A(net388),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[24].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[24].inv_gate_3/_0_  (.A(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[25].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[25].inv_gate_3/_0_  (.A(net731),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[26].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[26].inv_gate_3/_0_  (.A(net650),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[27].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[27].inv_gate_3/_0_  (.A(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[28].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[28].inv_gate_3/_0_  (.A(net308),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[29].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[29].inv_gate_3/_0_  (.A(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[2].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[2].inv_gate_3/_0_  (.A(net730),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[30].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[30].inv_gate_3/_0_  (.A(net645),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[31].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[31].inv_gate_3/_0_  (.A(net521),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[32].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[32].inv_gate_3/_0_  (.A(net265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[33].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[33].inv_gate_3/_0_  (.A(net247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[34].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[34].inv_gate_3/_0_  (.A(net283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[35].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[35].inv_gate_3/_0_  (.A(net587),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[36].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[36].inv_gate_3/_0_  (.A(net601),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[37].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[37].inv_gate_3/_0_  (.A(net695),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[38].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[38].inv_gate_3/_0_  (.A(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[39].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[39].inv_gate_3/_0_  (.A(net311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[3].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[3].inv_gate_3/_0_  (.A(net363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[40].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[40].inv_gate_3/_0_  (.A(net733),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[41].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[41].inv_gate_3/_0_  (.A(net419),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[42].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[42].inv_gate_3/_0_  (.A(net704),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[43].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[43].inv_gate_3/_0_  (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[44].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[44].inv_gate_3/_0_  (.A(net365),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[45].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[45].inv_gate_3/_0_  (.A(net512),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[46].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[46].inv_gate_3/_0_  (.A(net549),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[47].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[47].inv_gate_3/_0_  (.A(net623),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[48].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[48].inv_gate_3/_0_  (.A(net336),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[49].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[49].inv_gate_3/_0_  (.A(net374),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[4].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[4].inv_gate_3/_0_  (.A(net589),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[50].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[50].inv_gate_3/_0_  (.A(net523),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[51].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[51].inv_gate_3/_0_  (.A(net432),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[52].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[52].inv_gate_3/_0_  (.A(net715),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[53].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[53].inv_gate_3/_0_  (.A(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[54].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[54].inv_gate_3/_0_  (.A(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[55].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[55].inv_gate_3/_0_  (.A(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[56].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[56].inv_gate_3/_0_  (.A(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[57].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[57].inv_gate_3/_0_  (.A(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[58].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[58].inv_gate_3/_0_  (.A(net369),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[59].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[59].inv_gate_3/_0_  (.A(net231),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[5].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[5].inv_gate_3/_0_  (.A(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[60].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[60].inv_gate_3/_0_  (.A(net316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[61].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[61].inv_gate_3/_0_  (.A(net245),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[62].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[62].inv_gate_3/_0_  (.A(net328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[63].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[63].inv_gate_3/_0_  (.A(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[64].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[64].inv_gate_3/_0_  (.A(net690),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[65].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[65].inv_gate_3/_0_  (.A(net295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[66].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[66].inv_gate_3/_0_  (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[67].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[67].inv_gate_3/_0_  (.A(net696),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[68].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[68].inv_gate_3/_0_  (.A(net508),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[69].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[69].inv_gate_3/_0_  (.A(net657),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[6].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[6].inv_gate_3/_0_  (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[70].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[70].inv_gate_3/_0_  (.A(net348),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[71].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[71].inv_gate_3/_0_  (.A(net582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[72].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[72].inv_gate_3/_0_  (.A(net515),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[73].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[73].inv_gate_3/_0_  (.A(net705),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[74].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[74].inv_gate_3/_0_  (.A(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[75].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[75].inv_gate_3/_0_  (.A(net573),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[76].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[76].inv_gate_3/_0_  (.A(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[77].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[77].inv_gate_3/_0_  (.A(net667),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[78].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[78].inv_gate_3/_0_  (.A(net700),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[79].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[79].inv_gate_3/_0_  (.A(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[7].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[7].inv_gate_3/_0_  (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[8].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[8].inv_gate_3/_0_  (.A(net722),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[9].inv_gate_2/_0_  (.A(\thechain[7].chain1.flip2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip1[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[9].inv_gate_3/_0_  (.A(net160),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.flip2[9] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout49 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 fanout60 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout70 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout84 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__conb_1 tt_um_regfield_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net91));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_leaf_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_leaf_1_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_leaf_27_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_leaf_28_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_leaf_29_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_leaf_30_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_leaf_31_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload7 (.A(clknet_leaf_20_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_leaf_21_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload9 (.A(clknet_leaf_22_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_leaf_23_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload11 (.A(clknet_leaf_24_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload12 (.A(clknet_leaf_25_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload13 (.A(clknet_leaf_26_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_leaf_3_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload15 (.A(clknet_leaf_4_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload16 (.A(clknet_leaf_6_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload17 (.A(clknet_leaf_7_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_leaf_9_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload19 (.A(clknet_leaf_10_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload20 (.A(clknet_leaf_11_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload21 (.A(clknet_leaf_12_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload22 (.A(clknet_leaf_13_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload23 (.A(clknet_leaf_14_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_leaf_15_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload25 (.A(clknet_leaf_16_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload26 (.A(clknet_leaf_17_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\thechain[4].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\thechain[0].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\thechain[5].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\thechain[5].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\thechain[7].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\thechain[7].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\thechain[5].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\thechain[7].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\thechain[3].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\thechain[2].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\thechain[3].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\thechain[4].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\thechain[7].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\thechain[2].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\thechain[1].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\thechain[6].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\thechain[4].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\thechain[0].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\thechain[4].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\thechain[1].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\thechain[6].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\thechain[3].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\thechain[3].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\thechain[3].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\thechain[6].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\thechain[2].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\thechain[5].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\thechain[7].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\thechain[0].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\thechain[6].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\thechain[4].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\thechain[1].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\thechain[5].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\thechain[0].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\thechain[2].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\thechain[5].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\thechain[7].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\thechain[2].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\thechain[2].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\thechain[3].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\thechain[3].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\thechain[4].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\thechain[0].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\thechain[1].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\thechain[2].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\thechain[2].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\thechain[2].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\thechain[2].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\thechain[0].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\thechain[5].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\thechain[2].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\thechain[2].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\thechain[0].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\thechain[7].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\thechain[7].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\thechain[2].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\thechain[6].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\thechain[3].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\thechain[2].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\thechain[5].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\thechain[6].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\thechain[6].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\thechain[1].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\thechain[2].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\thechain[7].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\thechain[4].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\thechain[5].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\thechain[7].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\thechain[1].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\thechain[5].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\thechain[6].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\thechain[5].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\thechain[3].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\thechain[4].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\thechain[3].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\thechain[2].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\thechain[3].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\thechain[7].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\thechain[1].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\thechain[3].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\thechain[3].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\thechain[7].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\thechain[4].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\thechain[6].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\thechain[1].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\thechain[4].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\thechain[6].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\thechain[1].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\thechain[6].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\thechain[5].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\thechain[3].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\thechain[1].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\thechain[3].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\thechain[7].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\thechain[4].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\thechain[0].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\thechain[3].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\thechain[3].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\thechain[2].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\thechain[7].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\thechain[3].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\thechain[3].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\thechain[0].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\thechain[1].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\thechain[7].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\thechain[3].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\thechain[1].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\thechain[2].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\thechain[6].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\thechain[2].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\thechain[7].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\thechain[7].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\thechain[5].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\thechain[5].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\thechain[0].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\thechain[3].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\thechain[3].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\thechain[3].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\thechain[2].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\thechain[7].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\thechain[1].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\thechain[0].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\thechain[2].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\thechain[3].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\thechain[7].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\thechain[2].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\thechain[4].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\thechain[1].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\thechain[6].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\thechain[0].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\thechain[4].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\thechain[0].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\thechain[7].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\thechain[4].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\thechain[5].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\thechain[3].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\thechain[1].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\thechain[7].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\thechain[7].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\thechain[1].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\thechain[7].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\thechain[1].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\thechain[5].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\thechain[7].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\thechain[0].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\thechain[1].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\thechain[5].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\thechain[6].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\thechain[1].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\thechain[5].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\thechain[3].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\thechain[3].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\thechain[5].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\thechain[2].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\thechain[2].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\thechain[1].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\thechain[6].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\thechain[3].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\thechain[7].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\thechain[4].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\thechain[1].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\thechain[4].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\thechain[3].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\thechain[0].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\thechain[1].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\thechain[2].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\thechain[7].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\thechain[0].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\thechain[5].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\thechain[7].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\thechain[1].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\thechain[0].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\thechain[0].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\thechain[4].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\thechain[2].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\thechain[6].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\thechain[7].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\thechain[5].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\thechain[0].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\thechain[2].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\thechain[4].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\thechain[6].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\thechain[5].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\thechain[0].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\thechain[0].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\thechain[7].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\thechain[1].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\thechain[1].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\thechain[7].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\thechain[0].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\thechain[4].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\thechain[6].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\thechain[5].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\thechain[6].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\thechain[6].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\thechain[4].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\thechain[0].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\thechain[0].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\thechain[0].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\thechain[3].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\thechain[2].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\thechain[7].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\thechain[0].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\thechain[2].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\thechain[7].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\thechain[0].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\thechain[7].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\thechain[3].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\thechain[4].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\thechain[7].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\thechain[2].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\thechain[0].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\thechain[5].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\thechain[0].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\thechain[0].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\thechain[0].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\thechain[6].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\thechain[6].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\thechain[5].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\thechain[1].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\thechain[6].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\thechain[7].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\thechain[0].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\thechain[6].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\thechain[4].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\thechain[0].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\thechain[0].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\thechain[2].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\thechain[0].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\thechain[7].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\thechain[1].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\thechain[0].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\thechain[6].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\thechain[2].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\thechain[3].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\thechain[6].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\thechain[1].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\thechain[6].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\thechain[7].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\thechain[6].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\thechain[5].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\thechain[7].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\thechain[3].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\thechain[1].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\thechain[3].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\thechain[5].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\thechain[6].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\thechain[3].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\thechain[2].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\thechain[4].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\thechain[1].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\thechain[2].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\thechain[2].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\thechain[7].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\thechain[2].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\thechain[5].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\thechain[7].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\thechain[6].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\thechain[7].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\thechain[7].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\thechain[1].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\thechain[0].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\thechain[7].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\thechain[0].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\thechain[5].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\thechain[0].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\thechain[7].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\thechain[7].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\thechain[0].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\thechain[0].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\thechain[6].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\thechain[6].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\thechain[5].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\thechain[2].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\thechain[5].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\thechain[6].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\thechain[2].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\thechain[1].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\thechain[4].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\thechain[3].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\thechain[5].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\thechain[7].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\thechain[4].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\thechain[3].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\thechain[4].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\thechain[1].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\thechain[1].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\thechain[0].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\thechain[0].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\thechain[1].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\thechain[5].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\thechain[3].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\thechain[4].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\thechain[0].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\thechain[1].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\thechain[2].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\thechain[0].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\thechain[2].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\thechain[1].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\thechain[0].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\thechain[6].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\thechain[0].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\thechain[1].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\thechain[1].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\thechain[4].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\thechain[4].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\thechain[6].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\thechain[4].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\thechain[4].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\thechain[3].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\thechain[5].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\thechain[7].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\thechain[7].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\thechain[6].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\thechain[0].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\thechain[5].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\thechain[2].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\thechain[2].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\thechain[6].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\thechain[2].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\thechain[4].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\thechain[3].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\thechain[6].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\thechain[1].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\thechain[3].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\thechain[7].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\thechain[4].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\thechain[4].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\thechain[3].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\thechain[1].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\thechain[6].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\thechain[3].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\thechain[4].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\thechain[2].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\thechain[6].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\thechain[3].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\thechain[1].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\thechain[1].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\thechain[0].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\thechain[6].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\thechain[6].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\thechain[2].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\thechain[5].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\thechain[6].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\thechain[6].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\thechain[1].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\thechain[2].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\thechain[3].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\thechain[0].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\thechain[4].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\thechain[4].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\thechain[5].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\thechain[4].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\thechain[5].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\thechain[1].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\thechain[6].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\thechain[1].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\thechain[4].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\thechain[5].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\thechain[1].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\thechain[5].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\thechain[3].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\thechain[0].chain1.ff[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\thechain[5].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\thechain[6].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\thechain[4].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\thechain[2].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\thechain[5].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\thechain[5].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\thechain[6].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\thechain[0].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\thechain[3].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\thechain[1].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\thechain[5].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\thechain[3].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\thechain[1].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\thechain[5].chain1.ff[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\thechain[4].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\thechain[2].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\thechain[1].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\thechain[5].chain1.ff[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\thechain[2].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\thechain[0].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\thechain[1].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\thechain[4].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\thechain[0].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\thechain[5].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\thechain[5].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\thechain[4].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\thechain[2].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\thechain[3].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\thechain[4].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\thechain[3].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\thechain[1].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\thechain[2].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\thechain[5].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\thechain[5].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\thechain[4].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\thechain[2].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\thechain[0].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\thechain[4].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\thechain[7].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\thechain[6].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\thechain[5].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\thechain[1].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\thechain[7].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\thechain[3].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\thechain[6].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\thechain[7].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\thechain[3].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\thechain[0].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\thechain[3].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\thechain[6].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\thechain[4].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\thechain[7].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\thechain[0].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\thechain[7].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\thechain[4].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\thechain[6].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\thechain[4].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\thechain[5].chain1.ff[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\thechain[6].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\thechain[6].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\thechain[3].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\thechain[3].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\thechain[6].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\thechain[0].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\thechain[4].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\thechain[3].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\thechain[6].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\thechain[2].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\thechain[2].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\thechain[5].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\thechain[5].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\thechain[1].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\thechain[0].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\thechain[6].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\thechain[3].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\thechain[6].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\thechain[6].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\thechain[5].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\thechain[1].chain1.ff[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\thechain[7].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\thechain[6].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\thechain[2].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\thechain[0].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\thechain[1].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\thechain[3].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\thechain[5].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\thechain[3].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\thechain[1].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\thechain[4].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\thechain[4].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\thechain[2].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\thechain[5].chain1.ff[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\thechain[1].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\thechain[5].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\thechain[5].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\thechain[1].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\thechain[3].chain1.ff[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\thechain[4].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\thechain[1].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\thechain[2].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\thechain[5].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\thechain[6].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\thechain[0].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\thechain[7].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\thechain[4].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\thechain[3].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\thechain[5].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\thechain[4].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\thechain[1].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\thechain[2].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\thechain[0].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\thechain[2].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\thechain[7].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\thechain[2].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\thechain[5].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\thechain[5].chain1.ff[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\thechain[1].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\thechain[7].chain1.ff[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\thechain[4].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\thechain[7].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\thechain[1].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\thechain[0].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\thechain[6].chain1.ff[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\thechain[6].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\thechain[6].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\thechain[4].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\thechain[6].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\thechain[0].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\thechain[2].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\thechain[4].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\thechain[2].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\thechain[7].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\thechain[3].chain1.ff[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\thechain[2].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\thechain[5].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\thechain[0].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\thechain[4].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\thechain[5].chain1.ff[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\thechain[5].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\thechain[7].chain1.ff[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\thechain[0].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\thechain[3].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\thechain[5].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\thechain[4].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\thechain[1].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\thechain[2].chain1.ff[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\thechain[6].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\thechain[0].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\thechain[1].chain1.ff[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\thechain[1].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\thechain[4].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\thechain[4].chain1.ff[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\thechain[6].chain1.ff[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\thechain[7].chain1.ff[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\thechain[1].chain1.ff[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\thechain[5].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\thechain[4].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\thechain[5].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\thechain[2].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\thechain[5].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\thechain[3].chain1.ff[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\thechain[3].chain1.ff[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\thechain[0].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\thechain[7].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\thechain[3].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\thechain[4].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\thechain[0].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\thechain[1].chain1.ff[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\thechain[6].chain1.ff[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\thechain[4].chain1.ff[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\thechain[2].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\thechain[2].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\thechain[4].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\thechain[6].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\thechain[2].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\thechain[7].chain1.ff[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\thechain[1].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\thechain[0].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\thechain[4].chain1.ff[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\thechain[3].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\thechain[7].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\thechain[3].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\thechain[4].chain1.ff[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\thechain[0].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\thechain[1].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\thechain[3].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\thechain[4].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\thechain[7].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\thechain[5].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\thechain[5].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\thechain[3].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\thechain[1].chain1.ff[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\thechain[3].chain1.ff[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\thechain[2].chain1.ff[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\thechain[2].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\thechain[0].chain1.ff[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\thechain[5].chain1.ff[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\thechain[7].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\thechain[5].chain1.ff[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\thechain[0].chain1.ff[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\thechain[0].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\thechain[6].chain1.ff[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\thechain[4].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\thechain[3].chain1.ff[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\thechain[4].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\thechain[1].chain1.ff[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\thechain[6].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\thechain[4].chain1.ff[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\thechain[2].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\thechain[4].chain1.ff[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\thechain[2].chain1.ff[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\thechain[1].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\thechain[6].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\thechain[5].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\thechain[6].chain1.ff[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\thechain[0].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\thechain[6].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\thechain[4].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\thechain[4].chain1.ff[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\thechain[6].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\thechain[7].chain1.ff[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\thechain[3].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\thechain[3].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\thechain[2].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\thechain[6].chain1.ff[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\thechain[7].chain1.ff[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\thechain[7].chain1.ff[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\thechain[1].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\thechain[2].chain1.ff[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\thechain[4].chain1.ff[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\thechain[7].chain1.ff[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\thechain[5].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\thechain[2].chain1.ff[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\thechain[3].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\thechain[7].chain1.ff[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\thechain[7].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\thechain[1].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\thechain[2].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\thechain[4].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\thechain[0].chain1.ff[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\thechain[5].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\thechain[2].chain1.ff[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\thechain[1].chain1.ff[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\thechain[2].chain1.ff[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\thechain[3].chain1.ff[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\thechain[7].chain1.ff[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\thechain[1].chain1.ff[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\thechain[2].chain1.ff[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\thechain[5].chain1.ff[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\thechain[6].chain1.ff[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\thechain[3].chain1.ff[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\thechain[1].chain1.ff[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\thechain[7].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\thechain[6].chain1.ff[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\thechain[4].chain1.ff[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\thechain[0].chain1.ff[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\thechain[4].chain1.ff[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\thechain[6].chain1.ff[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\thechain[0].chain1.ff[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\thechain[3].chain1.ff[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\thechain[7].chain1.ff[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\thechain[7].chain1.ff[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\thechain[5].chain1.ff[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\thechain[7].chain1.ff[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\thechain[3].chain1.ff[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\thechain[7].chain1.ff[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\thechain[1].chain1.ff[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\thechain[0].chain1.ff[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\thechain[6].chain1.ff[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net738));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_3_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_5_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_163 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_6_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_206 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_95 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_10_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_23 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_11_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_12_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_15_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_24_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_116 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_29_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_123 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_30_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_30_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_212 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_36_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_41_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_43_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_172 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_43_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_45_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_47_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_50_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_50_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_51_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_52_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_52_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_95 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_53_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_57_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_60_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_63_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_65_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_65_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_67_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_68_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_69_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_69_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_71_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_71_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_72_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_72_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_73_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_73_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_74_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_74_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_74_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_75_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_75_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_75_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_76_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_76_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_76_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_76_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_76_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_120 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_77_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_77_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_77_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_80_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_80_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_80_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_80_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_201 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_80_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net91;
 assign uio_oe[1] = net92;
 assign uio_oe[2] = net93;
 assign uio_oe[3] = net94;
 assign uio_oe[4] = net95;
 assign uio_oe[5] = net96;
 assign uio_oe[6] = net97;
 assign uio_oe[7] = net98;
 assign uio_out[0] = net99;
 assign uio_out[1] = net100;
 assign uio_out[2] = net101;
 assign uio_out[3] = net102;
 assign uio_out[4] = net103;
 assign uio_out[5] = net104;
 assign uio_out[6] = net105;
 assign uio_out[7] = net106;
endmodule
