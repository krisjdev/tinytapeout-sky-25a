VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rejunity_atari2600
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_atari2600 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1378.160 BY 225.760 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 18.820 2.060 20.420 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.690 2.060 59.290 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.560 2.060 98.160 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.430 2.060 137.030 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.300 2.060 175.900 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.170 2.060 214.770 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 252.040 2.060 253.640 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.910 2.060 292.510 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.780 2.060 331.380 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.650 2.060 370.250 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 407.520 2.060 409.120 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.390 2.060 447.990 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.260 2.060 486.860 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.130 2.060 525.730 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.000 2.060 564.600 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.870 2.060 603.470 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 640.740 2.060 642.340 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.610 2.060 681.210 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 718.480 2.060 720.080 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 757.350 2.060 758.950 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.220 2.060 797.820 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 835.090 2.060 836.690 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.960 2.060 875.560 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 912.830 2.060 914.430 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.700 2.060 953.300 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 990.570 2.060 992.170 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1029.440 2.060 1031.040 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1068.310 2.060 1069.910 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.180 2.060 1108.780 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.050 2.060 1147.650 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.920 2.060 1186.520 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1262.660 2.060 1264.260 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.530 2.060 1303.130 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.400 2.060 1342.000 223.700 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.520 2.060 17.120 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.390 2.060 55.990 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.260 2.060 94.860 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.130 2.060 133.730 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.000 2.060 172.600 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.870 2.060 211.470 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.740 2.060 250.340 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 287.610 2.060 289.210 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.480 2.060 328.080 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 365.350 2.060 366.950 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.220 2.060 405.820 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.090 2.060 444.690 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.960 2.060 483.560 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 520.830 2.060 522.430 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 559.700 2.060 561.300 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 598.570 2.060 600.170 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 637.440 2.060 639.040 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.310 2.060 677.910 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 715.180 2.060 716.780 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 754.050 2.060 755.650 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.920 2.060 794.520 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.790 2.060 833.390 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 870.660 2.060 872.260 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.530 2.060 911.130 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 948.400 2.060 950.000 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 987.270 2.060 988.870 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.140 2.060 1027.740 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1065.010 2.060 1066.610 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.880 2.060 1105.480 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1142.750 2.060 1144.350 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1181.620 2.060 1183.220 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.360 2.060 1260.960 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1298.230 2.060 1299.830 223.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1337.100 2.060 1338.700 223.700 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.934000 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 1.650 0.330 1371.500 225.430 ;
      LAYER li1 ;
        RECT 1.840 0.450 1371.315 225.310 ;
      LAYER met1 ;
        RECT 1.840 0.040 1371.845 225.445 ;
      LAYER met2 ;
        RECT 7.920 0.010 1371.845 224.925 ;
      LAYER met3 ;
        RECT 12.945 0.315 1371.845 225.445 ;
      LAYER met4 ;
        RECT 31.370 224.360 33.030 224.905 ;
        RECT 34.130 224.360 35.790 224.905 ;
        RECT 36.890 224.360 38.550 224.905 ;
        RECT 39.650 224.360 41.310 224.905 ;
        RECT 42.410 224.360 44.070 224.905 ;
        RECT 45.170 224.360 46.830 224.905 ;
        RECT 47.930 224.360 49.590 224.905 ;
        RECT 50.690 224.360 52.350 224.905 ;
        RECT 53.450 224.360 55.110 224.905 ;
        RECT 56.210 224.360 57.870 224.905 ;
        RECT 58.970 224.360 60.630 224.905 ;
        RECT 61.730 224.360 63.390 224.905 ;
        RECT 64.490 224.360 66.150 224.905 ;
        RECT 67.250 224.360 68.910 224.905 ;
        RECT 70.010 224.360 71.670 224.905 ;
        RECT 72.770 224.360 74.430 224.905 ;
        RECT 75.530 224.360 77.190 224.905 ;
        RECT 78.290 224.360 79.950 224.905 ;
        RECT 81.050 224.360 82.710 224.905 ;
        RECT 83.810 224.360 85.470 224.905 ;
        RECT 86.570 224.360 88.230 224.905 ;
        RECT 89.330 224.360 90.990 224.905 ;
        RECT 92.090 224.360 93.750 224.905 ;
        RECT 94.850 224.360 96.510 224.905 ;
        RECT 97.610 224.360 99.270 224.905 ;
        RECT 100.370 224.360 102.030 224.905 ;
        RECT 103.130 224.360 104.790 224.905 ;
        RECT 105.890 224.360 107.550 224.905 ;
        RECT 108.650 224.360 110.310 224.905 ;
        RECT 111.410 224.360 113.070 224.905 ;
        RECT 114.170 224.360 115.830 224.905 ;
        RECT 116.930 224.360 118.590 224.905 ;
        RECT 119.690 224.360 121.350 224.905 ;
        RECT 122.450 224.360 124.110 224.905 ;
        RECT 125.210 224.360 126.870 224.905 ;
        RECT 127.970 224.360 129.630 224.905 ;
        RECT 130.730 224.360 132.390 224.905 ;
        RECT 133.490 224.360 135.150 224.905 ;
        RECT 136.250 224.360 137.910 224.905 ;
        RECT 139.010 224.360 140.670 224.905 ;
        RECT 141.770 224.360 143.430 224.905 ;
        RECT 144.530 224.360 146.190 224.905 ;
        RECT 147.290 224.360 1219.625 224.905 ;
        RECT 30.655 224.100 1219.625 224.360 ;
        RECT 30.655 6.295 53.990 224.100 ;
        RECT 56.390 6.295 57.290 224.100 ;
        RECT 59.690 6.295 92.860 224.100 ;
        RECT 95.260 6.295 96.160 224.100 ;
        RECT 98.560 6.295 131.730 224.100 ;
        RECT 134.130 6.295 135.030 224.100 ;
        RECT 137.430 6.295 170.600 224.100 ;
        RECT 173.000 6.295 173.900 224.100 ;
        RECT 176.300 6.295 209.470 224.100 ;
        RECT 211.870 6.295 212.770 224.100 ;
        RECT 215.170 6.295 248.340 224.100 ;
        RECT 250.740 6.295 251.640 224.100 ;
        RECT 254.040 6.295 287.210 224.100 ;
        RECT 289.610 6.295 290.510 224.100 ;
        RECT 292.910 6.295 326.080 224.100 ;
        RECT 328.480 6.295 329.380 224.100 ;
        RECT 331.780 6.295 364.950 224.100 ;
        RECT 367.350 6.295 368.250 224.100 ;
        RECT 370.650 6.295 403.820 224.100 ;
        RECT 406.220 6.295 407.120 224.100 ;
        RECT 409.520 6.295 442.690 224.100 ;
        RECT 445.090 6.295 445.990 224.100 ;
        RECT 448.390 6.295 481.560 224.100 ;
        RECT 483.960 6.295 484.860 224.100 ;
        RECT 487.260 6.295 520.430 224.100 ;
        RECT 522.830 6.295 523.730 224.100 ;
        RECT 526.130 6.295 559.300 224.100 ;
        RECT 561.700 6.295 562.600 224.100 ;
        RECT 565.000 6.295 598.170 224.100 ;
        RECT 600.570 6.295 601.470 224.100 ;
        RECT 603.870 6.295 637.040 224.100 ;
        RECT 639.440 6.295 640.340 224.100 ;
        RECT 642.740 6.295 675.910 224.100 ;
        RECT 678.310 6.295 679.210 224.100 ;
        RECT 681.610 6.295 714.780 224.100 ;
        RECT 717.180 6.295 718.080 224.100 ;
        RECT 720.480 6.295 753.650 224.100 ;
        RECT 756.050 6.295 756.950 224.100 ;
        RECT 759.350 6.295 792.520 224.100 ;
        RECT 794.920 6.295 795.820 224.100 ;
        RECT 798.220 6.295 831.390 224.100 ;
        RECT 833.790 6.295 834.690 224.100 ;
        RECT 837.090 6.295 870.260 224.100 ;
        RECT 872.660 6.295 873.560 224.100 ;
        RECT 875.960 6.295 909.130 224.100 ;
        RECT 911.530 6.295 912.430 224.100 ;
        RECT 914.830 6.295 948.000 224.100 ;
        RECT 950.400 6.295 951.300 224.100 ;
        RECT 953.700 6.295 986.870 224.100 ;
        RECT 989.270 6.295 990.170 224.100 ;
        RECT 992.570 6.295 1025.740 224.100 ;
        RECT 1028.140 6.295 1029.040 224.100 ;
        RECT 1031.440 6.295 1064.610 224.100 ;
        RECT 1067.010 6.295 1067.910 224.100 ;
        RECT 1070.310 6.295 1103.480 224.100 ;
        RECT 1105.880 6.295 1106.780 224.100 ;
        RECT 1109.180 6.295 1142.350 224.100 ;
        RECT 1144.750 6.295 1145.650 224.100 ;
        RECT 1148.050 6.295 1181.220 224.100 ;
        RECT 1183.620 6.295 1184.520 224.100 ;
        RECT 1186.920 6.295 1219.625 224.100 ;
  END
END tt_um_rejunity_atari2600
END LIBRARY

