VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_cw_vref
  CLASS BLOCK ;
  FOREIGN tt_um_cw_vref ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 4.640000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNADIFFAREA 4.640000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 320.000000 ;
    ANTENNADIFFAREA 9.280000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 12.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1134.794312 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 85.259995 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.600 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.600 5.000 5.200 220.760 ;
    END
  END VGND
  PIN VAPWR
    ANTENNAGATEAREA 2912.000000 ;
    ANTENNADIFFAREA 2005.394531 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.200 5.000 7.800 220.760 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 3.250 220.980 103.675 223.480 ;
        RECT 3.250 5.750 5.750 220.980 ;
        RECT 8.935 180.290 45.725 212.250 ;
        RECT 48.860 187.290 56.700 210.740 ;
      LAYER pwell ;
        RECT 9.140 168.330 52.250 178.810 ;
      LAYER nwell ;
        RECT 62.865 170.855 99.075 217.105 ;
        RECT 101.175 182.070 103.675 220.980 ;
        RECT 108.240 216.015 153.520 220.985 ;
        RECT 108.240 203.045 153.520 214.015 ;
      LAYER pwell ;
        RECT 108.440 184.690 153.320 201.100 ;
      LAYER nwell ;
        RECT 101.175 179.570 156.750 182.070 ;
      LAYER pwell ;
        RECT 9.140 147.810 51.970 168.220 ;
      LAYER nwell ;
        RECT 63.050 164.975 97.990 167.475 ;
      LAYER pwell ;
        RECT 9.600 134.835 20.550 138.315 ;
        RECT 23.425 135.385 58.475 143.515 ;
      LAYER nwell ;
        RECT 63.050 135.035 65.550 164.975 ;
        RECT 69.300 160.385 91.740 161.225 ;
        RECT 69.300 139.625 70.140 160.385 ;
      LAYER pwell ;
        RECT 71.090 158.670 89.950 159.435 ;
        RECT 71.090 156.220 71.855 158.670 ;
        RECT 74.305 156.220 75.575 158.670 ;
        RECT 78.025 156.220 79.295 158.670 ;
        RECT 81.745 156.220 83.015 158.670 ;
        RECT 85.465 156.220 86.735 158.670 ;
        RECT 89.185 156.220 89.950 158.670 ;
        RECT 71.090 154.950 89.950 156.220 ;
        RECT 71.090 152.500 71.855 154.950 ;
        RECT 74.305 152.500 75.575 154.950 ;
        RECT 78.025 152.500 79.295 154.950 ;
        RECT 81.745 152.500 83.015 154.950 ;
        RECT 85.465 152.500 86.735 154.950 ;
        RECT 89.185 152.500 89.950 154.950 ;
        RECT 71.090 151.230 89.950 152.500 ;
        RECT 71.090 148.780 71.855 151.230 ;
        RECT 74.305 148.780 75.575 151.230 ;
        RECT 78.025 148.780 79.295 151.230 ;
        RECT 81.745 148.780 83.015 151.230 ;
        RECT 85.465 148.780 86.735 151.230 ;
        RECT 89.185 148.780 89.950 151.230 ;
        RECT 71.090 147.510 89.950 148.780 ;
        RECT 71.090 145.060 71.855 147.510 ;
        RECT 74.305 145.060 75.575 147.510 ;
        RECT 78.025 145.060 79.295 147.510 ;
        RECT 81.745 145.060 83.015 147.510 ;
        RECT 85.465 145.060 86.735 147.510 ;
        RECT 89.185 145.060 89.950 147.510 ;
        RECT 71.090 143.790 89.950 145.060 ;
        RECT 71.090 141.340 71.855 143.790 ;
        RECT 74.305 141.340 75.575 143.790 ;
        RECT 78.025 141.340 79.295 143.790 ;
        RECT 81.745 141.340 83.015 143.790 ;
        RECT 85.465 141.340 86.735 143.790 ;
        RECT 89.185 141.340 89.950 143.790 ;
        RECT 71.090 140.575 89.950 141.340 ;
      LAYER nwell ;
        RECT 90.900 139.625 91.740 160.385 ;
        RECT 69.300 138.785 91.740 139.625 ;
        RECT 95.490 135.035 97.990 164.975 ;
      LAYER pwell ;
        RECT 102.550 158.280 111.160 172.690 ;
        RECT 114.030 166.235 151.540 176.715 ;
      LAYER nwell ;
        RECT 102.350 141.345 111.360 156.335 ;
        RECT 115.985 139.690 149.475 158.060 ;
        RECT 63.050 132.535 97.990 135.035 ;
        RECT 138.080 129.720 145.960 134.690 ;
      LAYER pwell ;
        RECT 138.280 124.290 145.760 128.770 ;
      LAYER nwell ;
        RECT 10.025 41.635 128.935 124.285 ;
      LAYER pwell ;
        RECT 10.225 9.090 74.495 39.430 ;
        RECT 79.865 9.090 128.735 39.430 ;
      LAYER nwell ;
        RECT 135.120 13.460 149.570 109.050 ;
        RECT 154.250 5.750 156.750 179.570 ;
        RECT 3.250 3.250 156.750 5.750 ;
      LAYER li1 ;
        RECT 4.300 222.030 102.625 222.430 ;
        RECT 4.300 4.700 4.700 222.030 ;
        RECT 62.895 216.545 99.045 217.075 ;
        RECT 62.895 213.695 63.425 216.545 ;
        RECT 63.925 215.855 80.385 216.025 ;
        RECT 63.925 214.385 64.155 215.855 ;
        RECT 80.155 214.385 80.385 215.855 ;
        RECT 63.925 214.215 80.385 214.385 ;
        RECT 80.885 213.695 81.055 216.545 ;
        RECT 81.555 215.855 98.015 216.025 ;
        RECT 81.555 214.385 81.785 215.855 ;
        RECT 97.785 214.385 98.015 215.855 ;
        RECT 81.555 214.215 98.015 214.385 ;
        RECT 98.515 213.695 99.045 216.545 ;
        RECT 62.895 213.525 99.045 213.695 ;
        RECT 9.325 211.690 45.335 211.860 ;
        RECT 9.325 201.840 9.495 211.690 ;
        RECT 10.225 211.000 18.225 211.170 ;
        RECT 18.515 211.000 26.515 211.170 ;
        RECT 9.995 202.745 10.165 210.785 ;
        RECT 18.285 202.745 18.455 210.785 ;
        RECT 26.575 202.745 26.745 210.785 ;
        RECT 10.225 202.360 18.225 202.530 ;
        RECT 18.515 202.360 26.515 202.530 ;
        RECT 27.245 201.840 27.415 211.690 ;
        RECT 28.145 211.000 36.145 211.170 ;
        RECT 36.435 211.000 44.435 211.170 ;
        RECT 27.915 202.745 28.085 210.785 ;
        RECT 36.205 202.745 36.375 210.785 ;
        RECT 44.495 202.745 44.665 210.785 ;
        RECT 28.145 202.360 36.145 202.530 ;
        RECT 36.435 202.360 44.435 202.530 ;
        RECT 45.165 201.840 45.335 211.690 ;
        RECT 62.895 210.675 63.425 213.525 ;
        RECT 64.155 212.835 80.155 213.005 ;
        RECT 63.925 211.580 64.095 212.620 ;
        RECT 80.215 211.580 80.385 212.620 ;
        RECT 64.155 211.195 80.155 211.365 ;
        RECT 80.885 210.675 81.055 213.525 ;
        RECT 81.785 212.835 97.785 213.005 ;
        RECT 81.555 211.580 81.725 212.620 ;
        RECT 97.845 211.580 98.015 212.620 ;
        RECT 81.785 211.195 97.785 211.365 ;
        RECT 98.515 210.675 99.045 213.525 ;
        RECT 62.895 210.505 99.045 210.675 ;
        RECT 9.325 201.670 45.335 201.840 ;
        RECT 9.325 191.820 9.495 201.670 ;
        RECT 10.225 200.980 18.225 201.150 ;
        RECT 18.515 200.980 26.515 201.150 ;
        RECT 9.995 192.725 10.165 200.765 ;
        RECT 18.285 192.725 18.455 200.765 ;
        RECT 26.575 192.725 26.745 200.765 ;
        RECT 10.225 192.340 18.225 192.510 ;
        RECT 18.515 192.340 26.515 192.510 ;
        RECT 27.245 191.820 27.415 201.670 ;
        RECT 28.145 200.980 36.145 201.150 ;
        RECT 36.435 200.980 44.435 201.150 ;
        RECT 27.915 192.725 28.085 200.765 ;
        RECT 36.205 192.725 36.375 200.765 ;
        RECT 44.495 192.725 44.665 200.765 ;
        RECT 28.145 192.340 36.145 192.510 ;
        RECT 36.435 192.340 44.435 192.510 ;
        RECT 45.165 191.820 45.335 201.670 ;
        RECT 9.325 191.650 45.335 191.820 ;
        RECT 49.250 210.180 56.310 210.350 ;
        RECT 9.325 190.700 15.415 190.870 ;
        RECT 9.325 180.850 9.495 190.700 ;
        RECT 10.225 190.010 12.225 190.180 ;
        RECT 12.515 190.010 14.515 190.180 ;
        RECT 9.995 181.755 10.165 189.795 ;
        RECT 12.285 181.755 12.455 189.795 ;
        RECT 14.575 181.755 14.745 189.795 ;
        RECT 10.225 181.370 12.225 181.540 ;
        RECT 12.515 181.370 14.515 181.540 ;
        RECT 15.245 180.850 15.415 190.700 ;
        RECT 9.325 180.680 15.415 180.850 ;
        RECT 16.345 190.700 45.335 190.870 ;
        RECT 16.345 180.850 16.515 190.700 ;
        RECT 17.245 190.010 19.245 190.180 ;
        RECT 19.535 190.010 21.535 190.180 ;
        RECT 21.825 190.010 23.825 190.180 ;
        RECT 24.115 190.010 26.115 190.180 ;
        RECT 26.405 190.010 28.405 190.180 ;
        RECT 28.695 190.010 30.695 190.180 ;
        RECT 30.985 190.010 32.985 190.180 ;
        RECT 33.275 190.010 35.275 190.180 ;
        RECT 35.565 190.010 37.565 190.180 ;
        RECT 37.855 190.010 39.855 190.180 ;
        RECT 40.145 190.010 42.145 190.180 ;
        RECT 42.435 190.010 44.435 190.180 ;
        RECT 17.015 181.755 17.185 189.795 ;
        RECT 19.305 181.755 19.475 189.795 ;
        RECT 21.595 181.755 21.765 189.795 ;
        RECT 23.885 181.755 24.055 189.795 ;
        RECT 26.175 181.755 26.345 189.795 ;
        RECT 28.465 181.755 28.635 189.795 ;
        RECT 30.755 181.755 30.925 189.795 ;
        RECT 33.045 181.755 33.215 189.795 ;
        RECT 35.335 181.755 35.505 189.795 ;
        RECT 37.625 181.755 37.795 189.795 ;
        RECT 39.915 181.755 40.085 189.795 ;
        RECT 42.205 181.755 42.375 189.795 ;
        RECT 44.495 181.755 44.665 189.795 ;
        RECT 17.245 181.370 19.245 181.540 ;
        RECT 19.535 181.370 21.535 181.540 ;
        RECT 21.825 181.370 23.825 181.540 ;
        RECT 24.115 181.370 26.115 181.540 ;
        RECT 26.405 181.370 28.405 181.540 ;
        RECT 28.695 181.370 30.695 181.540 ;
        RECT 30.985 181.370 32.985 181.540 ;
        RECT 33.275 181.370 35.275 181.540 ;
        RECT 35.565 181.370 37.565 181.540 ;
        RECT 37.855 181.370 39.855 181.540 ;
        RECT 40.145 181.370 42.145 181.540 ;
        RECT 42.435 181.370 44.435 181.540 ;
        RECT 45.165 180.850 45.335 190.700 ;
        RECT 49.250 187.850 49.420 210.180 ;
        RECT 50.095 207.435 50.785 209.595 ;
        RECT 51.265 207.435 51.955 209.595 ;
        RECT 52.435 207.435 53.125 209.595 ;
        RECT 53.605 207.435 54.295 209.595 ;
        RECT 54.775 207.435 55.465 209.595 ;
        RECT 50.095 188.435 50.785 190.595 ;
        RECT 51.265 188.435 51.955 190.595 ;
        RECT 52.435 188.435 53.125 190.595 ;
        RECT 53.605 188.435 54.295 190.595 ;
        RECT 54.775 188.435 55.465 190.595 ;
        RECT 56.140 187.850 56.310 210.180 ;
        RECT 49.250 187.680 56.310 187.850 ;
        RECT 62.895 207.655 63.425 210.505 ;
        RECT 64.155 209.815 80.155 209.985 ;
        RECT 63.925 208.560 64.095 209.600 ;
        RECT 80.215 208.560 80.385 209.600 ;
        RECT 64.155 208.175 80.155 208.345 ;
        RECT 80.885 207.655 81.055 210.505 ;
        RECT 81.785 209.815 97.785 209.985 ;
        RECT 81.555 208.560 81.725 209.600 ;
        RECT 97.845 208.560 98.015 209.600 ;
        RECT 81.785 208.175 97.785 208.345 ;
        RECT 98.515 207.655 99.045 210.505 ;
        RECT 62.895 207.485 99.045 207.655 ;
        RECT 62.895 204.635 63.425 207.485 ;
        RECT 64.155 206.795 80.155 206.965 ;
        RECT 63.925 205.540 64.095 206.580 ;
        RECT 80.215 205.540 80.385 206.580 ;
        RECT 64.155 205.155 80.155 205.325 ;
        RECT 80.885 204.635 81.055 207.485 ;
        RECT 81.785 206.795 97.785 206.965 ;
        RECT 81.555 205.540 81.725 206.580 ;
        RECT 97.845 205.540 98.015 206.580 ;
        RECT 81.785 205.155 97.785 205.325 ;
        RECT 98.515 204.635 99.045 207.485 ;
        RECT 62.895 204.465 99.045 204.635 ;
        RECT 62.895 201.615 63.425 204.465 ;
        RECT 64.155 203.775 80.155 203.945 ;
        RECT 63.925 202.520 64.095 203.560 ;
        RECT 80.215 202.520 80.385 203.560 ;
        RECT 64.155 202.135 80.155 202.305 ;
        RECT 80.885 201.615 81.055 204.465 ;
        RECT 81.785 203.775 97.785 203.945 ;
        RECT 81.555 202.520 81.725 203.560 ;
        RECT 97.845 202.520 98.015 203.560 ;
        RECT 81.785 202.135 97.785 202.305 ;
        RECT 98.515 201.615 99.045 204.465 ;
        RECT 62.895 201.445 99.045 201.615 ;
        RECT 62.895 198.595 63.425 201.445 ;
        RECT 64.155 200.755 80.155 200.925 ;
        RECT 63.925 199.500 64.095 200.540 ;
        RECT 80.215 199.500 80.385 200.540 ;
        RECT 64.155 199.115 80.155 199.285 ;
        RECT 80.885 198.595 81.055 201.445 ;
        RECT 81.785 200.755 97.785 200.925 ;
        RECT 81.555 199.500 81.725 200.540 ;
        RECT 97.845 199.500 98.015 200.540 ;
        RECT 81.785 199.115 97.785 199.285 ;
        RECT 98.515 198.595 99.045 201.445 ;
        RECT 62.895 198.425 99.045 198.595 ;
        RECT 62.895 195.575 63.425 198.425 ;
        RECT 64.155 197.735 80.155 197.905 ;
        RECT 63.925 196.480 64.095 197.520 ;
        RECT 80.215 196.480 80.385 197.520 ;
        RECT 64.155 196.095 80.155 196.265 ;
        RECT 80.885 195.575 81.055 198.425 ;
        RECT 81.785 197.735 97.785 197.905 ;
        RECT 81.555 196.480 81.725 197.520 ;
        RECT 97.845 196.480 98.015 197.520 ;
        RECT 81.785 196.095 97.785 196.265 ;
        RECT 98.515 195.575 99.045 198.425 ;
        RECT 62.895 195.405 99.045 195.575 ;
        RECT 62.895 192.555 63.425 195.405 ;
        RECT 64.155 194.715 80.155 194.885 ;
        RECT 63.925 193.460 64.095 194.500 ;
        RECT 80.215 193.460 80.385 194.500 ;
        RECT 64.155 193.075 80.155 193.245 ;
        RECT 80.885 192.555 81.055 195.405 ;
        RECT 81.785 194.715 97.785 194.885 ;
        RECT 81.555 193.460 81.725 194.500 ;
        RECT 97.845 193.460 98.015 194.500 ;
        RECT 81.785 193.075 97.785 193.245 ;
        RECT 98.515 192.555 99.045 195.405 ;
        RECT 62.895 192.385 99.045 192.555 ;
        RECT 62.895 189.535 63.425 192.385 ;
        RECT 64.155 191.695 80.155 191.865 ;
        RECT 63.925 190.440 64.095 191.480 ;
        RECT 80.215 190.440 80.385 191.480 ;
        RECT 64.155 190.055 80.155 190.225 ;
        RECT 80.885 189.535 81.055 192.385 ;
        RECT 81.785 191.695 97.785 191.865 ;
        RECT 81.555 190.440 81.725 191.480 ;
        RECT 97.845 190.440 98.015 191.480 ;
        RECT 81.785 190.055 97.785 190.225 ;
        RECT 98.515 189.535 99.045 192.385 ;
        RECT 62.895 189.365 99.045 189.535 ;
        RECT 16.345 180.680 45.335 180.850 ;
        RECT 62.895 186.515 63.425 189.365 ;
        RECT 64.155 188.675 80.155 188.845 ;
        RECT 63.925 187.420 64.095 188.460 ;
        RECT 80.215 187.420 80.385 188.460 ;
        RECT 64.155 187.035 80.155 187.205 ;
        RECT 80.885 186.515 81.055 189.365 ;
        RECT 81.785 188.675 97.785 188.845 ;
        RECT 81.555 187.420 81.725 188.460 ;
        RECT 97.845 187.420 98.015 188.460 ;
        RECT 81.785 187.035 97.785 187.205 ;
        RECT 98.515 186.515 99.045 189.365 ;
        RECT 62.895 186.345 99.045 186.515 ;
        RECT 62.895 183.495 63.425 186.345 ;
        RECT 64.155 185.655 80.155 185.825 ;
        RECT 63.925 184.400 64.095 185.440 ;
        RECT 80.215 184.400 80.385 185.440 ;
        RECT 64.155 184.015 80.155 184.185 ;
        RECT 80.885 183.495 81.055 186.345 ;
        RECT 81.785 185.655 97.785 185.825 ;
        RECT 81.555 184.400 81.725 185.440 ;
        RECT 97.845 184.400 98.015 185.440 ;
        RECT 81.785 184.015 97.785 184.185 ;
        RECT 98.515 183.495 99.045 186.345 ;
        RECT 62.895 183.325 99.045 183.495 ;
        RECT 62.895 180.475 63.425 183.325 ;
        RECT 64.155 182.635 80.155 182.805 ;
        RECT 63.925 181.380 64.095 182.420 ;
        RECT 80.215 181.380 80.385 182.420 ;
        RECT 64.155 180.995 80.155 181.165 ;
        RECT 80.885 180.475 81.055 183.325 ;
        RECT 81.785 182.635 97.785 182.805 ;
        RECT 81.555 181.380 81.725 182.420 ;
        RECT 97.845 181.380 98.015 182.420 ;
        RECT 81.785 180.995 97.785 181.165 ;
        RECT 98.515 180.475 99.045 183.325 ;
        RECT 102.225 181.020 102.625 222.030 ;
        RECT 108.630 220.425 153.130 220.595 ;
        RECT 108.630 216.575 108.800 220.425 ;
        RECT 109.585 219.735 110.585 219.905 ;
        RECT 110.875 219.735 111.875 219.905 ;
        RECT 109.355 217.480 109.525 219.520 ;
        RECT 110.645 217.480 110.815 219.520 ;
        RECT 111.935 217.480 112.105 219.520 ;
        RECT 109.585 217.095 110.585 217.265 ;
        RECT 110.875 217.095 111.875 217.265 ;
        RECT 112.660 216.575 112.830 220.425 ;
        RECT 113.615 219.735 114.615 219.905 ;
        RECT 114.905 219.735 115.905 219.905 ;
        RECT 113.385 217.480 113.555 219.520 ;
        RECT 114.675 217.480 114.845 219.520 ;
        RECT 115.965 217.480 116.135 219.520 ;
        RECT 113.615 217.095 114.615 217.265 ;
        RECT 114.905 217.095 115.905 217.265 ;
        RECT 116.690 216.575 116.860 220.425 ;
        RECT 117.645 219.735 118.645 219.905 ;
        RECT 118.935 219.735 119.935 219.905 ;
        RECT 117.415 217.480 117.585 219.520 ;
        RECT 118.705 217.480 118.875 219.520 ;
        RECT 119.995 217.480 120.165 219.520 ;
        RECT 117.645 217.095 118.645 217.265 ;
        RECT 118.935 217.095 119.935 217.265 ;
        RECT 120.720 216.575 120.890 220.425 ;
        RECT 121.675 219.735 122.675 219.905 ;
        RECT 122.965 219.735 123.965 219.905 ;
        RECT 121.445 217.480 121.615 219.520 ;
        RECT 122.735 217.480 122.905 219.520 ;
        RECT 124.025 217.480 124.195 219.520 ;
        RECT 121.675 217.095 122.675 217.265 ;
        RECT 122.965 217.095 123.965 217.265 ;
        RECT 124.750 216.575 124.920 220.425 ;
        RECT 125.705 219.735 126.705 219.905 ;
        RECT 126.995 219.735 127.995 219.905 ;
        RECT 125.475 217.480 125.645 219.520 ;
        RECT 126.765 217.480 126.935 219.520 ;
        RECT 128.055 217.480 128.225 219.520 ;
        RECT 125.705 217.095 126.705 217.265 ;
        RECT 126.995 217.095 127.995 217.265 ;
        RECT 128.780 216.575 128.950 220.425 ;
        RECT 129.735 219.735 130.735 219.905 ;
        RECT 131.025 219.735 132.025 219.905 ;
        RECT 129.505 217.480 129.675 219.520 ;
        RECT 130.795 217.480 130.965 219.520 ;
        RECT 132.085 217.480 132.255 219.520 ;
        RECT 129.735 217.095 130.735 217.265 ;
        RECT 131.025 217.095 132.025 217.265 ;
        RECT 132.810 216.575 132.980 220.425 ;
        RECT 133.765 219.735 134.765 219.905 ;
        RECT 135.055 219.735 136.055 219.905 ;
        RECT 133.535 217.480 133.705 219.520 ;
        RECT 134.825 217.480 134.995 219.520 ;
        RECT 136.115 217.480 136.285 219.520 ;
        RECT 133.765 217.095 134.765 217.265 ;
        RECT 135.055 217.095 136.055 217.265 ;
        RECT 136.840 216.575 137.010 220.425 ;
        RECT 137.795 219.735 138.795 219.905 ;
        RECT 139.085 219.735 140.085 219.905 ;
        RECT 137.565 217.480 137.735 219.520 ;
        RECT 138.855 217.480 139.025 219.520 ;
        RECT 140.145 217.480 140.315 219.520 ;
        RECT 137.795 217.095 138.795 217.265 ;
        RECT 139.085 217.095 140.085 217.265 ;
        RECT 140.870 216.575 141.040 220.425 ;
        RECT 141.825 219.735 142.825 219.905 ;
        RECT 143.115 219.735 144.115 219.905 ;
        RECT 141.595 217.480 141.765 219.520 ;
        RECT 142.885 217.480 143.055 219.520 ;
        RECT 144.175 217.480 144.345 219.520 ;
        RECT 141.825 217.095 142.825 217.265 ;
        RECT 143.115 217.095 144.115 217.265 ;
        RECT 144.900 216.575 145.070 220.425 ;
        RECT 145.855 219.735 146.855 219.905 ;
        RECT 147.145 219.735 148.145 219.905 ;
        RECT 145.625 217.480 145.795 219.520 ;
        RECT 146.915 217.480 147.085 219.520 ;
        RECT 148.205 217.480 148.375 219.520 ;
        RECT 145.855 217.095 146.855 217.265 ;
        RECT 147.145 217.095 148.145 217.265 ;
        RECT 148.930 216.575 149.100 220.425 ;
        RECT 149.885 219.735 150.885 219.905 ;
        RECT 151.175 219.735 152.175 219.905 ;
        RECT 149.655 217.480 149.825 219.520 ;
        RECT 150.945 217.480 151.115 219.520 ;
        RECT 152.235 217.480 152.405 219.520 ;
        RECT 149.885 217.095 150.885 217.265 ;
        RECT 151.175 217.095 152.175 217.265 ;
        RECT 152.960 216.575 153.130 220.425 ;
        RECT 108.630 216.405 153.130 216.575 ;
        RECT 108.630 213.455 153.130 213.625 ;
        RECT 108.630 203.605 108.800 213.455 ;
        RECT 109.585 212.765 110.585 212.935 ;
        RECT 110.875 212.765 111.875 212.935 ;
        RECT 109.355 204.510 109.525 212.550 ;
        RECT 110.645 204.510 110.815 212.550 ;
        RECT 111.935 204.510 112.105 212.550 ;
        RECT 109.585 204.125 110.585 204.295 ;
        RECT 110.875 204.125 111.875 204.295 ;
        RECT 112.660 203.605 112.830 213.455 ;
        RECT 113.615 212.765 114.615 212.935 ;
        RECT 114.905 212.765 115.905 212.935 ;
        RECT 113.385 204.510 113.555 212.550 ;
        RECT 114.675 204.510 114.845 212.550 ;
        RECT 115.965 204.510 116.135 212.550 ;
        RECT 113.615 204.125 114.615 204.295 ;
        RECT 114.905 204.125 115.905 204.295 ;
        RECT 116.690 203.605 116.860 213.455 ;
        RECT 117.645 212.765 118.645 212.935 ;
        RECT 118.935 212.765 119.935 212.935 ;
        RECT 117.415 204.510 117.585 212.550 ;
        RECT 118.705 204.510 118.875 212.550 ;
        RECT 119.995 204.510 120.165 212.550 ;
        RECT 117.645 204.125 118.645 204.295 ;
        RECT 118.935 204.125 119.935 204.295 ;
        RECT 120.720 203.605 120.890 213.455 ;
        RECT 121.675 212.765 122.675 212.935 ;
        RECT 122.965 212.765 123.965 212.935 ;
        RECT 121.445 204.510 121.615 212.550 ;
        RECT 122.735 204.510 122.905 212.550 ;
        RECT 124.025 204.510 124.195 212.550 ;
        RECT 121.675 204.125 122.675 204.295 ;
        RECT 122.965 204.125 123.965 204.295 ;
        RECT 124.750 203.605 124.920 213.455 ;
        RECT 125.705 212.765 126.705 212.935 ;
        RECT 126.995 212.765 127.995 212.935 ;
        RECT 125.475 204.510 125.645 212.550 ;
        RECT 126.765 204.510 126.935 212.550 ;
        RECT 128.055 204.510 128.225 212.550 ;
        RECT 125.705 204.125 126.705 204.295 ;
        RECT 126.995 204.125 127.995 204.295 ;
        RECT 128.780 203.605 128.950 213.455 ;
        RECT 129.735 212.765 130.735 212.935 ;
        RECT 131.025 212.765 132.025 212.935 ;
        RECT 129.505 204.510 129.675 212.550 ;
        RECT 130.795 204.510 130.965 212.550 ;
        RECT 132.085 204.510 132.255 212.550 ;
        RECT 129.735 204.125 130.735 204.295 ;
        RECT 131.025 204.125 132.025 204.295 ;
        RECT 132.810 203.605 132.980 213.455 ;
        RECT 133.765 212.765 134.765 212.935 ;
        RECT 135.055 212.765 136.055 212.935 ;
        RECT 133.535 204.510 133.705 212.550 ;
        RECT 134.825 204.510 134.995 212.550 ;
        RECT 136.115 204.510 136.285 212.550 ;
        RECT 133.765 204.125 134.765 204.295 ;
        RECT 135.055 204.125 136.055 204.295 ;
        RECT 136.840 203.605 137.010 213.455 ;
        RECT 137.795 212.765 138.795 212.935 ;
        RECT 139.085 212.765 140.085 212.935 ;
        RECT 137.565 204.510 137.735 212.550 ;
        RECT 138.855 204.510 139.025 212.550 ;
        RECT 140.145 204.510 140.315 212.550 ;
        RECT 137.795 204.125 138.795 204.295 ;
        RECT 139.085 204.125 140.085 204.295 ;
        RECT 140.870 203.605 141.040 213.455 ;
        RECT 141.825 212.765 142.825 212.935 ;
        RECT 143.115 212.765 144.115 212.935 ;
        RECT 141.595 204.510 141.765 212.550 ;
        RECT 142.885 204.510 143.055 212.550 ;
        RECT 144.175 204.510 144.345 212.550 ;
        RECT 141.825 204.125 142.825 204.295 ;
        RECT 143.115 204.125 144.115 204.295 ;
        RECT 144.900 203.605 145.070 213.455 ;
        RECT 145.855 212.765 146.855 212.935 ;
        RECT 147.145 212.765 148.145 212.935 ;
        RECT 145.625 204.510 145.795 212.550 ;
        RECT 146.915 204.510 147.085 212.550 ;
        RECT 148.205 204.510 148.375 212.550 ;
        RECT 145.855 204.125 146.855 204.295 ;
        RECT 147.145 204.125 148.145 204.295 ;
        RECT 148.930 203.605 149.100 213.455 ;
        RECT 149.885 212.765 150.885 212.935 ;
        RECT 151.175 212.765 152.175 212.935 ;
        RECT 149.655 204.510 149.825 212.550 ;
        RECT 150.945 204.510 151.115 212.550 ;
        RECT 152.235 204.510 152.405 212.550 ;
        RECT 149.885 204.125 150.885 204.295 ;
        RECT 151.175 204.125 152.175 204.295 ;
        RECT 152.960 203.605 153.130 213.455 ;
        RECT 108.630 203.435 153.130 203.605 ;
        RECT 108.630 200.740 153.130 200.910 ;
        RECT 108.630 194.980 108.800 200.740 ;
        RECT 109.585 200.050 110.585 200.220 ;
        RECT 110.875 200.050 111.875 200.220 ;
        RECT 109.355 195.840 109.525 199.880 ;
        RECT 110.645 195.840 110.815 199.880 ;
        RECT 111.935 195.840 112.105 199.880 ;
        RECT 109.585 195.500 110.585 195.670 ;
        RECT 110.875 195.500 111.875 195.670 ;
        RECT 112.660 194.980 112.830 200.740 ;
        RECT 113.615 200.050 114.615 200.220 ;
        RECT 114.905 200.050 115.905 200.220 ;
        RECT 113.385 195.840 113.555 199.880 ;
        RECT 114.675 195.840 114.845 199.880 ;
        RECT 115.965 195.840 116.135 199.880 ;
        RECT 113.615 195.500 114.615 195.670 ;
        RECT 114.905 195.500 115.905 195.670 ;
        RECT 116.690 194.980 116.860 200.740 ;
        RECT 117.645 200.050 118.645 200.220 ;
        RECT 118.935 200.050 119.935 200.220 ;
        RECT 117.415 195.840 117.585 199.880 ;
        RECT 118.705 195.840 118.875 199.880 ;
        RECT 119.995 195.840 120.165 199.880 ;
        RECT 117.645 195.500 118.645 195.670 ;
        RECT 118.935 195.500 119.935 195.670 ;
        RECT 120.720 194.980 120.890 200.740 ;
        RECT 121.675 200.050 122.675 200.220 ;
        RECT 122.965 200.050 123.965 200.220 ;
        RECT 121.445 195.840 121.615 199.880 ;
        RECT 122.735 195.840 122.905 199.880 ;
        RECT 124.025 195.840 124.195 199.880 ;
        RECT 121.675 195.500 122.675 195.670 ;
        RECT 122.965 195.500 123.965 195.670 ;
        RECT 124.750 194.980 124.920 200.740 ;
        RECT 125.705 200.050 126.705 200.220 ;
        RECT 126.995 200.050 127.995 200.220 ;
        RECT 125.475 195.840 125.645 199.880 ;
        RECT 126.765 195.840 126.935 199.880 ;
        RECT 128.055 195.840 128.225 199.880 ;
        RECT 125.705 195.500 126.705 195.670 ;
        RECT 126.995 195.500 127.995 195.670 ;
        RECT 128.780 194.980 128.950 200.740 ;
        RECT 129.735 200.050 130.735 200.220 ;
        RECT 131.025 200.050 132.025 200.220 ;
        RECT 129.505 195.840 129.675 199.880 ;
        RECT 130.795 195.840 130.965 199.880 ;
        RECT 132.085 195.840 132.255 199.880 ;
        RECT 129.735 195.500 130.735 195.670 ;
        RECT 131.025 195.500 132.025 195.670 ;
        RECT 132.810 194.980 132.980 200.740 ;
        RECT 133.765 200.050 134.765 200.220 ;
        RECT 135.055 200.050 136.055 200.220 ;
        RECT 133.535 195.840 133.705 199.880 ;
        RECT 134.825 195.840 134.995 199.880 ;
        RECT 136.115 195.840 136.285 199.880 ;
        RECT 133.765 195.500 134.765 195.670 ;
        RECT 135.055 195.500 136.055 195.670 ;
        RECT 136.840 194.980 137.010 200.740 ;
        RECT 137.795 200.050 138.795 200.220 ;
        RECT 139.085 200.050 140.085 200.220 ;
        RECT 137.565 195.840 137.735 199.880 ;
        RECT 138.855 195.840 139.025 199.880 ;
        RECT 140.145 195.840 140.315 199.880 ;
        RECT 137.795 195.500 138.795 195.670 ;
        RECT 139.085 195.500 140.085 195.670 ;
        RECT 140.870 194.980 141.040 200.740 ;
        RECT 141.825 200.050 142.825 200.220 ;
        RECT 143.115 200.050 144.115 200.220 ;
        RECT 141.595 195.840 141.765 199.880 ;
        RECT 142.885 195.840 143.055 199.880 ;
        RECT 144.175 195.840 144.345 199.880 ;
        RECT 141.825 195.500 142.825 195.670 ;
        RECT 143.115 195.500 144.115 195.670 ;
        RECT 144.900 194.980 145.070 200.740 ;
        RECT 145.855 200.050 146.855 200.220 ;
        RECT 147.145 200.050 148.145 200.220 ;
        RECT 145.625 195.840 145.795 199.880 ;
        RECT 146.915 195.840 147.085 199.880 ;
        RECT 148.205 195.840 148.375 199.880 ;
        RECT 145.855 195.500 146.855 195.670 ;
        RECT 147.145 195.500 148.145 195.670 ;
        RECT 148.930 194.980 149.100 200.740 ;
        RECT 149.885 200.050 150.885 200.220 ;
        RECT 151.175 200.050 152.175 200.220 ;
        RECT 149.655 195.840 149.825 199.880 ;
        RECT 150.945 195.840 151.115 199.880 ;
        RECT 152.235 195.840 152.405 199.880 ;
        RECT 149.885 195.500 150.885 195.670 ;
        RECT 151.175 195.500 152.175 195.670 ;
        RECT 152.960 194.980 153.130 200.740 ;
        RECT 108.630 194.810 153.130 194.980 ;
        RECT 108.630 185.050 108.800 194.810 ;
        RECT 109.585 194.120 110.585 194.290 ;
        RECT 110.875 194.120 111.875 194.290 ;
        RECT 109.355 185.910 109.525 193.950 ;
        RECT 110.645 185.910 110.815 193.950 ;
        RECT 111.935 185.910 112.105 193.950 ;
        RECT 109.585 185.570 110.585 185.740 ;
        RECT 110.875 185.570 111.875 185.740 ;
        RECT 112.660 185.050 112.830 194.810 ;
        RECT 113.615 194.120 114.615 194.290 ;
        RECT 114.905 194.120 115.905 194.290 ;
        RECT 113.385 185.910 113.555 193.950 ;
        RECT 114.675 185.910 114.845 193.950 ;
        RECT 115.965 185.910 116.135 193.950 ;
        RECT 113.615 185.570 114.615 185.740 ;
        RECT 114.905 185.570 115.905 185.740 ;
        RECT 116.690 185.050 116.860 194.810 ;
        RECT 117.645 194.120 118.645 194.290 ;
        RECT 118.935 194.120 119.935 194.290 ;
        RECT 117.415 185.910 117.585 193.950 ;
        RECT 118.705 185.910 118.875 193.950 ;
        RECT 119.995 185.910 120.165 193.950 ;
        RECT 117.645 185.570 118.645 185.740 ;
        RECT 118.935 185.570 119.935 185.740 ;
        RECT 120.720 185.050 120.890 194.810 ;
        RECT 121.675 194.120 122.675 194.290 ;
        RECT 122.965 194.120 123.965 194.290 ;
        RECT 121.445 185.910 121.615 193.950 ;
        RECT 122.735 185.910 122.905 193.950 ;
        RECT 124.025 185.910 124.195 193.950 ;
        RECT 121.675 185.570 122.675 185.740 ;
        RECT 122.965 185.570 123.965 185.740 ;
        RECT 124.750 185.050 124.920 194.810 ;
        RECT 125.705 194.120 126.705 194.290 ;
        RECT 126.995 194.120 127.995 194.290 ;
        RECT 125.475 185.910 125.645 193.950 ;
        RECT 126.765 185.910 126.935 193.950 ;
        RECT 128.055 185.910 128.225 193.950 ;
        RECT 125.705 185.570 126.705 185.740 ;
        RECT 126.995 185.570 127.995 185.740 ;
        RECT 128.780 185.050 128.950 194.810 ;
        RECT 129.735 194.120 130.735 194.290 ;
        RECT 131.025 194.120 132.025 194.290 ;
        RECT 129.505 185.910 129.675 193.950 ;
        RECT 130.795 185.910 130.965 193.950 ;
        RECT 132.085 185.910 132.255 193.950 ;
        RECT 129.735 185.570 130.735 185.740 ;
        RECT 131.025 185.570 132.025 185.740 ;
        RECT 132.810 185.050 132.980 194.810 ;
        RECT 133.765 194.120 134.765 194.290 ;
        RECT 135.055 194.120 136.055 194.290 ;
        RECT 133.535 185.910 133.705 193.950 ;
        RECT 134.825 185.910 134.995 193.950 ;
        RECT 136.115 185.910 136.285 193.950 ;
        RECT 133.765 185.570 134.765 185.740 ;
        RECT 135.055 185.570 136.055 185.740 ;
        RECT 136.840 185.050 137.010 194.810 ;
        RECT 137.795 194.120 138.795 194.290 ;
        RECT 139.085 194.120 140.085 194.290 ;
        RECT 137.565 185.910 137.735 193.950 ;
        RECT 138.855 185.910 139.025 193.950 ;
        RECT 140.145 185.910 140.315 193.950 ;
        RECT 137.795 185.570 138.795 185.740 ;
        RECT 139.085 185.570 140.085 185.740 ;
        RECT 140.870 185.050 141.040 194.810 ;
        RECT 141.825 194.120 142.825 194.290 ;
        RECT 143.115 194.120 144.115 194.290 ;
        RECT 141.595 185.910 141.765 193.950 ;
        RECT 142.885 185.910 143.055 193.950 ;
        RECT 144.175 185.910 144.345 193.950 ;
        RECT 141.825 185.570 142.825 185.740 ;
        RECT 143.115 185.570 144.115 185.740 ;
        RECT 144.900 185.050 145.070 194.810 ;
        RECT 145.855 194.120 146.855 194.290 ;
        RECT 147.145 194.120 148.145 194.290 ;
        RECT 145.625 185.910 145.795 193.950 ;
        RECT 146.915 185.910 147.085 193.950 ;
        RECT 148.205 185.910 148.375 193.950 ;
        RECT 145.855 185.570 146.855 185.740 ;
        RECT 147.145 185.570 148.145 185.740 ;
        RECT 148.930 185.050 149.100 194.810 ;
        RECT 149.885 194.120 150.885 194.290 ;
        RECT 151.175 194.120 152.175 194.290 ;
        RECT 149.655 185.910 149.825 193.950 ;
        RECT 150.945 185.910 151.115 193.950 ;
        RECT 152.235 185.910 152.405 193.950 ;
        RECT 149.885 185.570 150.885 185.740 ;
        RECT 151.175 185.570 152.175 185.740 ;
        RECT 152.960 185.050 153.130 194.810 ;
        RECT 108.630 184.880 153.130 185.050 ;
        RECT 102.225 180.620 155.700 181.020 ;
        RECT 62.895 180.305 99.045 180.475 ;
        RECT 9.330 178.450 52.060 178.620 ;
        RECT 9.330 168.690 9.500 178.450 ;
        RECT 10.230 177.760 12.230 177.930 ;
        RECT 12.520 177.760 14.520 177.930 ;
        RECT 14.810 177.760 16.810 177.930 ;
        RECT 17.100 177.760 19.100 177.930 ;
        RECT 19.390 177.760 21.390 177.930 ;
        RECT 21.680 177.760 23.680 177.930 ;
        RECT 23.970 177.760 25.970 177.930 ;
        RECT 26.260 177.760 28.260 177.930 ;
        RECT 28.550 177.760 30.550 177.930 ;
        RECT 30.840 177.760 32.840 177.930 ;
        RECT 33.130 177.760 35.130 177.930 ;
        RECT 35.420 177.760 37.420 177.930 ;
        RECT 37.710 177.760 39.710 177.930 ;
        RECT 40.000 177.760 42.000 177.930 ;
        RECT 42.290 177.760 44.290 177.930 ;
        RECT 44.580 177.760 46.580 177.930 ;
        RECT 46.870 177.760 48.870 177.930 ;
        RECT 49.160 177.760 51.160 177.930 ;
        RECT 10.000 169.550 10.170 177.590 ;
        RECT 12.290 169.550 12.460 177.590 ;
        RECT 14.580 169.550 14.750 177.590 ;
        RECT 16.870 169.550 17.040 177.590 ;
        RECT 19.160 169.550 19.330 177.590 ;
        RECT 21.450 169.550 21.620 177.590 ;
        RECT 23.740 169.550 23.910 177.590 ;
        RECT 26.030 169.550 26.200 177.590 ;
        RECT 28.320 169.550 28.490 177.590 ;
        RECT 30.610 169.550 30.780 177.590 ;
        RECT 32.900 169.550 33.070 177.590 ;
        RECT 35.190 169.550 35.360 177.590 ;
        RECT 37.480 169.550 37.650 177.590 ;
        RECT 39.770 169.550 39.940 177.590 ;
        RECT 42.060 169.550 42.230 177.590 ;
        RECT 44.350 169.550 44.520 177.590 ;
        RECT 46.640 169.550 46.810 177.590 ;
        RECT 48.930 169.550 49.100 177.590 ;
        RECT 51.220 169.550 51.390 177.590 ;
        RECT 10.230 169.210 12.230 169.380 ;
        RECT 12.520 169.210 14.520 169.380 ;
        RECT 14.810 169.210 16.810 169.380 ;
        RECT 17.100 169.210 19.100 169.380 ;
        RECT 19.390 169.210 21.390 169.380 ;
        RECT 21.680 169.210 23.680 169.380 ;
        RECT 23.970 169.210 25.970 169.380 ;
        RECT 26.260 169.210 28.260 169.380 ;
        RECT 28.550 169.210 30.550 169.380 ;
        RECT 30.840 169.210 32.840 169.380 ;
        RECT 33.130 169.210 35.130 169.380 ;
        RECT 35.420 169.210 37.420 169.380 ;
        RECT 37.710 169.210 39.710 169.380 ;
        RECT 40.000 169.210 42.000 169.380 ;
        RECT 42.290 169.210 44.290 169.380 ;
        RECT 44.580 169.210 46.580 169.380 ;
        RECT 46.870 169.210 48.870 169.380 ;
        RECT 49.160 169.210 51.160 169.380 ;
        RECT 51.890 168.690 52.060 178.450 ;
        RECT 62.895 177.455 63.425 180.305 ;
        RECT 64.155 179.615 80.155 179.785 ;
        RECT 63.925 178.360 64.095 179.400 ;
        RECT 80.215 178.360 80.385 179.400 ;
        RECT 64.155 177.975 80.155 178.145 ;
        RECT 80.885 177.455 81.055 180.305 ;
        RECT 81.785 179.615 97.785 179.785 ;
        RECT 81.555 178.360 81.725 179.400 ;
        RECT 97.845 178.360 98.015 179.400 ;
        RECT 81.785 177.975 97.785 178.145 ;
        RECT 98.515 177.455 99.045 180.305 ;
        RECT 62.895 177.285 99.045 177.455 ;
        RECT 62.895 174.435 63.425 177.285 ;
        RECT 64.155 176.595 80.155 176.765 ;
        RECT 63.925 175.340 64.095 176.380 ;
        RECT 80.215 175.340 80.385 176.380 ;
        RECT 64.155 174.955 80.155 175.125 ;
        RECT 80.885 174.435 81.055 177.285 ;
        RECT 81.785 176.595 97.785 176.765 ;
        RECT 81.555 175.340 81.725 176.380 ;
        RECT 97.845 175.340 98.015 176.380 ;
        RECT 81.785 174.955 97.785 175.125 ;
        RECT 98.515 174.435 99.045 177.285 ;
        RECT 62.895 174.265 99.045 174.435 ;
        RECT 62.895 171.415 63.425 174.265 ;
        RECT 63.925 173.575 80.385 173.745 ;
        RECT 63.925 172.105 64.155 173.575 ;
        RECT 80.155 172.105 80.385 173.575 ;
        RECT 63.925 171.935 80.385 172.105 ;
        RECT 80.885 171.415 81.055 174.265 ;
        RECT 81.555 173.575 98.015 173.745 ;
        RECT 81.555 172.105 81.785 173.575 ;
        RECT 97.785 172.105 98.015 173.575 ;
        RECT 81.555 171.935 98.015 172.105 ;
        RECT 98.515 171.415 99.045 174.265 ;
        RECT 113.860 176.355 151.710 176.885 ;
        RECT 62.895 170.885 99.045 171.415 ;
        RECT 102.740 172.330 110.970 172.500 ;
        RECT 9.330 168.520 52.060 168.690 ;
        RECT 9.330 167.860 51.780 168.030 ;
        RECT 9.330 158.100 9.500 167.860 ;
        RECT 10.290 167.170 12.290 167.340 ;
        RECT 12.580 167.170 14.580 167.340 ;
        RECT 10.060 158.960 10.230 167.000 ;
        RECT 12.350 158.960 12.520 167.000 ;
        RECT 14.640 158.960 14.810 167.000 ;
        RECT 10.290 158.620 12.290 158.790 ;
        RECT 12.580 158.620 14.580 158.790 ;
        RECT 15.370 158.100 15.540 167.860 ;
        RECT 16.330 167.170 18.330 167.340 ;
        RECT 18.620 167.170 20.620 167.340 ;
        RECT 16.100 158.960 16.270 167.000 ;
        RECT 18.390 158.960 18.560 167.000 ;
        RECT 20.680 158.960 20.850 167.000 ;
        RECT 16.330 158.620 18.330 158.790 ;
        RECT 18.620 158.620 20.620 158.790 ;
        RECT 21.410 158.100 21.580 167.860 ;
        RECT 22.370 167.170 24.370 167.340 ;
        RECT 24.660 167.170 26.660 167.340 ;
        RECT 22.140 158.960 22.310 167.000 ;
        RECT 24.430 158.960 24.600 167.000 ;
        RECT 26.720 158.960 26.890 167.000 ;
        RECT 22.370 158.620 24.370 158.790 ;
        RECT 24.660 158.620 26.660 158.790 ;
        RECT 27.450 158.100 27.620 167.860 ;
        RECT 28.410 167.170 30.410 167.340 ;
        RECT 30.700 167.170 32.700 167.340 ;
        RECT 28.180 158.960 28.350 167.000 ;
        RECT 30.470 158.960 30.640 167.000 ;
        RECT 32.760 158.960 32.930 167.000 ;
        RECT 28.410 158.620 30.410 158.790 ;
        RECT 30.700 158.620 32.700 158.790 ;
        RECT 33.490 158.100 33.660 167.860 ;
        RECT 34.450 167.170 36.450 167.340 ;
        RECT 36.740 167.170 38.740 167.340 ;
        RECT 34.220 158.960 34.390 167.000 ;
        RECT 36.510 158.960 36.680 167.000 ;
        RECT 38.800 158.960 38.970 167.000 ;
        RECT 34.450 158.620 36.450 158.790 ;
        RECT 36.740 158.620 38.740 158.790 ;
        RECT 39.530 158.100 39.700 167.860 ;
        RECT 40.490 167.170 42.490 167.340 ;
        RECT 42.780 167.170 44.780 167.340 ;
        RECT 40.260 158.960 40.430 167.000 ;
        RECT 42.550 158.960 42.720 167.000 ;
        RECT 44.840 158.960 45.010 167.000 ;
        RECT 40.490 158.620 42.490 158.790 ;
        RECT 42.780 158.620 44.780 158.790 ;
        RECT 45.570 158.100 45.740 167.860 ;
        RECT 46.530 167.170 48.530 167.340 ;
        RECT 48.820 167.170 50.820 167.340 ;
        RECT 46.300 158.960 46.470 167.000 ;
        RECT 48.590 158.960 48.760 167.000 ;
        RECT 50.880 158.960 51.050 167.000 ;
        RECT 46.530 158.620 48.530 158.790 ;
        RECT 48.820 158.620 50.820 158.790 ;
        RECT 51.610 158.100 51.780 167.860 ;
        RECT 9.330 157.930 51.780 158.100 ;
        RECT 9.330 148.170 9.500 157.930 ;
        RECT 10.290 157.240 12.290 157.410 ;
        RECT 12.580 157.240 14.580 157.410 ;
        RECT 10.060 149.030 10.230 157.070 ;
        RECT 12.350 149.030 12.520 157.070 ;
        RECT 14.640 149.030 14.810 157.070 ;
        RECT 10.290 148.690 12.290 148.860 ;
        RECT 12.580 148.690 14.580 148.860 ;
        RECT 15.370 148.170 15.540 157.930 ;
        RECT 16.330 157.240 18.330 157.410 ;
        RECT 18.620 157.240 20.620 157.410 ;
        RECT 16.100 149.030 16.270 157.070 ;
        RECT 18.390 149.030 18.560 157.070 ;
        RECT 20.680 149.030 20.850 157.070 ;
        RECT 16.330 148.690 18.330 148.860 ;
        RECT 18.620 148.690 20.620 148.860 ;
        RECT 21.410 148.170 21.580 157.930 ;
        RECT 22.370 157.240 24.370 157.410 ;
        RECT 24.660 157.240 26.660 157.410 ;
        RECT 22.140 149.030 22.310 157.070 ;
        RECT 24.430 149.030 24.600 157.070 ;
        RECT 26.720 149.030 26.890 157.070 ;
        RECT 22.370 148.690 24.370 148.860 ;
        RECT 24.660 148.690 26.660 148.860 ;
        RECT 27.450 148.170 27.620 157.930 ;
        RECT 28.410 157.240 30.410 157.410 ;
        RECT 30.700 157.240 32.700 157.410 ;
        RECT 28.180 149.030 28.350 157.070 ;
        RECT 30.470 149.030 30.640 157.070 ;
        RECT 32.760 149.030 32.930 157.070 ;
        RECT 28.410 148.690 30.410 148.860 ;
        RECT 30.700 148.690 32.700 148.860 ;
        RECT 33.490 148.170 33.660 157.930 ;
        RECT 34.450 157.240 36.450 157.410 ;
        RECT 36.740 157.240 38.740 157.410 ;
        RECT 34.220 149.030 34.390 157.070 ;
        RECT 36.510 149.030 36.680 157.070 ;
        RECT 38.800 149.030 38.970 157.070 ;
        RECT 34.450 148.690 36.450 148.860 ;
        RECT 36.740 148.690 38.740 148.860 ;
        RECT 39.530 148.170 39.700 157.930 ;
        RECT 40.490 157.240 42.490 157.410 ;
        RECT 42.780 157.240 44.780 157.410 ;
        RECT 40.260 149.030 40.430 157.070 ;
        RECT 42.550 149.030 42.720 157.070 ;
        RECT 44.840 149.030 45.010 157.070 ;
        RECT 40.490 148.690 42.490 148.860 ;
        RECT 42.780 148.690 44.780 148.860 ;
        RECT 45.570 148.170 45.740 157.930 ;
        RECT 46.530 157.240 48.530 157.410 ;
        RECT 48.820 157.240 50.820 157.410 ;
        RECT 46.300 149.030 46.470 157.070 ;
        RECT 48.590 149.030 48.760 157.070 ;
        RECT 50.880 149.030 51.050 157.070 ;
        RECT 46.530 148.690 48.530 148.860 ;
        RECT 48.820 148.690 50.820 148.860 ;
        RECT 51.610 148.170 51.780 157.930 ;
        RECT 9.330 148.000 51.780 148.170 ;
        RECT 64.100 166.025 96.940 166.425 ;
        RECT 23.195 143.155 58.705 143.745 ;
        RECT 23.195 140.745 23.785 143.155 ;
        RECT 24.515 142.465 32.515 142.635 ;
        RECT 32.805 142.465 40.805 142.635 ;
        RECT 41.095 142.465 49.095 142.635 ;
        RECT 49.385 142.465 57.385 142.635 ;
        RECT 24.285 141.255 24.455 142.295 ;
        RECT 32.575 141.255 32.745 142.295 ;
        RECT 40.865 141.255 41.035 142.295 ;
        RECT 49.155 141.255 49.325 142.295 ;
        RECT 57.445 141.255 57.615 142.295 ;
        RECT 24.515 140.915 32.515 141.085 ;
        RECT 32.805 140.915 40.805 141.085 ;
        RECT 41.095 140.915 49.095 141.085 ;
        RECT 49.385 140.915 57.385 141.085 ;
        RECT 23.195 139.705 24.455 140.745 ;
        RECT 32.575 139.705 32.745 140.745 ;
        RECT 40.865 139.705 41.035 140.745 ;
        RECT 49.155 139.705 49.325 140.745 ;
        RECT 57.445 139.705 57.615 140.745 ;
        RECT 23.195 139.195 23.785 139.705 ;
        RECT 24.515 139.365 32.515 139.535 ;
        RECT 32.805 139.365 40.805 139.535 ;
        RECT 41.095 139.365 49.095 139.535 ;
        RECT 49.385 139.365 57.385 139.535 ;
        RECT 9.430 137.955 20.720 138.485 ;
        RECT 9.430 135.195 9.960 137.955 ;
        RECT 10.995 137.265 11.995 137.435 ;
        RECT 10.765 136.055 10.935 137.095 ;
        RECT 12.055 136.055 12.225 137.095 ;
        RECT 13.030 135.195 13.200 137.955 ;
        RECT 13.930 137.265 14.930 137.435 ;
        RECT 15.220 137.265 16.220 137.435 ;
        RECT 13.700 136.055 13.870 137.095 ;
        RECT 14.990 136.055 15.160 137.095 ;
        RECT 16.280 136.055 16.450 137.095 ;
        RECT 16.950 135.195 17.120 137.955 ;
        RECT 18.155 137.265 19.155 137.435 ;
        RECT 17.925 136.055 18.095 137.095 ;
        RECT 19.215 136.055 19.385 137.095 ;
        RECT 20.190 135.195 20.720 137.955 ;
        RECT 9.430 134.665 20.720 135.195 ;
        RECT 23.195 138.155 24.455 139.195 ;
        RECT 32.575 138.155 32.745 139.195 ;
        RECT 40.865 138.155 41.035 139.195 ;
        RECT 49.155 138.155 49.325 139.195 ;
        RECT 57.445 138.155 57.615 139.195 ;
        RECT 23.195 135.745 23.785 138.155 ;
        RECT 24.515 137.815 32.515 137.985 ;
        RECT 32.805 137.815 40.805 137.985 ;
        RECT 41.095 137.815 49.095 137.985 ;
        RECT 49.385 137.815 57.385 137.985 ;
        RECT 24.285 136.605 24.455 137.645 ;
        RECT 32.575 136.605 32.745 137.645 ;
        RECT 40.865 136.605 41.035 137.645 ;
        RECT 49.155 136.605 49.325 137.645 ;
        RECT 57.445 136.605 57.615 137.645 ;
        RECT 24.515 136.265 32.515 136.435 ;
        RECT 32.805 136.265 40.805 136.435 ;
        RECT 41.095 136.265 49.095 136.435 ;
        RECT 49.385 136.265 57.385 136.435 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 23.195 135.155 58.705 135.745 ;
        RECT 64.100 133.985 64.500 166.025 ;
        RECT 69.635 160.720 91.405 160.890 ;
        RECT 69.635 139.290 69.805 160.720 ;
        RECT 71.220 158.800 89.820 159.305 ;
        RECT 71.220 156.090 71.725 158.800 ;
        RECT 72.035 158.130 74.125 158.490 ;
        RECT 72.035 156.760 72.395 158.130 ;
        RECT 72.685 157.050 73.475 157.840 ;
        RECT 73.765 156.760 74.125 158.130 ;
        RECT 72.035 156.400 74.125 156.760 ;
        RECT 74.435 156.090 75.445 158.800 ;
        RECT 75.755 158.130 77.845 158.490 ;
        RECT 75.755 156.760 76.115 158.130 ;
        RECT 76.405 157.050 77.195 157.840 ;
        RECT 77.485 156.760 77.845 158.130 ;
        RECT 75.755 156.400 77.845 156.760 ;
        RECT 78.155 156.090 79.165 158.800 ;
        RECT 79.475 158.130 81.565 158.490 ;
        RECT 79.475 156.760 79.835 158.130 ;
        RECT 80.125 157.050 80.915 157.840 ;
        RECT 81.205 156.760 81.565 158.130 ;
        RECT 79.475 156.400 81.565 156.760 ;
        RECT 81.875 156.090 82.885 158.800 ;
        RECT 83.195 158.130 85.285 158.490 ;
        RECT 83.195 156.760 83.555 158.130 ;
        RECT 83.845 157.050 84.635 157.840 ;
        RECT 84.925 156.760 85.285 158.130 ;
        RECT 83.195 156.400 85.285 156.760 ;
        RECT 85.595 156.090 86.605 158.800 ;
        RECT 86.915 158.130 89.005 158.490 ;
        RECT 86.915 156.760 87.275 158.130 ;
        RECT 87.565 157.050 88.355 157.840 ;
        RECT 88.645 156.760 89.005 158.130 ;
        RECT 86.915 156.400 89.005 156.760 ;
        RECT 89.315 156.090 89.820 158.800 ;
        RECT 71.220 155.080 89.820 156.090 ;
        RECT 71.220 152.370 71.725 155.080 ;
        RECT 72.035 154.410 74.125 154.770 ;
        RECT 72.035 153.040 72.395 154.410 ;
        RECT 72.685 153.330 73.475 154.120 ;
        RECT 73.765 153.040 74.125 154.410 ;
        RECT 72.035 152.680 74.125 153.040 ;
        RECT 74.435 152.370 75.445 155.080 ;
        RECT 75.755 154.410 77.845 154.770 ;
        RECT 75.755 153.040 76.115 154.410 ;
        RECT 76.405 153.330 77.195 154.120 ;
        RECT 77.485 153.040 77.845 154.410 ;
        RECT 75.755 152.680 77.845 153.040 ;
        RECT 78.155 152.370 79.165 155.080 ;
        RECT 79.475 154.410 81.565 154.770 ;
        RECT 79.475 153.040 79.835 154.410 ;
        RECT 80.125 153.330 80.915 154.120 ;
        RECT 81.205 153.040 81.565 154.410 ;
        RECT 79.475 152.680 81.565 153.040 ;
        RECT 81.875 152.370 82.885 155.080 ;
        RECT 83.195 154.410 85.285 154.770 ;
        RECT 83.195 153.040 83.555 154.410 ;
        RECT 83.845 153.330 84.635 154.120 ;
        RECT 84.925 153.040 85.285 154.410 ;
        RECT 83.195 152.680 85.285 153.040 ;
        RECT 85.595 152.370 86.605 155.080 ;
        RECT 86.915 154.410 89.005 154.770 ;
        RECT 86.915 153.040 87.275 154.410 ;
        RECT 87.565 153.330 88.355 154.120 ;
        RECT 88.645 153.040 89.005 154.410 ;
        RECT 86.915 152.680 89.005 153.040 ;
        RECT 89.315 152.370 89.820 155.080 ;
        RECT 71.220 151.360 89.820 152.370 ;
        RECT 71.220 148.650 71.725 151.360 ;
        RECT 72.035 150.690 74.125 151.050 ;
        RECT 72.035 149.320 72.395 150.690 ;
        RECT 72.685 149.610 73.475 150.400 ;
        RECT 73.765 149.320 74.125 150.690 ;
        RECT 72.035 148.960 74.125 149.320 ;
        RECT 74.435 148.650 75.445 151.360 ;
        RECT 75.755 150.690 77.845 151.050 ;
        RECT 75.755 149.320 76.115 150.690 ;
        RECT 76.405 149.610 77.195 150.400 ;
        RECT 77.485 149.320 77.845 150.690 ;
        RECT 75.755 148.960 77.845 149.320 ;
        RECT 78.155 148.650 79.165 151.360 ;
        RECT 79.475 150.690 81.565 151.050 ;
        RECT 79.475 149.320 79.835 150.690 ;
        RECT 80.125 149.610 80.915 150.400 ;
        RECT 81.205 149.320 81.565 150.690 ;
        RECT 79.475 148.960 81.565 149.320 ;
        RECT 81.875 148.650 82.885 151.360 ;
        RECT 83.195 150.690 85.285 151.050 ;
        RECT 83.195 149.320 83.555 150.690 ;
        RECT 83.845 149.610 84.635 150.400 ;
        RECT 84.925 149.320 85.285 150.690 ;
        RECT 83.195 148.960 85.285 149.320 ;
        RECT 85.595 148.650 86.605 151.360 ;
        RECT 86.915 150.690 89.005 151.050 ;
        RECT 86.915 149.320 87.275 150.690 ;
        RECT 87.565 149.610 88.355 150.400 ;
        RECT 88.645 149.320 89.005 150.690 ;
        RECT 86.915 148.960 89.005 149.320 ;
        RECT 89.315 148.650 89.820 151.360 ;
        RECT 71.220 147.640 89.820 148.650 ;
        RECT 71.220 144.930 71.725 147.640 ;
        RECT 72.035 146.970 74.125 147.330 ;
        RECT 72.035 145.600 72.395 146.970 ;
        RECT 72.685 145.890 73.475 146.680 ;
        RECT 73.765 145.600 74.125 146.970 ;
        RECT 72.035 145.240 74.125 145.600 ;
        RECT 74.435 144.930 75.445 147.640 ;
        RECT 75.755 146.970 77.845 147.330 ;
        RECT 75.755 145.600 76.115 146.970 ;
        RECT 76.405 145.890 77.195 146.680 ;
        RECT 77.485 145.600 77.845 146.970 ;
        RECT 75.755 145.240 77.845 145.600 ;
        RECT 78.155 144.930 79.165 147.640 ;
        RECT 79.475 146.970 81.565 147.330 ;
        RECT 79.475 145.600 79.835 146.970 ;
        RECT 80.125 145.890 80.915 146.680 ;
        RECT 81.205 145.600 81.565 146.970 ;
        RECT 79.475 145.240 81.565 145.600 ;
        RECT 81.875 144.930 82.885 147.640 ;
        RECT 83.195 146.970 85.285 147.330 ;
        RECT 83.195 145.600 83.555 146.970 ;
        RECT 83.845 145.890 84.635 146.680 ;
        RECT 84.925 145.600 85.285 146.970 ;
        RECT 83.195 145.240 85.285 145.600 ;
        RECT 85.595 144.930 86.605 147.640 ;
        RECT 86.915 146.970 89.005 147.330 ;
        RECT 86.915 145.600 87.275 146.970 ;
        RECT 87.565 145.890 88.355 146.680 ;
        RECT 88.645 145.600 89.005 146.970 ;
        RECT 86.915 145.240 89.005 145.600 ;
        RECT 89.315 144.930 89.820 147.640 ;
        RECT 71.220 143.920 89.820 144.930 ;
        RECT 71.220 141.210 71.725 143.920 ;
        RECT 72.035 143.250 74.125 143.610 ;
        RECT 72.035 141.880 72.395 143.250 ;
        RECT 72.685 142.170 73.475 142.960 ;
        RECT 73.765 141.880 74.125 143.250 ;
        RECT 72.035 141.520 74.125 141.880 ;
        RECT 74.435 141.210 75.445 143.920 ;
        RECT 75.755 143.250 77.845 143.610 ;
        RECT 75.755 141.880 76.115 143.250 ;
        RECT 76.405 142.170 77.195 142.960 ;
        RECT 77.485 141.880 77.845 143.250 ;
        RECT 75.755 141.520 77.845 141.880 ;
        RECT 78.155 141.210 79.165 143.920 ;
        RECT 79.475 143.250 81.565 143.610 ;
        RECT 79.475 141.880 79.835 143.250 ;
        RECT 80.125 142.170 80.915 142.960 ;
        RECT 81.205 141.880 81.565 143.250 ;
        RECT 79.475 141.520 81.565 141.880 ;
        RECT 81.875 141.210 82.885 143.920 ;
        RECT 83.195 143.250 85.285 143.610 ;
        RECT 83.195 141.880 83.555 143.250 ;
        RECT 83.845 142.170 84.635 142.960 ;
        RECT 84.925 141.880 85.285 143.250 ;
        RECT 83.195 141.520 85.285 141.880 ;
        RECT 85.595 141.210 86.605 143.920 ;
        RECT 86.915 143.250 89.005 143.610 ;
        RECT 86.915 141.880 87.275 143.250 ;
        RECT 87.565 142.170 88.355 142.960 ;
        RECT 88.645 141.880 89.005 143.250 ;
        RECT 86.915 141.520 89.005 141.880 ;
        RECT 89.315 141.210 89.820 143.920 ;
        RECT 71.220 140.705 89.820 141.210 ;
        RECT 91.235 139.290 91.405 160.720 ;
        RECT 69.635 139.120 91.405 139.290 ;
        RECT 96.540 133.985 96.940 166.025 ;
        RECT 102.740 162.570 102.910 172.330 ;
        RECT 103.695 171.640 104.695 171.810 ;
        RECT 104.985 171.640 105.985 171.810 ;
        RECT 103.465 163.430 103.635 171.470 ;
        RECT 104.755 163.430 104.925 171.470 ;
        RECT 106.045 163.430 106.215 171.470 ;
        RECT 103.695 163.090 104.695 163.260 ;
        RECT 104.985 163.090 105.985 163.260 ;
        RECT 106.770 162.570 106.940 172.330 ;
        RECT 107.725 171.640 108.725 171.810 ;
        RECT 109.015 171.640 110.015 171.810 ;
        RECT 107.495 163.430 107.665 171.470 ;
        RECT 108.785 163.430 108.955 171.470 ;
        RECT 110.075 163.430 110.245 171.470 ;
        RECT 107.725 163.090 108.725 163.260 ;
        RECT 109.015 163.090 110.015 163.260 ;
        RECT 110.800 162.570 110.970 172.330 ;
        RECT 113.860 166.595 114.390 176.355 ;
        RECT 115.180 175.665 115.680 175.835 ;
        RECT 115.970 175.665 116.470 175.835 ;
        RECT 116.760 175.665 117.260 175.835 ;
        RECT 117.550 175.665 118.050 175.835 ;
        RECT 114.950 167.455 115.120 175.495 ;
        RECT 115.740 167.455 115.910 175.495 ;
        RECT 116.530 167.455 116.700 175.495 ;
        RECT 117.320 167.455 117.490 175.495 ;
        RECT 118.110 167.455 118.280 175.495 ;
        RECT 115.180 167.115 115.680 167.285 ;
        RECT 115.970 167.115 116.470 167.285 ;
        RECT 116.760 167.115 117.260 167.285 ;
        RECT 117.550 167.115 118.050 167.285 ;
        RECT 118.840 166.595 119.010 176.355 ;
        RECT 119.800 175.665 120.300 175.835 ;
        RECT 120.590 175.665 121.090 175.835 ;
        RECT 121.380 175.665 121.880 175.835 ;
        RECT 122.170 175.665 122.670 175.835 ;
        RECT 119.570 167.455 119.740 175.495 ;
        RECT 120.360 167.455 120.530 175.495 ;
        RECT 121.150 167.455 121.320 175.495 ;
        RECT 121.940 167.455 122.110 175.495 ;
        RECT 122.730 167.455 122.900 175.495 ;
        RECT 119.800 167.115 120.300 167.285 ;
        RECT 120.590 167.115 121.090 167.285 ;
        RECT 121.380 167.115 121.880 167.285 ;
        RECT 122.170 167.115 122.670 167.285 ;
        RECT 123.460 166.595 123.630 176.355 ;
        RECT 124.420 175.665 124.920 175.835 ;
        RECT 125.210 175.665 125.710 175.835 ;
        RECT 126.000 175.665 126.500 175.835 ;
        RECT 126.790 175.665 127.290 175.835 ;
        RECT 124.190 167.455 124.360 175.495 ;
        RECT 124.980 167.455 125.150 175.495 ;
        RECT 125.770 167.455 125.940 175.495 ;
        RECT 126.560 167.455 126.730 175.495 ;
        RECT 127.350 167.455 127.520 175.495 ;
        RECT 124.420 167.115 124.920 167.285 ;
        RECT 125.210 167.115 125.710 167.285 ;
        RECT 126.000 167.115 126.500 167.285 ;
        RECT 126.790 167.115 127.290 167.285 ;
        RECT 128.080 166.595 128.250 176.355 ;
        RECT 129.040 175.665 129.540 175.835 ;
        RECT 129.830 175.665 130.330 175.835 ;
        RECT 130.620 175.665 131.120 175.835 ;
        RECT 131.410 175.665 131.910 175.835 ;
        RECT 128.810 167.455 128.980 175.495 ;
        RECT 129.600 167.455 129.770 175.495 ;
        RECT 130.390 167.455 130.560 175.495 ;
        RECT 131.180 167.455 131.350 175.495 ;
        RECT 131.970 167.455 132.140 175.495 ;
        RECT 129.040 167.115 129.540 167.285 ;
        RECT 129.830 167.115 130.330 167.285 ;
        RECT 130.620 167.115 131.120 167.285 ;
        RECT 131.410 167.115 131.910 167.285 ;
        RECT 132.700 166.595 132.870 176.355 ;
        RECT 133.660 175.665 134.160 175.835 ;
        RECT 134.450 175.665 134.950 175.835 ;
        RECT 135.240 175.665 135.740 175.835 ;
        RECT 136.030 175.665 136.530 175.835 ;
        RECT 133.430 167.455 133.600 175.495 ;
        RECT 134.220 167.455 134.390 175.495 ;
        RECT 135.010 167.455 135.180 175.495 ;
        RECT 135.800 167.455 135.970 175.495 ;
        RECT 136.590 167.455 136.760 175.495 ;
        RECT 133.660 167.115 134.160 167.285 ;
        RECT 134.450 167.115 134.950 167.285 ;
        RECT 135.240 167.115 135.740 167.285 ;
        RECT 136.030 167.115 136.530 167.285 ;
        RECT 137.320 166.595 137.490 176.355 ;
        RECT 138.280 175.665 138.780 175.835 ;
        RECT 139.070 175.665 139.570 175.835 ;
        RECT 139.860 175.665 140.360 175.835 ;
        RECT 140.650 175.665 141.150 175.835 ;
        RECT 138.050 167.455 138.220 175.495 ;
        RECT 138.840 167.455 139.010 175.495 ;
        RECT 139.630 167.455 139.800 175.495 ;
        RECT 140.420 167.455 140.590 175.495 ;
        RECT 141.210 167.455 141.380 175.495 ;
        RECT 138.280 167.115 138.780 167.285 ;
        RECT 139.070 167.115 139.570 167.285 ;
        RECT 139.860 167.115 140.360 167.285 ;
        RECT 140.650 167.115 141.150 167.285 ;
        RECT 141.940 166.595 142.110 176.355 ;
        RECT 142.900 175.665 143.400 175.835 ;
        RECT 143.690 175.665 144.190 175.835 ;
        RECT 144.480 175.665 144.980 175.835 ;
        RECT 145.270 175.665 145.770 175.835 ;
        RECT 142.670 167.455 142.840 175.495 ;
        RECT 143.460 167.455 143.630 175.495 ;
        RECT 144.250 167.455 144.420 175.495 ;
        RECT 145.040 167.455 145.210 175.495 ;
        RECT 145.830 167.455 146.000 175.495 ;
        RECT 142.900 167.115 143.400 167.285 ;
        RECT 143.690 167.115 144.190 167.285 ;
        RECT 144.480 167.115 144.980 167.285 ;
        RECT 145.270 167.115 145.770 167.285 ;
        RECT 146.560 166.595 146.730 176.355 ;
        RECT 147.520 175.665 148.020 175.835 ;
        RECT 148.310 175.665 148.810 175.835 ;
        RECT 149.100 175.665 149.600 175.835 ;
        RECT 149.890 175.665 150.390 175.835 ;
        RECT 147.290 167.455 147.460 175.495 ;
        RECT 148.080 167.455 148.250 175.495 ;
        RECT 148.870 167.455 149.040 175.495 ;
        RECT 149.660 167.455 149.830 175.495 ;
        RECT 150.450 167.455 150.620 175.495 ;
        RECT 147.520 167.115 148.020 167.285 ;
        RECT 148.310 167.115 148.810 167.285 ;
        RECT 149.100 167.115 149.600 167.285 ;
        RECT 149.890 167.115 150.390 167.285 ;
        RECT 151.180 166.595 151.710 176.355 ;
        RECT 113.860 166.065 151.710 166.595 ;
        RECT 102.740 162.400 110.970 162.570 ;
        RECT 102.740 158.640 102.910 162.400 ;
        RECT 103.465 159.500 103.635 161.540 ;
        RECT 104.755 159.500 104.925 161.540 ;
        RECT 106.045 159.500 106.215 161.540 ;
        RECT 103.695 159.160 104.695 159.330 ;
        RECT 104.985 159.160 105.985 159.330 ;
        RECT 106.770 158.640 106.940 162.400 ;
        RECT 107.495 159.500 107.665 161.540 ;
        RECT 108.785 159.500 108.955 161.540 ;
        RECT 110.075 159.500 110.245 161.540 ;
        RECT 107.725 159.160 108.725 159.330 ;
        RECT 109.015 159.160 110.015 159.330 ;
        RECT 110.800 158.640 110.970 162.400 ;
        RECT 102.740 158.470 110.970 158.640 ;
        RECT 116.015 157.500 149.445 158.030 ;
        RECT 102.740 155.775 110.970 155.945 ;
        RECT 102.740 151.925 102.910 155.775 ;
        RECT 103.695 155.085 104.695 155.255 ;
        RECT 104.985 155.085 105.985 155.255 ;
        RECT 103.465 152.830 103.635 154.870 ;
        RECT 104.755 152.830 104.925 154.870 ;
        RECT 106.045 152.830 106.215 154.870 ;
        RECT 106.770 151.925 106.940 155.775 ;
        RECT 107.725 155.085 108.725 155.255 ;
        RECT 109.015 155.085 110.015 155.255 ;
        RECT 107.495 152.830 107.665 154.870 ;
        RECT 108.785 152.830 108.955 154.870 ;
        RECT 110.075 152.830 110.245 154.870 ;
        RECT 110.800 151.925 110.970 155.775 ;
        RECT 102.740 151.755 110.970 151.925 ;
        RECT 102.740 141.905 102.910 151.755 ;
        RECT 103.695 151.065 104.695 151.235 ;
        RECT 104.985 151.065 105.985 151.235 ;
        RECT 103.465 142.810 103.635 150.850 ;
        RECT 104.755 142.810 104.925 150.850 ;
        RECT 106.045 142.810 106.215 150.850 ;
        RECT 103.695 142.425 104.695 142.595 ;
        RECT 104.985 142.425 105.985 142.595 ;
        RECT 106.770 141.905 106.940 151.755 ;
        RECT 107.725 151.065 108.725 151.235 ;
        RECT 109.015 151.065 110.015 151.235 ;
        RECT 107.495 142.810 107.665 150.850 ;
        RECT 108.785 142.810 108.955 150.850 ;
        RECT 110.075 142.810 110.245 150.850 ;
        RECT 107.725 142.425 108.725 142.595 ;
        RECT 109.015 142.425 110.015 142.595 ;
        RECT 110.800 141.905 110.970 151.755 ;
        RECT 102.740 141.735 110.970 141.905 ;
        RECT 116.015 140.250 116.545 157.500 ;
        RECT 117.130 156.135 119.290 156.825 ;
        RECT 117.130 154.965 119.290 155.655 ;
        RECT 117.130 153.795 119.290 154.485 ;
        RECT 117.130 152.625 119.290 153.315 ;
        RECT 117.130 151.455 119.290 152.145 ;
        RECT 117.130 150.285 119.290 150.975 ;
        RECT 117.130 149.115 119.290 149.805 ;
        RECT 117.130 147.945 119.290 148.635 ;
        RECT 117.130 146.775 119.290 147.465 ;
        RECT 117.130 145.605 119.290 146.295 ;
        RECT 117.130 144.435 119.290 145.125 ;
        RECT 117.130 143.265 119.290 143.955 ;
        RECT 117.130 142.095 119.290 142.785 ;
        RECT 117.130 140.925 119.290 141.615 ;
        RECT 119.595 140.250 122.075 157.500 ;
        RECT 122.380 156.135 124.540 156.825 ;
        RECT 125.060 156.135 127.220 156.825 ;
        RECT 122.380 154.965 124.540 155.655 ;
        RECT 125.060 154.965 127.220 155.655 ;
        RECT 122.380 153.795 124.540 154.485 ;
        RECT 125.060 153.795 127.220 154.485 ;
        RECT 122.380 152.625 124.540 153.315 ;
        RECT 125.060 152.625 127.220 153.315 ;
        RECT 122.380 151.455 124.540 152.145 ;
        RECT 125.060 151.455 127.220 152.145 ;
        RECT 122.380 150.285 124.540 150.975 ;
        RECT 125.060 150.285 127.220 150.975 ;
        RECT 122.380 149.115 124.540 149.805 ;
        RECT 125.060 149.115 127.220 149.805 ;
        RECT 122.380 147.945 124.540 148.635 ;
        RECT 125.060 147.945 127.220 148.635 ;
        RECT 122.380 146.775 124.540 147.465 ;
        RECT 125.060 146.775 127.220 147.465 ;
        RECT 122.380 145.605 124.540 146.295 ;
        RECT 125.060 145.605 127.220 146.295 ;
        RECT 122.380 144.435 124.540 145.125 ;
        RECT 125.060 144.435 127.220 145.125 ;
        RECT 122.380 143.265 124.540 143.955 ;
        RECT 125.060 143.265 127.220 143.955 ;
        RECT 122.380 142.095 124.540 142.785 ;
        RECT 125.060 142.095 127.220 142.785 ;
        RECT 122.380 140.925 124.540 141.615 ;
        RECT 125.060 140.925 127.220 141.615 ;
        RECT 127.525 140.250 130.005 157.500 ;
        RECT 130.310 156.135 132.470 156.825 ;
        RECT 132.990 156.135 135.150 156.825 ;
        RECT 130.310 154.965 132.470 155.655 ;
        RECT 132.990 154.965 135.150 155.655 ;
        RECT 130.310 153.795 132.470 154.485 ;
        RECT 132.990 153.795 135.150 154.485 ;
        RECT 130.310 152.625 132.470 153.315 ;
        RECT 132.990 152.625 135.150 153.315 ;
        RECT 130.310 151.455 132.470 152.145 ;
        RECT 132.990 151.455 135.150 152.145 ;
        RECT 130.310 150.285 132.470 150.975 ;
        RECT 132.990 150.285 135.150 150.975 ;
        RECT 130.310 149.115 132.470 149.805 ;
        RECT 132.990 149.115 135.150 149.805 ;
        RECT 130.310 147.945 132.470 148.635 ;
        RECT 132.990 147.945 135.150 148.635 ;
        RECT 130.310 146.775 132.470 147.465 ;
        RECT 132.990 146.775 135.150 147.465 ;
        RECT 130.310 145.605 132.470 146.295 ;
        RECT 132.990 145.605 135.150 146.295 ;
        RECT 130.310 144.435 132.470 145.125 ;
        RECT 132.990 144.435 135.150 145.125 ;
        RECT 130.310 143.265 132.470 143.955 ;
        RECT 132.990 143.265 135.150 143.955 ;
        RECT 130.310 142.095 132.470 142.785 ;
        RECT 132.990 142.095 135.150 142.785 ;
        RECT 130.310 140.925 132.470 141.615 ;
        RECT 132.990 140.925 135.150 141.615 ;
        RECT 135.455 140.250 137.935 157.500 ;
        RECT 138.240 156.135 140.400 156.825 ;
        RECT 140.920 156.135 143.080 156.825 ;
        RECT 138.240 154.965 140.400 155.655 ;
        RECT 140.920 154.965 143.080 155.655 ;
        RECT 138.240 153.795 140.400 154.485 ;
        RECT 140.920 153.795 143.080 154.485 ;
        RECT 138.240 152.625 140.400 153.315 ;
        RECT 140.920 152.625 143.080 153.315 ;
        RECT 138.240 151.455 140.400 152.145 ;
        RECT 140.920 151.455 143.080 152.145 ;
        RECT 138.240 150.285 140.400 150.975 ;
        RECT 140.920 150.285 143.080 150.975 ;
        RECT 138.240 149.115 140.400 149.805 ;
        RECT 140.920 149.115 143.080 149.805 ;
        RECT 138.240 147.945 140.400 148.635 ;
        RECT 140.920 147.945 143.080 148.635 ;
        RECT 138.240 146.775 140.400 147.465 ;
        RECT 140.920 146.775 143.080 147.465 ;
        RECT 138.240 145.605 140.400 146.295 ;
        RECT 140.920 145.605 143.080 146.295 ;
        RECT 138.240 144.435 140.400 145.125 ;
        RECT 140.920 144.435 143.080 145.125 ;
        RECT 138.240 143.265 140.400 143.955 ;
        RECT 140.920 143.265 143.080 143.955 ;
        RECT 138.240 142.095 140.400 142.785 ;
        RECT 140.920 142.095 143.080 142.785 ;
        RECT 138.240 140.925 140.400 141.615 ;
        RECT 140.920 140.925 143.080 141.615 ;
        RECT 143.385 140.250 145.865 157.500 ;
        RECT 146.170 156.135 148.330 156.825 ;
        RECT 146.170 154.965 148.330 155.655 ;
        RECT 146.170 153.795 148.330 154.485 ;
        RECT 146.170 152.625 148.330 153.315 ;
        RECT 146.170 151.455 148.330 152.145 ;
        RECT 146.170 150.285 148.330 150.975 ;
        RECT 146.170 149.115 148.330 149.805 ;
        RECT 146.170 147.945 148.330 148.635 ;
        RECT 146.170 146.775 148.330 147.465 ;
        RECT 146.170 145.605 148.330 146.295 ;
        RECT 146.170 144.435 148.330 145.125 ;
        RECT 146.170 143.265 148.330 143.955 ;
        RECT 146.170 142.095 148.330 142.785 ;
        RECT 146.170 140.925 148.330 141.615 ;
        RECT 148.915 140.250 149.445 157.500 ;
        RECT 116.015 139.720 149.445 140.250 ;
        RECT 64.100 133.585 96.940 133.985 ;
        RECT 138.110 134.130 145.930 134.660 ;
        RECT 138.110 130.280 138.640 134.130 ;
        RECT 139.465 133.440 140.465 133.610 ;
        RECT 140.755 133.440 141.755 133.610 ;
        RECT 139.235 131.185 139.405 133.225 ;
        RECT 140.525 131.185 140.695 133.225 ;
        RECT 141.815 131.185 141.985 133.225 ;
        RECT 142.580 130.280 142.750 134.130 ;
        RECT 143.345 131.185 143.515 133.225 ;
        RECT 144.635 131.185 144.805 133.225 ;
        RECT 143.575 130.800 144.575 130.970 ;
        RECT 145.400 130.280 145.930 134.130 ;
        RECT 138.110 129.750 145.930 130.280 ;
        RECT 138.110 128.410 145.930 128.940 ;
        RECT 138.110 124.650 138.640 128.410 ;
        RECT 139.235 125.510 139.405 127.550 ;
        RECT 140.525 125.510 140.695 127.550 ;
        RECT 141.815 125.510 141.985 127.550 ;
        RECT 139.465 125.170 140.465 125.340 ;
        RECT 140.755 125.170 141.755 125.340 ;
        RECT 142.580 124.650 142.750 128.410 ;
        RECT 143.575 127.720 144.575 127.890 ;
        RECT 143.345 125.510 143.515 127.550 ;
        RECT 144.635 125.510 144.805 127.550 ;
        RECT 145.400 124.650 145.930 128.410 ;
        RECT 10.055 123.725 70.145 124.255 ;
        RECT 10.055 113.875 10.585 123.725 ;
        RECT 11.315 123.035 13.315 123.205 ;
        RECT 13.605 123.035 15.605 123.205 ;
        RECT 11.085 114.780 11.255 122.820 ;
        RECT 13.375 114.780 13.545 122.820 ;
        RECT 15.665 114.780 15.835 122.820 ;
        RECT 11.315 114.395 13.315 114.565 ;
        RECT 13.605 114.395 15.605 114.565 ;
        RECT 16.335 113.875 16.505 123.725 ;
        RECT 17.235 123.035 19.235 123.205 ;
        RECT 19.525 123.035 21.525 123.205 ;
        RECT 17.005 114.780 17.175 122.820 ;
        RECT 19.295 114.780 19.465 122.820 ;
        RECT 21.585 114.780 21.755 122.820 ;
        RECT 17.235 114.395 19.235 114.565 ;
        RECT 19.525 114.395 21.525 114.565 ;
        RECT 22.255 113.875 22.425 123.725 ;
        RECT 23.155 123.035 25.155 123.205 ;
        RECT 25.445 123.035 27.445 123.205 ;
        RECT 22.925 114.780 23.095 122.820 ;
        RECT 25.215 114.780 25.385 122.820 ;
        RECT 27.505 114.780 27.675 122.820 ;
        RECT 23.155 114.395 25.155 114.565 ;
        RECT 25.445 114.395 27.445 114.565 ;
        RECT 28.175 113.875 28.345 123.725 ;
        RECT 29.075 123.035 31.075 123.205 ;
        RECT 31.365 123.035 33.365 123.205 ;
        RECT 28.845 114.780 29.015 122.820 ;
        RECT 31.135 114.780 31.305 122.820 ;
        RECT 33.425 114.780 33.595 122.820 ;
        RECT 29.075 114.395 31.075 114.565 ;
        RECT 31.365 114.395 33.365 114.565 ;
        RECT 34.095 113.875 34.265 123.725 ;
        RECT 34.995 123.035 36.995 123.205 ;
        RECT 37.285 123.035 39.285 123.205 ;
        RECT 34.765 114.780 34.935 122.820 ;
        RECT 37.055 114.780 37.225 122.820 ;
        RECT 39.345 114.780 39.515 122.820 ;
        RECT 34.995 114.395 36.995 114.565 ;
        RECT 37.285 114.395 39.285 114.565 ;
        RECT 40.015 113.875 40.185 123.725 ;
        RECT 40.915 123.035 42.915 123.205 ;
        RECT 43.205 123.035 45.205 123.205 ;
        RECT 40.685 114.780 40.855 122.820 ;
        RECT 42.975 114.780 43.145 122.820 ;
        RECT 45.265 114.780 45.435 122.820 ;
        RECT 40.915 114.395 42.915 114.565 ;
        RECT 43.205 114.395 45.205 114.565 ;
        RECT 45.935 113.875 46.105 123.725 ;
        RECT 46.835 123.035 48.835 123.205 ;
        RECT 49.125 123.035 51.125 123.205 ;
        RECT 46.605 114.780 46.775 122.820 ;
        RECT 48.895 114.780 49.065 122.820 ;
        RECT 51.185 114.780 51.355 122.820 ;
        RECT 46.835 114.395 48.835 114.565 ;
        RECT 49.125 114.395 51.125 114.565 ;
        RECT 51.855 113.875 52.025 123.725 ;
        RECT 52.755 123.035 54.755 123.205 ;
        RECT 55.045 123.035 57.045 123.205 ;
        RECT 52.525 114.780 52.695 122.820 ;
        RECT 54.815 114.780 54.985 122.820 ;
        RECT 57.105 114.780 57.275 122.820 ;
        RECT 52.755 114.395 54.755 114.565 ;
        RECT 55.045 114.395 57.045 114.565 ;
        RECT 57.775 113.875 57.945 123.725 ;
        RECT 58.675 123.035 60.675 123.205 ;
        RECT 60.965 123.035 62.965 123.205 ;
        RECT 58.445 114.780 58.615 122.820 ;
        RECT 60.735 114.780 60.905 122.820 ;
        RECT 63.025 114.780 63.195 122.820 ;
        RECT 58.675 114.395 60.675 114.565 ;
        RECT 60.965 114.395 62.965 114.565 ;
        RECT 63.695 113.875 63.865 123.725 ;
        RECT 64.595 123.035 66.595 123.205 ;
        RECT 66.885 123.035 68.885 123.205 ;
        RECT 64.365 114.780 64.535 122.820 ;
        RECT 66.655 114.780 66.825 122.820 ;
        RECT 68.945 114.780 69.115 122.820 ;
        RECT 64.595 114.395 66.595 114.565 ;
        RECT 66.885 114.395 68.885 114.565 ;
        RECT 69.615 113.875 70.145 123.725 ;
        RECT 10.055 113.705 70.145 113.875 ;
        RECT 10.055 103.855 10.585 113.705 ;
        RECT 11.315 113.015 13.315 113.185 ;
        RECT 13.605 113.015 15.605 113.185 ;
        RECT 11.085 104.760 11.255 112.800 ;
        RECT 13.375 104.760 13.545 112.800 ;
        RECT 15.665 104.760 15.835 112.800 ;
        RECT 11.315 104.375 13.315 104.545 ;
        RECT 13.605 104.375 15.605 104.545 ;
        RECT 16.335 103.855 16.505 113.705 ;
        RECT 17.235 113.015 19.235 113.185 ;
        RECT 19.525 113.015 21.525 113.185 ;
        RECT 17.005 104.760 17.175 112.800 ;
        RECT 19.295 104.760 19.465 112.800 ;
        RECT 21.585 104.760 21.755 112.800 ;
        RECT 17.235 104.375 19.235 104.545 ;
        RECT 19.525 104.375 21.525 104.545 ;
        RECT 22.255 103.855 22.425 113.705 ;
        RECT 23.155 113.015 25.155 113.185 ;
        RECT 25.445 113.015 27.445 113.185 ;
        RECT 22.925 104.760 23.095 112.800 ;
        RECT 25.215 104.760 25.385 112.800 ;
        RECT 27.505 104.760 27.675 112.800 ;
        RECT 23.155 104.375 25.155 104.545 ;
        RECT 25.445 104.375 27.445 104.545 ;
        RECT 28.175 103.855 28.345 113.705 ;
        RECT 29.075 113.015 31.075 113.185 ;
        RECT 31.365 113.015 33.365 113.185 ;
        RECT 28.845 104.760 29.015 112.800 ;
        RECT 31.135 104.760 31.305 112.800 ;
        RECT 33.425 104.760 33.595 112.800 ;
        RECT 29.075 104.375 31.075 104.545 ;
        RECT 31.365 104.375 33.365 104.545 ;
        RECT 34.095 103.855 34.265 113.705 ;
        RECT 34.995 113.015 36.995 113.185 ;
        RECT 37.285 113.015 39.285 113.185 ;
        RECT 34.765 104.760 34.935 112.800 ;
        RECT 37.055 104.760 37.225 112.800 ;
        RECT 39.345 104.760 39.515 112.800 ;
        RECT 34.995 104.375 36.995 104.545 ;
        RECT 37.285 104.375 39.285 104.545 ;
        RECT 40.015 103.855 40.185 113.705 ;
        RECT 40.915 113.015 42.915 113.185 ;
        RECT 43.205 113.015 45.205 113.185 ;
        RECT 40.685 104.760 40.855 112.800 ;
        RECT 42.975 104.760 43.145 112.800 ;
        RECT 45.265 104.760 45.435 112.800 ;
        RECT 40.915 104.375 42.915 104.545 ;
        RECT 43.205 104.375 45.205 104.545 ;
        RECT 45.935 103.855 46.105 113.705 ;
        RECT 46.835 113.015 48.835 113.185 ;
        RECT 49.125 113.015 51.125 113.185 ;
        RECT 46.605 104.760 46.775 112.800 ;
        RECT 48.895 104.760 49.065 112.800 ;
        RECT 51.185 104.760 51.355 112.800 ;
        RECT 46.835 104.375 48.835 104.545 ;
        RECT 49.125 104.375 51.125 104.545 ;
        RECT 51.855 103.855 52.025 113.705 ;
        RECT 52.755 113.015 54.755 113.185 ;
        RECT 55.045 113.015 57.045 113.185 ;
        RECT 52.525 104.760 52.695 112.800 ;
        RECT 54.815 104.760 54.985 112.800 ;
        RECT 57.105 104.760 57.275 112.800 ;
        RECT 52.755 104.375 54.755 104.545 ;
        RECT 55.045 104.375 57.045 104.545 ;
        RECT 57.775 103.855 57.945 113.705 ;
        RECT 58.675 113.015 60.675 113.185 ;
        RECT 60.965 113.015 62.965 113.185 ;
        RECT 58.445 104.760 58.615 112.800 ;
        RECT 60.735 104.760 60.905 112.800 ;
        RECT 63.025 104.760 63.195 112.800 ;
        RECT 58.675 104.375 60.675 104.545 ;
        RECT 60.965 104.375 62.965 104.545 ;
        RECT 63.695 103.855 63.865 113.705 ;
        RECT 64.595 113.015 66.595 113.185 ;
        RECT 66.885 113.015 68.885 113.185 ;
        RECT 64.365 104.760 64.535 112.800 ;
        RECT 66.655 104.760 66.825 112.800 ;
        RECT 68.945 104.760 69.115 112.800 ;
        RECT 64.595 104.375 66.595 104.545 ;
        RECT 66.885 104.375 68.885 104.545 ;
        RECT 69.615 103.855 70.145 113.705 ;
        RECT 10.055 103.325 70.145 103.855 ;
        RECT 71.805 123.725 114.135 124.255 ;
        RECT 138.110 124.120 145.930 124.650 ;
        RECT 71.805 113.875 72.335 123.725 ;
        RECT 72.835 122.820 77.585 123.725 ;
        RECT 72.835 114.780 73.005 122.820 ;
        RECT 75.125 114.780 75.295 122.820 ;
        RECT 77.415 114.780 77.585 122.820 ;
        RECT 73.065 114.395 75.065 114.565 ;
        RECT 75.355 114.395 77.355 114.565 ;
        RECT 78.085 113.875 78.255 123.725 ;
        RECT 78.985 123.035 80.985 123.205 ;
        RECT 81.275 123.035 83.275 123.205 ;
        RECT 78.755 114.780 78.925 122.820 ;
        RECT 81.045 114.780 81.215 122.820 ;
        RECT 83.335 114.780 83.505 122.820 ;
        RECT 78.985 114.395 80.985 114.565 ;
        RECT 81.275 114.395 83.275 114.565 ;
        RECT 84.005 113.875 84.175 123.725 ;
        RECT 84.905 123.035 86.905 123.205 ;
        RECT 87.195 123.035 89.195 123.205 ;
        RECT 84.675 114.780 84.845 122.820 ;
        RECT 86.965 114.780 87.135 122.820 ;
        RECT 89.255 114.780 89.425 122.820 ;
        RECT 84.905 114.395 86.905 114.565 ;
        RECT 87.195 114.395 89.195 114.565 ;
        RECT 89.925 113.875 90.095 123.725 ;
        RECT 90.825 123.035 92.825 123.205 ;
        RECT 93.115 123.035 95.115 123.205 ;
        RECT 90.595 114.780 90.765 122.820 ;
        RECT 92.885 114.780 93.055 122.820 ;
        RECT 95.175 114.780 95.345 122.820 ;
        RECT 90.825 114.395 92.825 114.565 ;
        RECT 93.115 114.395 95.115 114.565 ;
        RECT 95.845 113.875 96.015 123.725 ;
        RECT 96.745 123.035 98.745 123.205 ;
        RECT 99.035 123.035 101.035 123.205 ;
        RECT 96.515 114.780 96.685 122.820 ;
        RECT 98.805 114.780 98.975 122.820 ;
        RECT 101.095 114.780 101.265 122.820 ;
        RECT 96.745 114.395 98.745 114.565 ;
        RECT 99.035 114.395 101.035 114.565 ;
        RECT 101.765 113.875 101.935 123.725 ;
        RECT 102.665 123.035 104.665 123.205 ;
        RECT 104.955 123.035 106.955 123.205 ;
        RECT 102.435 114.780 102.605 122.820 ;
        RECT 104.725 114.780 104.895 122.820 ;
        RECT 107.015 114.780 107.185 122.820 ;
        RECT 102.665 114.395 104.665 114.565 ;
        RECT 104.955 114.395 106.955 114.565 ;
        RECT 107.685 113.875 107.855 123.725 ;
        RECT 108.355 122.820 113.105 123.725 ;
        RECT 108.355 114.780 108.525 122.820 ;
        RECT 110.645 114.780 110.815 122.820 ;
        RECT 112.935 114.780 113.105 122.820 ;
        RECT 108.585 114.395 110.585 114.565 ;
        RECT 110.875 114.395 112.875 114.565 ;
        RECT 113.605 113.875 114.135 123.725 ;
        RECT 71.805 113.705 114.135 113.875 ;
        RECT 71.805 103.855 72.335 113.705 ;
        RECT 73.065 113.015 75.065 113.185 ;
        RECT 75.355 113.015 77.355 113.185 ;
        RECT 72.835 104.760 73.005 112.800 ;
        RECT 75.125 104.760 75.295 112.800 ;
        RECT 77.415 104.760 77.585 112.800 ;
        RECT 72.835 103.855 77.585 104.760 ;
        RECT 78.085 103.855 78.255 113.705 ;
        RECT 78.985 113.015 80.985 113.185 ;
        RECT 81.275 113.015 83.275 113.185 ;
        RECT 78.755 104.760 78.925 112.800 ;
        RECT 81.045 104.760 81.215 112.800 ;
        RECT 83.335 104.760 83.505 112.800 ;
        RECT 78.985 104.375 80.985 104.545 ;
        RECT 81.275 104.375 83.275 104.545 ;
        RECT 84.005 103.855 84.175 113.705 ;
        RECT 84.905 113.015 86.905 113.185 ;
        RECT 87.195 113.015 89.195 113.185 ;
        RECT 84.675 104.760 84.845 112.800 ;
        RECT 86.965 104.760 87.135 112.800 ;
        RECT 89.255 104.760 89.425 112.800 ;
        RECT 84.905 104.375 86.905 104.545 ;
        RECT 87.195 104.375 89.195 104.545 ;
        RECT 89.925 103.855 90.095 113.705 ;
        RECT 90.825 113.015 92.825 113.185 ;
        RECT 93.115 113.015 95.115 113.185 ;
        RECT 90.595 104.760 90.765 112.800 ;
        RECT 92.885 104.760 93.055 112.800 ;
        RECT 95.175 104.760 95.345 112.800 ;
        RECT 90.825 104.375 92.825 104.545 ;
        RECT 93.115 104.375 95.115 104.545 ;
        RECT 95.845 103.855 96.015 113.705 ;
        RECT 96.745 113.015 98.745 113.185 ;
        RECT 99.035 113.015 101.035 113.185 ;
        RECT 96.515 104.760 96.685 112.800 ;
        RECT 98.805 104.760 98.975 112.800 ;
        RECT 101.095 104.760 101.265 112.800 ;
        RECT 96.745 104.375 98.745 104.545 ;
        RECT 99.035 104.375 101.035 104.545 ;
        RECT 101.765 103.855 101.935 113.705 ;
        RECT 102.665 113.015 104.665 113.185 ;
        RECT 104.955 113.015 106.955 113.185 ;
        RECT 102.435 104.760 102.605 112.800 ;
        RECT 104.725 104.760 104.895 112.800 ;
        RECT 107.015 104.760 107.185 112.800 ;
        RECT 102.665 104.375 104.665 104.545 ;
        RECT 104.955 104.375 106.955 104.545 ;
        RECT 107.685 103.855 107.855 113.705 ;
        RECT 108.585 113.015 110.585 113.185 ;
        RECT 110.875 113.015 112.875 113.185 ;
        RECT 108.355 104.760 108.525 112.800 ;
        RECT 110.645 104.760 110.815 112.800 ;
        RECT 112.935 104.760 113.105 112.800 ;
        RECT 108.355 103.855 113.105 104.760 ;
        RECT 113.605 103.855 114.135 113.705 ;
        RECT 71.805 103.325 114.135 103.855 ;
        RECT 115.935 122.945 128.905 123.475 ;
        RECT 115.935 113.485 116.465 122.945 ;
        RECT 117.370 122.275 118.410 122.445 ;
        RECT 116.985 114.215 117.155 122.215 ;
        RECT 118.625 114.215 118.795 122.215 ;
        RECT 117.370 113.985 118.410 114.155 ;
        RECT 119.315 113.485 119.485 122.945 ;
        RECT 120.390 122.275 121.430 122.445 ;
        RECT 120.005 114.215 120.175 122.215 ;
        RECT 121.645 114.215 121.815 122.215 ;
        RECT 120.390 113.985 121.430 114.155 ;
        RECT 122.335 113.485 122.505 122.945 ;
        RECT 123.410 122.275 124.450 122.445 ;
        RECT 123.025 114.215 123.195 122.215 ;
        RECT 124.665 114.215 124.835 122.215 ;
        RECT 123.410 113.985 124.450 114.155 ;
        RECT 125.355 113.485 125.525 122.945 ;
        RECT 126.430 122.275 127.470 122.445 ;
        RECT 126.045 114.215 126.215 122.215 ;
        RECT 127.685 114.215 127.855 122.215 ;
        RECT 126.430 113.985 127.470 114.155 ;
        RECT 128.375 113.485 128.905 122.945 ;
        RECT 115.935 113.315 128.905 113.485 ;
        RECT 115.935 103.855 116.465 113.315 ;
        RECT 117.370 112.645 118.410 112.815 ;
        RECT 116.985 104.585 117.155 112.585 ;
        RECT 118.625 104.585 118.795 112.585 ;
        RECT 117.370 104.355 118.410 104.525 ;
        RECT 119.315 103.855 119.485 113.315 ;
        RECT 120.390 112.645 121.430 112.815 ;
        RECT 120.005 104.585 120.175 112.585 ;
        RECT 121.645 104.585 121.815 112.585 ;
        RECT 120.390 104.355 121.430 104.525 ;
        RECT 122.335 103.855 122.505 113.315 ;
        RECT 123.410 112.645 124.450 112.815 ;
        RECT 123.025 104.585 123.195 112.585 ;
        RECT 124.665 104.585 124.835 112.585 ;
        RECT 123.410 104.355 124.450 104.525 ;
        RECT 125.355 103.855 125.525 113.315 ;
        RECT 126.430 112.645 127.470 112.815 ;
        RECT 126.045 104.585 126.215 112.585 ;
        RECT 127.685 104.585 127.855 112.585 ;
        RECT 126.430 104.355 127.470 104.525 ;
        RECT 128.375 103.855 128.905 113.315 ;
        RECT 115.935 103.325 128.905 103.855 ;
        RECT 135.150 104.785 149.540 108.660 ;
        RECT 10.055 102.145 128.905 102.675 ;
        RECT 10.055 92.295 10.585 102.145 ;
        RECT 11.315 101.455 13.315 101.625 ;
        RECT 13.605 101.455 15.605 101.625 ;
        RECT 15.895 101.455 17.895 101.625 ;
        RECT 18.185 101.455 20.185 101.625 ;
        RECT 20.475 101.455 22.475 101.625 ;
        RECT 22.765 101.455 24.765 101.625 ;
        RECT 25.055 101.455 27.055 101.625 ;
        RECT 27.345 101.455 29.345 101.625 ;
        RECT 11.085 93.200 11.255 101.240 ;
        RECT 13.375 93.200 13.545 101.240 ;
        RECT 15.665 93.200 15.835 101.240 ;
        RECT 17.955 93.200 18.125 101.240 ;
        RECT 20.245 93.200 20.415 101.240 ;
        RECT 22.535 93.200 22.705 101.240 ;
        RECT 24.825 93.200 24.995 101.240 ;
        RECT 27.115 93.200 27.285 101.240 ;
        RECT 29.405 93.200 29.575 101.240 ;
        RECT 11.315 92.815 13.315 92.985 ;
        RECT 13.605 92.815 15.605 92.985 ;
        RECT 15.895 92.815 17.895 92.985 ;
        RECT 18.185 92.815 20.185 92.985 ;
        RECT 20.475 92.815 22.475 92.985 ;
        RECT 22.765 92.815 24.765 92.985 ;
        RECT 25.055 92.815 27.055 92.985 ;
        RECT 27.345 92.815 29.345 92.985 ;
        RECT 30.075 92.295 30.245 102.145 ;
        RECT 30.975 101.455 32.975 101.625 ;
        RECT 33.265 101.455 35.265 101.625 ;
        RECT 35.555 101.455 37.555 101.625 ;
        RECT 37.845 101.455 39.845 101.625 ;
        RECT 40.135 101.455 42.135 101.625 ;
        RECT 42.425 101.455 44.425 101.625 ;
        RECT 44.715 101.455 46.715 101.625 ;
        RECT 47.005 101.455 49.005 101.625 ;
        RECT 30.745 93.200 30.915 101.240 ;
        RECT 33.035 93.200 33.205 101.240 ;
        RECT 35.325 93.200 35.495 101.240 ;
        RECT 37.615 93.200 37.785 101.240 ;
        RECT 39.905 93.200 40.075 101.240 ;
        RECT 42.195 93.200 42.365 101.240 ;
        RECT 44.485 93.200 44.655 101.240 ;
        RECT 46.775 93.200 46.945 101.240 ;
        RECT 49.065 93.200 49.235 101.240 ;
        RECT 30.975 92.815 32.975 92.985 ;
        RECT 33.265 92.815 35.265 92.985 ;
        RECT 35.555 92.815 37.555 92.985 ;
        RECT 37.845 92.815 39.845 92.985 ;
        RECT 40.135 92.815 42.135 92.985 ;
        RECT 42.425 92.815 44.425 92.985 ;
        RECT 44.715 92.815 46.715 92.985 ;
        RECT 47.005 92.815 49.005 92.985 ;
        RECT 49.735 92.295 49.905 102.145 ;
        RECT 50.635 101.455 52.635 101.625 ;
        RECT 52.925 101.455 54.925 101.625 ;
        RECT 55.215 101.455 57.215 101.625 ;
        RECT 57.505 101.455 59.505 101.625 ;
        RECT 59.795 101.455 61.795 101.625 ;
        RECT 62.085 101.455 64.085 101.625 ;
        RECT 64.375 101.455 66.375 101.625 ;
        RECT 66.665 101.455 68.665 101.625 ;
        RECT 50.405 93.200 50.575 101.240 ;
        RECT 52.695 93.200 52.865 101.240 ;
        RECT 54.985 93.200 55.155 101.240 ;
        RECT 57.275 93.200 57.445 101.240 ;
        RECT 59.565 93.200 59.735 101.240 ;
        RECT 61.855 93.200 62.025 101.240 ;
        RECT 64.145 93.200 64.315 101.240 ;
        RECT 66.435 93.200 66.605 101.240 ;
        RECT 68.725 93.200 68.895 101.240 ;
        RECT 50.635 92.815 52.635 92.985 ;
        RECT 52.925 92.815 54.925 92.985 ;
        RECT 55.215 92.815 57.215 92.985 ;
        RECT 57.505 92.815 59.505 92.985 ;
        RECT 59.795 92.815 61.795 92.985 ;
        RECT 62.085 92.815 64.085 92.985 ;
        RECT 64.375 92.815 66.375 92.985 ;
        RECT 66.665 92.815 68.665 92.985 ;
        RECT 69.395 92.295 69.565 102.145 ;
        RECT 70.295 101.455 72.295 101.625 ;
        RECT 72.585 101.455 74.585 101.625 ;
        RECT 74.875 101.455 76.875 101.625 ;
        RECT 77.165 101.455 79.165 101.625 ;
        RECT 79.455 101.455 81.455 101.625 ;
        RECT 81.745 101.455 83.745 101.625 ;
        RECT 84.035 101.455 86.035 101.625 ;
        RECT 86.325 101.455 88.325 101.625 ;
        RECT 70.065 93.200 70.235 101.240 ;
        RECT 72.355 93.200 72.525 101.240 ;
        RECT 74.645 93.200 74.815 101.240 ;
        RECT 76.935 93.200 77.105 101.240 ;
        RECT 79.225 93.200 79.395 101.240 ;
        RECT 81.515 93.200 81.685 101.240 ;
        RECT 83.805 93.200 83.975 101.240 ;
        RECT 86.095 93.200 86.265 101.240 ;
        RECT 88.385 93.200 88.555 101.240 ;
        RECT 70.295 92.815 72.295 92.985 ;
        RECT 72.585 92.815 74.585 92.985 ;
        RECT 74.875 92.815 76.875 92.985 ;
        RECT 77.165 92.815 79.165 92.985 ;
        RECT 79.455 92.815 81.455 92.985 ;
        RECT 81.745 92.815 83.745 92.985 ;
        RECT 84.035 92.815 86.035 92.985 ;
        RECT 86.325 92.815 88.325 92.985 ;
        RECT 89.055 92.295 89.225 102.145 ;
        RECT 89.955 101.455 91.955 101.625 ;
        RECT 92.245 101.455 94.245 101.625 ;
        RECT 94.535 101.455 96.535 101.625 ;
        RECT 96.825 101.455 98.825 101.625 ;
        RECT 99.115 101.455 101.115 101.625 ;
        RECT 101.405 101.455 103.405 101.625 ;
        RECT 103.695 101.455 105.695 101.625 ;
        RECT 105.985 101.455 107.985 101.625 ;
        RECT 89.725 93.200 89.895 101.240 ;
        RECT 92.015 93.200 92.185 101.240 ;
        RECT 94.305 93.200 94.475 101.240 ;
        RECT 96.595 93.200 96.765 101.240 ;
        RECT 98.885 93.200 99.055 101.240 ;
        RECT 101.175 93.200 101.345 101.240 ;
        RECT 103.465 93.200 103.635 101.240 ;
        RECT 105.755 93.200 105.925 101.240 ;
        RECT 108.045 93.200 108.215 101.240 ;
        RECT 89.955 92.815 91.955 92.985 ;
        RECT 92.245 92.815 94.245 92.985 ;
        RECT 94.535 92.815 96.535 92.985 ;
        RECT 96.825 92.815 98.825 92.985 ;
        RECT 99.115 92.815 101.115 92.985 ;
        RECT 101.405 92.815 103.405 92.985 ;
        RECT 103.695 92.815 105.695 92.985 ;
        RECT 105.985 92.815 107.985 92.985 ;
        RECT 108.715 92.295 108.885 102.145 ;
        RECT 109.615 101.455 111.615 101.625 ;
        RECT 111.905 101.455 113.905 101.625 ;
        RECT 114.195 101.455 116.195 101.625 ;
        RECT 116.485 101.455 118.485 101.625 ;
        RECT 118.775 101.455 120.775 101.625 ;
        RECT 121.065 101.455 123.065 101.625 ;
        RECT 123.355 101.455 125.355 101.625 ;
        RECT 125.645 101.455 127.645 101.625 ;
        RECT 109.385 93.200 109.555 101.240 ;
        RECT 111.675 93.200 111.845 101.240 ;
        RECT 113.965 93.200 114.135 101.240 ;
        RECT 116.255 93.200 116.425 101.240 ;
        RECT 118.545 93.200 118.715 101.240 ;
        RECT 120.835 93.200 121.005 101.240 ;
        RECT 123.125 93.200 123.295 101.240 ;
        RECT 125.415 93.200 125.585 101.240 ;
        RECT 127.705 93.200 127.875 101.240 ;
        RECT 109.615 92.815 111.615 92.985 ;
        RECT 111.905 92.815 113.905 92.985 ;
        RECT 114.195 92.815 116.195 92.985 ;
        RECT 116.485 92.815 118.485 92.985 ;
        RECT 118.775 92.815 120.775 92.985 ;
        RECT 121.065 92.815 123.065 92.985 ;
        RECT 123.355 92.815 125.355 92.985 ;
        RECT 125.645 92.815 127.645 92.985 ;
        RECT 128.375 92.295 128.905 102.145 ;
        RECT 10.055 92.125 128.905 92.295 ;
        RECT 10.055 82.275 10.585 92.125 ;
        RECT 11.315 91.435 13.315 91.605 ;
        RECT 13.605 91.435 15.605 91.605 ;
        RECT 15.895 91.435 17.895 91.605 ;
        RECT 18.185 91.435 20.185 91.605 ;
        RECT 20.475 91.435 22.475 91.605 ;
        RECT 22.765 91.435 24.765 91.605 ;
        RECT 25.055 91.435 27.055 91.605 ;
        RECT 27.345 91.435 29.345 91.605 ;
        RECT 11.085 83.180 11.255 91.220 ;
        RECT 13.375 83.180 13.545 91.220 ;
        RECT 15.665 83.180 15.835 91.220 ;
        RECT 17.955 83.180 18.125 91.220 ;
        RECT 20.245 83.180 20.415 91.220 ;
        RECT 22.535 83.180 22.705 91.220 ;
        RECT 24.825 83.180 24.995 91.220 ;
        RECT 27.115 83.180 27.285 91.220 ;
        RECT 29.405 83.180 29.575 91.220 ;
        RECT 11.315 82.795 13.315 82.965 ;
        RECT 13.605 82.795 15.605 82.965 ;
        RECT 15.895 82.795 17.895 82.965 ;
        RECT 18.185 82.795 20.185 82.965 ;
        RECT 20.475 82.795 22.475 82.965 ;
        RECT 22.765 82.795 24.765 82.965 ;
        RECT 25.055 82.795 27.055 82.965 ;
        RECT 27.345 82.795 29.345 82.965 ;
        RECT 30.075 82.275 30.245 92.125 ;
        RECT 30.975 91.435 32.975 91.605 ;
        RECT 33.265 91.435 35.265 91.605 ;
        RECT 35.555 91.435 37.555 91.605 ;
        RECT 37.845 91.435 39.845 91.605 ;
        RECT 40.135 91.435 42.135 91.605 ;
        RECT 42.425 91.435 44.425 91.605 ;
        RECT 44.715 91.435 46.715 91.605 ;
        RECT 47.005 91.435 49.005 91.605 ;
        RECT 30.745 83.180 30.915 91.220 ;
        RECT 33.035 83.180 33.205 91.220 ;
        RECT 35.325 83.180 35.495 91.220 ;
        RECT 37.615 83.180 37.785 91.220 ;
        RECT 39.905 83.180 40.075 91.220 ;
        RECT 42.195 83.180 42.365 91.220 ;
        RECT 44.485 83.180 44.655 91.220 ;
        RECT 46.775 83.180 46.945 91.220 ;
        RECT 49.065 83.180 49.235 91.220 ;
        RECT 30.975 82.795 32.975 82.965 ;
        RECT 33.265 82.795 35.265 82.965 ;
        RECT 35.555 82.795 37.555 82.965 ;
        RECT 37.845 82.795 39.845 82.965 ;
        RECT 40.135 82.795 42.135 82.965 ;
        RECT 42.425 82.795 44.425 82.965 ;
        RECT 44.715 82.795 46.715 82.965 ;
        RECT 47.005 82.795 49.005 82.965 ;
        RECT 49.735 82.275 49.905 92.125 ;
        RECT 50.635 91.435 52.635 91.605 ;
        RECT 52.925 91.435 54.925 91.605 ;
        RECT 55.215 91.435 57.215 91.605 ;
        RECT 57.505 91.435 59.505 91.605 ;
        RECT 59.795 91.435 61.795 91.605 ;
        RECT 62.085 91.435 64.085 91.605 ;
        RECT 64.375 91.435 66.375 91.605 ;
        RECT 66.665 91.435 68.665 91.605 ;
        RECT 50.405 83.180 50.575 91.220 ;
        RECT 52.695 83.180 52.865 91.220 ;
        RECT 54.985 83.180 55.155 91.220 ;
        RECT 57.275 83.180 57.445 91.220 ;
        RECT 59.565 83.180 59.735 91.220 ;
        RECT 61.855 83.180 62.025 91.220 ;
        RECT 64.145 83.180 64.315 91.220 ;
        RECT 66.435 83.180 66.605 91.220 ;
        RECT 68.725 83.180 68.895 91.220 ;
        RECT 50.635 82.795 52.635 82.965 ;
        RECT 52.925 82.795 54.925 82.965 ;
        RECT 55.215 82.795 57.215 82.965 ;
        RECT 57.505 82.795 59.505 82.965 ;
        RECT 59.795 82.795 61.795 82.965 ;
        RECT 62.085 82.795 64.085 82.965 ;
        RECT 64.375 82.795 66.375 82.965 ;
        RECT 66.665 82.795 68.665 82.965 ;
        RECT 69.395 82.275 69.565 92.125 ;
        RECT 70.295 91.435 72.295 91.605 ;
        RECT 72.585 91.435 74.585 91.605 ;
        RECT 74.875 91.435 76.875 91.605 ;
        RECT 77.165 91.435 79.165 91.605 ;
        RECT 79.455 91.435 81.455 91.605 ;
        RECT 81.745 91.435 83.745 91.605 ;
        RECT 84.035 91.435 86.035 91.605 ;
        RECT 86.325 91.435 88.325 91.605 ;
        RECT 70.065 83.180 70.235 91.220 ;
        RECT 72.355 83.180 72.525 91.220 ;
        RECT 74.645 83.180 74.815 91.220 ;
        RECT 76.935 83.180 77.105 91.220 ;
        RECT 79.225 83.180 79.395 91.220 ;
        RECT 81.515 83.180 81.685 91.220 ;
        RECT 83.805 83.180 83.975 91.220 ;
        RECT 86.095 83.180 86.265 91.220 ;
        RECT 88.385 83.180 88.555 91.220 ;
        RECT 70.295 82.795 72.295 82.965 ;
        RECT 72.585 82.795 74.585 82.965 ;
        RECT 74.875 82.795 76.875 82.965 ;
        RECT 77.165 82.795 79.165 82.965 ;
        RECT 79.455 82.795 81.455 82.965 ;
        RECT 81.745 82.795 83.745 82.965 ;
        RECT 84.035 82.795 86.035 82.965 ;
        RECT 86.325 82.795 88.325 82.965 ;
        RECT 89.055 82.275 89.225 92.125 ;
        RECT 89.955 91.435 91.955 91.605 ;
        RECT 92.245 91.435 94.245 91.605 ;
        RECT 94.535 91.435 96.535 91.605 ;
        RECT 96.825 91.435 98.825 91.605 ;
        RECT 99.115 91.435 101.115 91.605 ;
        RECT 101.405 91.435 103.405 91.605 ;
        RECT 103.695 91.435 105.695 91.605 ;
        RECT 105.985 91.435 107.985 91.605 ;
        RECT 89.725 83.180 89.895 91.220 ;
        RECT 92.015 83.180 92.185 91.220 ;
        RECT 94.305 83.180 94.475 91.220 ;
        RECT 96.595 83.180 96.765 91.220 ;
        RECT 98.885 83.180 99.055 91.220 ;
        RECT 101.175 83.180 101.345 91.220 ;
        RECT 103.465 83.180 103.635 91.220 ;
        RECT 105.755 83.180 105.925 91.220 ;
        RECT 108.045 83.180 108.215 91.220 ;
        RECT 89.955 82.795 91.955 82.965 ;
        RECT 92.245 82.795 94.245 82.965 ;
        RECT 94.535 82.795 96.535 82.965 ;
        RECT 96.825 82.795 98.825 82.965 ;
        RECT 99.115 82.795 101.115 82.965 ;
        RECT 101.405 82.795 103.405 82.965 ;
        RECT 103.695 82.795 105.695 82.965 ;
        RECT 105.985 82.795 107.985 82.965 ;
        RECT 108.715 82.275 108.885 92.125 ;
        RECT 109.615 91.435 111.615 91.605 ;
        RECT 111.905 91.435 113.905 91.605 ;
        RECT 114.195 91.435 116.195 91.605 ;
        RECT 116.485 91.435 118.485 91.605 ;
        RECT 118.775 91.435 120.775 91.605 ;
        RECT 121.065 91.435 123.065 91.605 ;
        RECT 123.355 91.435 125.355 91.605 ;
        RECT 125.645 91.435 127.645 91.605 ;
        RECT 109.385 83.180 109.555 91.220 ;
        RECT 111.675 83.180 111.845 91.220 ;
        RECT 113.965 83.180 114.135 91.220 ;
        RECT 116.255 83.180 116.425 91.220 ;
        RECT 118.545 83.180 118.715 91.220 ;
        RECT 120.835 83.180 121.005 91.220 ;
        RECT 123.125 83.180 123.295 91.220 ;
        RECT 125.415 83.180 125.585 91.220 ;
        RECT 127.705 83.180 127.875 91.220 ;
        RECT 109.615 82.795 111.615 82.965 ;
        RECT 111.905 82.795 113.905 82.965 ;
        RECT 114.195 82.795 116.195 82.965 ;
        RECT 116.485 82.795 118.485 82.965 ;
        RECT 118.775 82.795 120.775 82.965 ;
        RECT 121.065 82.795 123.065 82.965 ;
        RECT 123.355 82.795 125.355 82.965 ;
        RECT 125.645 82.795 127.645 82.965 ;
        RECT 128.375 82.275 128.905 92.125 ;
        RECT 10.055 82.105 128.905 82.275 ;
        RECT 10.055 72.255 10.585 82.105 ;
        RECT 11.315 81.415 13.315 81.585 ;
        RECT 13.605 81.415 15.605 81.585 ;
        RECT 15.895 81.415 17.895 81.585 ;
        RECT 18.185 81.415 20.185 81.585 ;
        RECT 20.475 81.415 22.475 81.585 ;
        RECT 22.765 81.415 24.765 81.585 ;
        RECT 25.055 81.415 27.055 81.585 ;
        RECT 27.345 81.415 29.345 81.585 ;
        RECT 11.085 73.160 11.255 81.200 ;
        RECT 13.375 73.160 13.545 81.200 ;
        RECT 15.665 73.160 15.835 81.200 ;
        RECT 17.955 73.160 18.125 81.200 ;
        RECT 20.245 73.160 20.415 81.200 ;
        RECT 22.535 73.160 22.705 81.200 ;
        RECT 24.825 73.160 24.995 81.200 ;
        RECT 27.115 73.160 27.285 81.200 ;
        RECT 29.405 73.160 29.575 81.200 ;
        RECT 11.315 72.775 13.315 72.945 ;
        RECT 13.605 72.775 15.605 72.945 ;
        RECT 15.895 72.775 17.895 72.945 ;
        RECT 18.185 72.775 20.185 72.945 ;
        RECT 20.475 72.775 22.475 72.945 ;
        RECT 22.765 72.775 24.765 72.945 ;
        RECT 25.055 72.775 27.055 72.945 ;
        RECT 27.345 72.775 29.345 72.945 ;
        RECT 30.075 72.255 30.245 82.105 ;
        RECT 30.975 81.415 32.975 81.585 ;
        RECT 33.265 81.415 35.265 81.585 ;
        RECT 35.555 81.415 37.555 81.585 ;
        RECT 37.845 81.415 39.845 81.585 ;
        RECT 40.135 81.415 42.135 81.585 ;
        RECT 42.425 81.415 44.425 81.585 ;
        RECT 44.715 81.415 46.715 81.585 ;
        RECT 47.005 81.415 49.005 81.585 ;
        RECT 30.745 73.160 30.915 81.200 ;
        RECT 33.035 73.160 33.205 81.200 ;
        RECT 35.325 73.160 35.495 81.200 ;
        RECT 37.615 73.160 37.785 81.200 ;
        RECT 39.905 73.160 40.075 81.200 ;
        RECT 42.195 73.160 42.365 81.200 ;
        RECT 44.485 73.160 44.655 81.200 ;
        RECT 46.775 73.160 46.945 81.200 ;
        RECT 49.065 73.160 49.235 81.200 ;
        RECT 30.975 72.775 32.975 72.945 ;
        RECT 33.265 72.775 35.265 72.945 ;
        RECT 35.555 72.775 37.555 72.945 ;
        RECT 37.845 72.775 39.845 72.945 ;
        RECT 40.135 72.775 42.135 72.945 ;
        RECT 42.425 72.775 44.425 72.945 ;
        RECT 44.715 72.775 46.715 72.945 ;
        RECT 47.005 72.775 49.005 72.945 ;
        RECT 49.735 72.255 49.905 82.105 ;
        RECT 50.635 81.415 52.635 81.585 ;
        RECT 52.925 81.415 54.925 81.585 ;
        RECT 55.215 81.415 57.215 81.585 ;
        RECT 57.505 81.415 59.505 81.585 ;
        RECT 59.795 81.415 61.795 81.585 ;
        RECT 62.085 81.415 64.085 81.585 ;
        RECT 64.375 81.415 66.375 81.585 ;
        RECT 66.665 81.415 68.665 81.585 ;
        RECT 50.405 73.160 50.575 81.200 ;
        RECT 52.695 73.160 52.865 81.200 ;
        RECT 54.985 73.160 55.155 81.200 ;
        RECT 57.275 73.160 57.445 81.200 ;
        RECT 59.565 73.160 59.735 81.200 ;
        RECT 61.855 73.160 62.025 81.200 ;
        RECT 64.145 73.160 64.315 81.200 ;
        RECT 66.435 73.160 66.605 81.200 ;
        RECT 68.725 73.160 68.895 81.200 ;
        RECT 50.635 72.775 52.635 72.945 ;
        RECT 52.925 72.775 54.925 72.945 ;
        RECT 55.215 72.775 57.215 72.945 ;
        RECT 57.505 72.775 59.505 72.945 ;
        RECT 59.795 72.775 61.795 72.945 ;
        RECT 62.085 72.775 64.085 72.945 ;
        RECT 64.375 72.775 66.375 72.945 ;
        RECT 66.665 72.775 68.665 72.945 ;
        RECT 69.395 72.255 69.565 82.105 ;
        RECT 70.295 81.415 72.295 81.585 ;
        RECT 72.585 81.415 74.585 81.585 ;
        RECT 74.875 81.415 76.875 81.585 ;
        RECT 77.165 81.415 79.165 81.585 ;
        RECT 79.455 81.415 81.455 81.585 ;
        RECT 81.745 81.415 83.745 81.585 ;
        RECT 84.035 81.415 86.035 81.585 ;
        RECT 86.325 81.415 88.325 81.585 ;
        RECT 70.065 73.160 70.235 81.200 ;
        RECT 72.355 73.160 72.525 81.200 ;
        RECT 74.645 73.160 74.815 81.200 ;
        RECT 76.935 73.160 77.105 81.200 ;
        RECT 79.225 73.160 79.395 81.200 ;
        RECT 81.515 73.160 81.685 81.200 ;
        RECT 83.805 73.160 83.975 81.200 ;
        RECT 86.095 73.160 86.265 81.200 ;
        RECT 88.385 73.160 88.555 81.200 ;
        RECT 70.295 72.775 72.295 72.945 ;
        RECT 72.585 72.775 74.585 72.945 ;
        RECT 74.875 72.775 76.875 72.945 ;
        RECT 77.165 72.775 79.165 72.945 ;
        RECT 79.455 72.775 81.455 72.945 ;
        RECT 81.745 72.775 83.745 72.945 ;
        RECT 84.035 72.775 86.035 72.945 ;
        RECT 86.325 72.775 88.325 72.945 ;
        RECT 89.055 72.255 89.225 82.105 ;
        RECT 89.955 81.415 91.955 81.585 ;
        RECT 92.245 81.415 94.245 81.585 ;
        RECT 94.535 81.415 96.535 81.585 ;
        RECT 96.825 81.415 98.825 81.585 ;
        RECT 99.115 81.415 101.115 81.585 ;
        RECT 101.405 81.415 103.405 81.585 ;
        RECT 103.695 81.415 105.695 81.585 ;
        RECT 105.985 81.415 107.985 81.585 ;
        RECT 89.725 73.160 89.895 81.200 ;
        RECT 92.015 73.160 92.185 81.200 ;
        RECT 94.305 73.160 94.475 81.200 ;
        RECT 96.595 73.160 96.765 81.200 ;
        RECT 98.885 73.160 99.055 81.200 ;
        RECT 101.175 73.160 101.345 81.200 ;
        RECT 103.465 73.160 103.635 81.200 ;
        RECT 105.755 73.160 105.925 81.200 ;
        RECT 108.045 73.160 108.215 81.200 ;
        RECT 89.955 72.775 91.955 72.945 ;
        RECT 92.245 72.775 94.245 72.945 ;
        RECT 94.535 72.775 96.535 72.945 ;
        RECT 96.825 72.775 98.825 72.945 ;
        RECT 99.115 72.775 101.115 72.945 ;
        RECT 101.405 72.775 103.405 72.945 ;
        RECT 103.695 72.775 105.695 72.945 ;
        RECT 105.985 72.775 107.985 72.945 ;
        RECT 108.715 72.255 108.885 82.105 ;
        RECT 109.615 81.415 111.615 81.585 ;
        RECT 111.905 81.415 113.905 81.585 ;
        RECT 114.195 81.415 116.195 81.585 ;
        RECT 116.485 81.415 118.485 81.585 ;
        RECT 118.775 81.415 120.775 81.585 ;
        RECT 121.065 81.415 123.065 81.585 ;
        RECT 123.355 81.415 125.355 81.585 ;
        RECT 125.645 81.415 127.645 81.585 ;
        RECT 109.385 73.160 109.555 81.200 ;
        RECT 111.675 73.160 111.845 81.200 ;
        RECT 113.965 73.160 114.135 81.200 ;
        RECT 116.255 73.160 116.425 81.200 ;
        RECT 118.545 73.160 118.715 81.200 ;
        RECT 120.835 73.160 121.005 81.200 ;
        RECT 123.125 73.160 123.295 81.200 ;
        RECT 125.415 73.160 125.585 81.200 ;
        RECT 127.705 73.160 127.875 81.200 ;
        RECT 109.615 72.775 111.615 72.945 ;
        RECT 111.905 72.775 113.905 72.945 ;
        RECT 114.195 72.775 116.195 72.945 ;
        RECT 116.485 72.775 118.485 72.945 ;
        RECT 118.775 72.775 120.775 72.945 ;
        RECT 121.065 72.775 123.065 72.945 ;
        RECT 123.355 72.775 125.355 72.945 ;
        RECT 125.645 72.775 127.645 72.945 ;
        RECT 128.375 72.255 128.905 82.105 ;
        RECT 10.055 72.085 128.905 72.255 ;
        RECT 10.055 62.235 10.585 72.085 ;
        RECT 11.315 71.395 13.315 71.565 ;
        RECT 13.605 71.395 15.605 71.565 ;
        RECT 15.895 71.395 17.895 71.565 ;
        RECT 18.185 71.395 20.185 71.565 ;
        RECT 20.475 71.395 22.475 71.565 ;
        RECT 22.765 71.395 24.765 71.565 ;
        RECT 25.055 71.395 27.055 71.565 ;
        RECT 27.345 71.395 29.345 71.565 ;
        RECT 11.085 63.140 11.255 71.180 ;
        RECT 13.375 63.140 13.545 71.180 ;
        RECT 15.665 63.140 15.835 71.180 ;
        RECT 17.955 63.140 18.125 71.180 ;
        RECT 20.245 63.140 20.415 71.180 ;
        RECT 22.535 63.140 22.705 71.180 ;
        RECT 24.825 63.140 24.995 71.180 ;
        RECT 27.115 63.140 27.285 71.180 ;
        RECT 29.405 63.140 29.575 71.180 ;
        RECT 11.315 62.755 13.315 62.925 ;
        RECT 13.605 62.755 15.605 62.925 ;
        RECT 15.895 62.755 17.895 62.925 ;
        RECT 18.185 62.755 20.185 62.925 ;
        RECT 20.475 62.755 22.475 62.925 ;
        RECT 22.765 62.755 24.765 62.925 ;
        RECT 25.055 62.755 27.055 62.925 ;
        RECT 27.345 62.755 29.345 62.925 ;
        RECT 30.075 62.235 30.245 72.085 ;
        RECT 30.975 71.395 32.975 71.565 ;
        RECT 33.265 71.395 35.265 71.565 ;
        RECT 35.555 71.395 37.555 71.565 ;
        RECT 37.845 71.395 39.845 71.565 ;
        RECT 40.135 71.395 42.135 71.565 ;
        RECT 42.425 71.395 44.425 71.565 ;
        RECT 44.715 71.395 46.715 71.565 ;
        RECT 47.005 71.395 49.005 71.565 ;
        RECT 30.745 63.140 30.915 71.180 ;
        RECT 33.035 63.140 33.205 71.180 ;
        RECT 35.325 63.140 35.495 71.180 ;
        RECT 37.615 63.140 37.785 71.180 ;
        RECT 39.905 63.140 40.075 71.180 ;
        RECT 42.195 63.140 42.365 71.180 ;
        RECT 44.485 63.140 44.655 71.180 ;
        RECT 46.775 63.140 46.945 71.180 ;
        RECT 49.065 63.140 49.235 71.180 ;
        RECT 30.975 62.755 32.975 62.925 ;
        RECT 33.265 62.755 35.265 62.925 ;
        RECT 35.555 62.755 37.555 62.925 ;
        RECT 37.845 62.755 39.845 62.925 ;
        RECT 40.135 62.755 42.135 62.925 ;
        RECT 42.425 62.755 44.425 62.925 ;
        RECT 44.715 62.755 46.715 62.925 ;
        RECT 47.005 62.755 49.005 62.925 ;
        RECT 49.735 62.235 49.905 72.085 ;
        RECT 50.635 71.395 52.635 71.565 ;
        RECT 52.925 71.395 54.925 71.565 ;
        RECT 55.215 71.395 57.215 71.565 ;
        RECT 57.505 71.395 59.505 71.565 ;
        RECT 59.795 71.395 61.795 71.565 ;
        RECT 62.085 71.395 64.085 71.565 ;
        RECT 64.375 71.395 66.375 71.565 ;
        RECT 66.665 71.395 68.665 71.565 ;
        RECT 50.405 63.140 50.575 71.180 ;
        RECT 52.695 63.140 52.865 71.180 ;
        RECT 54.985 63.140 55.155 71.180 ;
        RECT 57.275 63.140 57.445 71.180 ;
        RECT 59.565 63.140 59.735 71.180 ;
        RECT 61.855 63.140 62.025 71.180 ;
        RECT 64.145 63.140 64.315 71.180 ;
        RECT 66.435 63.140 66.605 71.180 ;
        RECT 68.725 63.140 68.895 71.180 ;
        RECT 50.635 62.755 52.635 62.925 ;
        RECT 52.925 62.755 54.925 62.925 ;
        RECT 55.215 62.755 57.215 62.925 ;
        RECT 57.505 62.755 59.505 62.925 ;
        RECT 59.795 62.755 61.795 62.925 ;
        RECT 62.085 62.755 64.085 62.925 ;
        RECT 64.375 62.755 66.375 62.925 ;
        RECT 66.665 62.755 68.665 62.925 ;
        RECT 69.395 62.235 69.565 72.085 ;
        RECT 70.295 71.395 72.295 71.565 ;
        RECT 72.585 71.395 74.585 71.565 ;
        RECT 74.875 71.395 76.875 71.565 ;
        RECT 77.165 71.395 79.165 71.565 ;
        RECT 79.455 71.395 81.455 71.565 ;
        RECT 81.745 71.395 83.745 71.565 ;
        RECT 84.035 71.395 86.035 71.565 ;
        RECT 86.325 71.395 88.325 71.565 ;
        RECT 70.065 63.140 70.235 71.180 ;
        RECT 72.355 63.140 72.525 71.180 ;
        RECT 74.645 63.140 74.815 71.180 ;
        RECT 76.935 63.140 77.105 71.180 ;
        RECT 79.225 63.140 79.395 71.180 ;
        RECT 81.515 63.140 81.685 71.180 ;
        RECT 83.805 63.140 83.975 71.180 ;
        RECT 86.095 63.140 86.265 71.180 ;
        RECT 88.385 63.140 88.555 71.180 ;
        RECT 70.295 62.755 72.295 62.925 ;
        RECT 72.585 62.755 74.585 62.925 ;
        RECT 74.875 62.755 76.875 62.925 ;
        RECT 77.165 62.755 79.165 62.925 ;
        RECT 79.455 62.755 81.455 62.925 ;
        RECT 81.745 62.755 83.745 62.925 ;
        RECT 84.035 62.755 86.035 62.925 ;
        RECT 86.325 62.755 88.325 62.925 ;
        RECT 89.055 62.235 89.225 72.085 ;
        RECT 89.955 71.395 91.955 71.565 ;
        RECT 92.245 71.395 94.245 71.565 ;
        RECT 94.535 71.395 96.535 71.565 ;
        RECT 96.825 71.395 98.825 71.565 ;
        RECT 99.115 71.395 101.115 71.565 ;
        RECT 101.405 71.395 103.405 71.565 ;
        RECT 103.695 71.395 105.695 71.565 ;
        RECT 105.985 71.395 107.985 71.565 ;
        RECT 89.725 63.140 89.895 71.180 ;
        RECT 92.015 63.140 92.185 71.180 ;
        RECT 94.305 63.140 94.475 71.180 ;
        RECT 96.595 63.140 96.765 71.180 ;
        RECT 98.885 63.140 99.055 71.180 ;
        RECT 101.175 63.140 101.345 71.180 ;
        RECT 103.465 63.140 103.635 71.180 ;
        RECT 105.755 63.140 105.925 71.180 ;
        RECT 108.045 63.140 108.215 71.180 ;
        RECT 89.955 62.755 91.955 62.925 ;
        RECT 92.245 62.755 94.245 62.925 ;
        RECT 94.535 62.755 96.535 62.925 ;
        RECT 96.825 62.755 98.825 62.925 ;
        RECT 99.115 62.755 101.115 62.925 ;
        RECT 101.405 62.755 103.405 62.925 ;
        RECT 103.695 62.755 105.695 62.925 ;
        RECT 105.985 62.755 107.985 62.925 ;
        RECT 108.715 62.235 108.885 72.085 ;
        RECT 109.615 71.395 111.615 71.565 ;
        RECT 111.905 71.395 113.905 71.565 ;
        RECT 114.195 71.395 116.195 71.565 ;
        RECT 116.485 71.395 118.485 71.565 ;
        RECT 118.775 71.395 120.775 71.565 ;
        RECT 121.065 71.395 123.065 71.565 ;
        RECT 123.355 71.395 125.355 71.565 ;
        RECT 125.645 71.395 127.645 71.565 ;
        RECT 109.385 63.140 109.555 71.180 ;
        RECT 111.675 63.140 111.845 71.180 ;
        RECT 113.965 63.140 114.135 71.180 ;
        RECT 116.255 63.140 116.425 71.180 ;
        RECT 118.545 63.140 118.715 71.180 ;
        RECT 120.835 63.140 121.005 71.180 ;
        RECT 123.125 63.140 123.295 71.180 ;
        RECT 125.415 63.140 125.585 71.180 ;
        RECT 127.705 63.140 127.875 71.180 ;
        RECT 109.615 62.755 111.615 62.925 ;
        RECT 111.905 62.755 113.905 62.925 ;
        RECT 114.195 62.755 116.195 62.925 ;
        RECT 116.485 62.755 118.485 62.925 ;
        RECT 118.775 62.755 120.775 62.925 ;
        RECT 121.065 62.755 123.065 62.925 ;
        RECT 123.355 62.755 125.355 62.925 ;
        RECT 125.645 62.755 127.645 62.925 ;
        RECT 128.375 62.235 128.905 72.085 ;
        RECT 10.055 62.065 128.905 62.235 ;
        RECT 10.055 52.215 10.585 62.065 ;
        RECT 11.315 61.375 13.315 61.545 ;
        RECT 13.605 61.375 15.605 61.545 ;
        RECT 15.895 61.375 17.895 61.545 ;
        RECT 18.185 61.375 20.185 61.545 ;
        RECT 20.475 61.375 22.475 61.545 ;
        RECT 22.765 61.375 24.765 61.545 ;
        RECT 25.055 61.375 27.055 61.545 ;
        RECT 27.345 61.375 29.345 61.545 ;
        RECT 11.085 53.120 11.255 61.160 ;
        RECT 13.375 53.120 13.545 61.160 ;
        RECT 15.665 53.120 15.835 61.160 ;
        RECT 17.955 53.120 18.125 61.160 ;
        RECT 20.245 53.120 20.415 61.160 ;
        RECT 22.535 53.120 22.705 61.160 ;
        RECT 24.825 53.120 24.995 61.160 ;
        RECT 27.115 53.120 27.285 61.160 ;
        RECT 29.405 53.120 29.575 61.160 ;
        RECT 11.315 52.735 13.315 52.905 ;
        RECT 13.605 52.735 15.605 52.905 ;
        RECT 15.895 52.735 17.895 52.905 ;
        RECT 18.185 52.735 20.185 52.905 ;
        RECT 20.475 52.735 22.475 52.905 ;
        RECT 22.765 52.735 24.765 52.905 ;
        RECT 25.055 52.735 27.055 52.905 ;
        RECT 27.345 52.735 29.345 52.905 ;
        RECT 30.075 52.215 30.245 62.065 ;
        RECT 30.975 61.375 32.975 61.545 ;
        RECT 33.265 61.375 35.265 61.545 ;
        RECT 35.555 61.375 37.555 61.545 ;
        RECT 37.845 61.375 39.845 61.545 ;
        RECT 40.135 61.375 42.135 61.545 ;
        RECT 42.425 61.375 44.425 61.545 ;
        RECT 44.715 61.375 46.715 61.545 ;
        RECT 47.005 61.375 49.005 61.545 ;
        RECT 30.745 53.120 30.915 61.160 ;
        RECT 33.035 53.120 33.205 61.160 ;
        RECT 35.325 53.120 35.495 61.160 ;
        RECT 37.615 53.120 37.785 61.160 ;
        RECT 39.905 53.120 40.075 61.160 ;
        RECT 42.195 53.120 42.365 61.160 ;
        RECT 44.485 53.120 44.655 61.160 ;
        RECT 46.775 53.120 46.945 61.160 ;
        RECT 49.065 53.120 49.235 61.160 ;
        RECT 30.975 52.735 32.975 52.905 ;
        RECT 33.265 52.735 35.265 52.905 ;
        RECT 35.555 52.735 37.555 52.905 ;
        RECT 37.845 52.735 39.845 52.905 ;
        RECT 40.135 52.735 42.135 52.905 ;
        RECT 42.425 52.735 44.425 52.905 ;
        RECT 44.715 52.735 46.715 52.905 ;
        RECT 47.005 52.735 49.005 52.905 ;
        RECT 49.735 52.215 49.905 62.065 ;
        RECT 50.635 61.375 52.635 61.545 ;
        RECT 52.925 61.375 54.925 61.545 ;
        RECT 55.215 61.375 57.215 61.545 ;
        RECT 57.505 61.375 59.505 61.545 ;
        RECT 59.795 61.375 61.795 61.545 ;
        RECT 62.085 61.375 64.085 61.545 ;
        RECT 64.375 61.375 66.375 61.545 ;
        RECT 66.665 61.375 68.665 61.545 ;
        RECT 50.405 53.120 50.575 61.160 ;
        RECT 52.695 53.120 52.865 61.160 ;
        RECT 54.985 53.120 55.155 61.160 ;
        RECT 57.275 53.120 57.445 61.160 ;
        RECT 59.565 53.120 59.735 61.160 ;
        RECT 61.855 53.120 62.025 61.160 ;
        RECT 64.145 53.120 64.315 61.160 ;
        RECT 66.435 53.120 66.605 61.160 ;
        RECT 68.725 53.120 68.895 61.160 ;
        RECT 50.635 52.735 52.635 52.905 ;
        RECT 52.925 52.735 54.925 52.905 ;
        RECT 55.215 52.735 57.215 52.905 ;
        RECT 57.505 52.735 59.505 52.905 ;
        RECT 59.795 52.735 61.795 52.905 ;
        RECT 62.085 52.735 64.085 52.905 ;
        RECT 64.375 52.735 66.375 52.905 ;
        RECT 66.665 52.735 68.665 52.905 ;
        RECT 69.395 52.215 69.565 62.065 ;
        RECT 70.295 61.375 72.295 61.545 ;
        RECT 72.585 61.375 74.585 61.545 ;
        RECT 74.875 61.375 76.875 61.545 ;
        RECT 77.165 61.375 79.165 61.545 ;
        RECT 79.455 61.375 81.455 61.545 ;
        RECT 81.745 61.375 83.745 61.545 ;
        RECT 84.035 61.375 86.035 61.545 ;
        RECT 86.325 61.375 88.325 61.545 ;
        RECT 70.065 53.120 70.235 61.160 ;
        RECT 72.355 53.120 72.525 61.160 ;
        RECT 74.645 53.120 74.815 61.160 ;
        RECT 76.935 53.120 77.105 61.160 ;
        RECT 79.225 53.120 79.395 61.160 ;
        RECT 81.515 53.120 81.685 61.160 ;
        RECT 83.805 53.120 83.975 61.160 ;
        RECT 86.095 53.120 86.265 61.160 ;
        RECT 88.385 53.120 88.555 61.160 ;
        RECT 70.295 52.735 72.295 52.905 ;
        RECT 72.585 52.735 74.585 52.905 ;
        RECT 74.875 52.735 76.875 52.905 ;
        RECT 77.165 52.735 79.165 52.905 ;
        RECT 79.455 52.735 81.455 52.905 ;
        RECT 81.745 52.735 83.745 52.905 ;
        RECT 84.035 52.735 86.035 52.905 ;
        RECT 86.325 52.735 88.325 52.905 ;
        RECT 89.055 52.215 89.225 62.065 ;
        RECT 89.955 61.375 91.955 61.545 ;
        RECT 92.245 61.375 94.245 61.545 ;
        RECT 94.535 61.375 96.535 61.545 ;
        RECT 96.825 61.375 98.825 61.545 ;
        RECT 99.115 61.375 101.115 61.545 ;
        RECT 101.405 61.375 103.405 61.545 ;
        RECT 103.695 61.375 105.695 61.545 ;
        RECT 105.985 61.375 107.985 61.545 ;
        RECT 89.725 53.120 89.895 61.160 ;
        RECT 92.015 53.120 92.185 61.160 ;
        RECT 94.305 53.120 94.475 61.160 ;
        RECT 96.595 53.120 96.765 61.160 ;
        RECT 98.885 53.120 99.055 61.160 ;
        RECT 101.175 53.120 101.345 61.160 ;
        RECT 103.465 53.120 103.635 61.160 ;
        RECT 105.755 53.120 105.925 61.160 ;
        RECT 108.045 53.120 108.215 61.160 ;
        RECT 89.955 52.735 91.955 52.905 ;
        RECT 92.245 52.735 94.245 52.905 ;
        RECT 94.535 52.735 96.535 52.905 ;
        RECT 96.825 52.735 98.825 52.905 ;
        RECT 99.115 52.735 101.115 52.905 ;
        RECT 101.405 52.735 103.405 52.905 ;
        RECT 103.695 52.735 105.695 52.905 ;
        RECT 105.985 52.735 107.985 52.905 ;
        RECT 108.715 52.215 108.885 62.065 ;
        RECT 109.615 61.375 111.615 61.545 ;
        RECT 111.905 61.375 113.905 61.545 ;
        RECT 114.195 61.375 116.195 61.545 ;
        RECT 116.485 61.375 118.485 61.545 ;
        RECT 118.775 61.375 120.775 61.545 ;
        RECT 121.065 61.375 123.065 61.545 ;
        RECT 123.355 61.375 125.355 61.545 ;
        RECT 125.645 61.375 127.645 61.545 ;
        RECT 109.385 53.120 109.555 61.160 ;
        RECT 111.675 53.120 111.845 61.160 ;
        RECT 113.965 53.120 114.135 61.160 ;
        RECT 116.255 53.120 116.425 61.160 ;
        RECT 118.545 53.120 118.715 61.160 ;
        RECT 120.835 53.120 121.005 61.160 ;
        RECT 123.125 53.120 123.295 61.160 ;
        RECT 125.415 53.120 125.585 61.160 ;
        RECT 127.705 53.120 127.875 61.160 ;
        RECT 109.615 52.735 111.615 52.905 ;
        RECT 111.905 52.735 113.905 52.905 ;
        RECT 114.195 52.735 116.195 52.905 ;
        RECT 116.485 52.735 118.485 52.905 ;
        RECT 118.775 52.735 120.775 52.905 ;
        RECT 121.065 52.735 123.065 52.905 ;
        RECT 123.355 52.735 125.355 52.905 ;
        RECT 125.645 52.735 127.645 52.905 ;
        RECT 128.375 52.215 128.905 62.065 ;
        RECT 10.055 52.045 128.905 52.215 ;
        RECT 10.055 42.195 10.585 52.045 ;
        RECT 11.315 51.355 13.315 51.525 ;
        RECT 13.605 51.355 15.605 51.525 ;
        RECT 15.895 51.355 17.895 51.525 ;
        RECT 18.185 51.355 20.185 51.525 ;
        RECT 20.475 51.355 22.475 51.525 ;
        RECT 22.765 51.355 24.765 51.525 ;
        RECT 25.055 51.355 27.055 51.525 ;
        RECT 27.345 51.355 29.345 51.525 ;
        RECT 11.085 43.100 11.255 51.140 ;
        RECT 13.375 43.100 13.545 51.140 ;
        RECT 15.665 43.100 15.835 51.140 ;
        RECT 17.955 43.100 18.125 51.140 ;
        RECT 20.245 43.100 20.415 51.140 ;
        RECT 22.535 43.100 22.705 51.140 ;
        RECT 24.825 43.100 24.995 51.140 ;
        RECT 27.115 43.100 27.285 51.140 ;
        RECT 29.405 43.100 29.575 51.140 ;
        RECT 11.315 42.715 13.315 42.885 ;
        RECT 13.605 42.715 15.605 42.885 ;
        RECT 15.895 42.715 17.895 42.885 ;
        RECT 18.185 42.715 20.185 42.885 ;
        RECT 20.475 42.715 22.475 42.885 ;
        RECT 22.765 42.715 24.765 42.885 ;
        RECT 25.055 42.715 27.055 42.885 ;
        RECT 27.345 42.715 29.345 42.885 ;
        RECT 30.075 42.195 30.245 52.045 ;
        RECT 30.975 51.355 32.975 51.525 ;
        RECT 33.265 51.355 35.265 51.525 ;
        RECT 35.555 51.355 37.555 51.525 ;
        RECT 37.845 51.355 39.845 51.525 ;
        RECT 40.135 51.355 42.135 51.525 ;
        RECT 42.425 51.355 44.425 51.525 ;
        RECT 44.715 51.355 46.715 51.525 ;
        RECT 47.005 51.355 49.005 51.525 ;
        RECT 30.745 43.100 30.915 51.140 ;
        RECT 33.035 43.100 33.205 51.140 ;
        RECT 35.325 43.100 35.495 51.140 ;
        RECT 37.615 43.100 37.785 51.140 ;
        RECT 39.905 43.100 40.075 51.140 ;
        RECT 42.195 43.100 42.365 51.140 ;
        RECT 44.485 43.100 44.655 51.140 ;
        RECT 46.775 43.100 46.945 51.140 ;
        RECT 49.065 43.100 49.235 51.140 ;
        RECT 30.975 42.715 32.975 42.885 ;
        RECT 33.265 42.715 35.265 42.885 ;
        RECT 35.555 42.715 37.555 42.885 ;
        RECT 37.845 42.715 39.845 42.885 ;
        RECT 40.135 42.715 42.135 42.885 ;
        RECT 42.425 42.715 44.425 42.885 ;
        RECT 44.715 42.715 46.715 42.885 ;
        RECT 47.005 42.715 49.005 42.885 ;
        RECT 49.735 42.195 49.905 52.045 ;
        RECT 50.635 51.355 52.635 51.525 ;
        RECT 52.925 51.355 54.925 51.525 ;
        RECT 55.215 51.355 57.215 51.525 ;
        RECT 57.505 51.355 59.505 51.525 ;
        RECT 59.795 51.355 61.795 51.525 ;
        RECT 62.085 51.355 64.085 51.525 ;
        RECT 64.375 51.355 66.375 51.525 ;
        RECT 66.665 51.355 68.665 51.525 ;
        RECT 50.405 43.100 50.575 51.140 ;
        RECT 52.695 43.100 52.865 51.140 ;
        RECT 54.985 43.100 55.155 51.140 ;
        RECT 57.275 43.100 57.445 51.140 ;
        RECT 59.565 43.100 59.735 51.140 ;
        RECT 61.855 43.100 62.025 51.140 ;
        RECT 64.145 43.100 64.315 51.140 ;
        RECT 66.435 43.100 66.605 51.140 ;
        RECT 68.725 43.100 68.895 51.140 ;
        RECT 50.635 42.715 52.635 42.885 ;
        RECT 52.925 42.715 54.925 42.885 ;
        RECT 55.215 42.715 57.215 42.885 ;
        RECT 57.505 42.715 59.505 42.885 ;
        RECT 59.795 42.715 61.795 42.885 ;
        RECT 62.085 42.715 64.085 42.885 ;
        RECT 64.375 42.715 66.375 42.885 ;
        RECT 66.665 42.715 68.665 42.885 ;
        RECT 69.395 42.195 69.565 52.045 ;
        RECT 70.295 51.355 72.295 51.525 ;
        RECT 72.585 51.355 74.585 51.525 ;
        RECT 74.875 51.355 76.875 51.525 ;
        RECT 77.165 51.355 79.165 51.525 ;
        RECT 79.455 51.355 81.455 51.525 ;
        RECT 81.745 51.355 83.745 51.525 ;
        RECT 84.035 51.355 86.035 51.525 ;
        RECT 86.325 51.355 88.325 51.525 ;
        RECT 70.065 43.100 70.235 51.140 ;
        RECT 72.355 43.100 72.525 51.140 ;
        RECT 74.645 43.100 74.815 51.140 ;
        RECT 76.935 43.100 77.105 51.140 ;
        RECT 79.225 43.100 79.395 51.140 ;
        RECT 81.515 43.100 81.685 51.140 ;
        RECT 83.805 43.100 83.975 51.140 ;
        RECT 86.095 43.100 86.265 51.140 ;
        RECT 88.385 43.100 88.555 51.140 ;
        RECT 70.295 42.715 72.295 42.885 ;
        RECT 72.585 42.715 74.585 42.885 ;
        RECT 74.875 42.715 76.875 42.885 ;
        RECT 77.165 42.715 79.165 42.885 ;
        RECT 79.455 42.715 81.455 42.885 ;
        RECT 81.745 42.715 83.745 42.885 ;
        RECT 84.035 42.715 86.035 42.885 ;
        RECT 86.325 42.715 88.325 42.885 ;
        RECT 89.055 42.195 89.225 52.045 ;
        RECT 89.955 51.355 91.955 51.525 ;
        RECT 92.245 51.355 94.245 51.525 ;
        RECT 94.535 51.355 96.535 51.525 ;
        RECT 96.825 51.355 98.825 51.525 ;
        RECT 99.115 51.355 101.115 51.525 ;
        RECT 101.405 51.355 103.405 51.525 ;
        RECT 103.695 51.355 105.695 51.525 ;
        RECT 105.985 51.355 107.985 51.525 ;
        RECT 89.725 43.100 89.895 51.140 ;
        RECT 92.015 43.100 92.185 51.140 ;
        RECT 94.305 43.100 94.475 51.140 ;
        RECT 96.595 43.100 96.765 51.140 ;
        RECT 98.885 43.100 99.055 51.140 ;
        RECT 101.175 43.100 101.345 51.140 ;
        RECT 103.465 43.100 103.635 51.140 ;
        RECT 105.755 43.100 105.925 51.140 ;
        RECT 108.045 43.100 108.215 51.140 ;
        RECT 89.955 42.715 91.955 42.885 ;
        RECT 92.245 42.715 94.245 42.885 ;
        RECT 94.535 42.715 96.535 42.885 ;
        RECT 96.825 42.715 98.825 42.885 ;
        RECT 99.115 42.715 101.115 42.885 ;
        RECT 101.405 42.715 103.405 42.885 ;
        RECT 103.695 42.715 105.695 42.885 ;
        RECT 105.985 42.715 107.985 42.885 ;
        RECT 108.715 42.195 108.885 52.045 ;
        RECT 109.615 51.355 111.615 51.525 ;
        RECT 111.905 51.355 113.905 51.525 ;
        RECT 114.195 51.355 116.195 51.525 ;
        RECT 116.485 51.355 118.485 51.525 ;
        RECT 118.775 51.355 120.775 51.525 ;
        RECT 121.065 51.355 123.065 51.525 ;
        RECT 123.355 51.355 125.355 51.525 ;
        RECT 125.645 51.355 127.645 51.525 ;
        RECT 109.385 43.100 109.555 51.140 ;
        RECT 111.675 43.100 111.845 51.140 ;
        RECT 113.965 43.100 114.135 51.140 ;
        RECT 116.255 43.100 116.425 51.140 ;
        RECT 118.545 43.100 118.715 51.140 ;
        RECT 120.835 43.100 121.005 51.140 ;
        RECT 123.125 43.100 123.295 51.140 ;
        RECT 125.415 43.100 125.585 51.140 ;
        RECT 127.705 43.100 127.875 51.140 ;
        RECT 109.615 42.715 111.615 42.885 ;
        RECT 111.905 42.715 113.905 42.885 ;
        RECT 114.195 42.715 116.195 42.885 ;
        RECT 116.485 42.715 118.485 42.885 ;
        RECT 118.775 42.715 120.775 42.885 ;
        RECT 121.065 42.715 123.065 42.885 ;
        RECT 123.355 42.715 125.355 42.885 ;
        RECT 125.645 42.715 127.645 42.885 ;
        RECT 128.375 42.195 128.905 52.045 ;
        RECT 10.055 41.665 128.905 42.195 ;
        RECT 10.055 39.070 74.665 39.600 ;
        RECT 10.055 29.310 10.585 39.070 ;
        RECT 11.375 38.380 13.375 38.550 ;
        RECT 13.665 38.380 15.665 38.550 ;
        RECT 15.955 38.380 17.955 38.550 ;
        RECT 18.245 38.380 20.245 38.550 ;
        RECT 11.145 30.170 11.315 38.210 ;
        RECT 13.435 30.170 13.605 38.210 ;
        RECT 15.725 30.170 15.895 38.210 ;
        RECT 18.015 30.170 18.185 38.210 ;
        RECT 20.305 30.170 20.475 38.210 ;
        RECT 11.375 29.830 13.375 30.000 ;
        RECT 13.665 29.830 15.665 30.000 ;
        RECT 15.955 29.830 17.955 30.000 ;
        RECT 18.245 29.830 20.245 30.000 ;
        RECT 21.035 29.310 21.205 39.070 ;
        RECT 21.995 38.380 23.995 38.550 ;
        RECT 24.285 38.380 26.285 38.550 ;
        RECT 26.575 38.380 28.575 38.550 ;
        RECT 28.865 38.380 30.865 38.550 ;
        RECT 21.765 30.170 21.935 38.210 ;
        RECT 24.055 30.170 24.225 38.210 ;
        RECT 26.345 30.170 26.515 38.210 ;
        RECT 28.635 30.170 28.805 38.210 ;
        RECT 30.925 30.170 31.095 38.210 ;
        RECT 21.995 29.830 23.995 30.000 ;
        RECT 24.285 29.830 26.285 30.000 ;
        RECT 26.575 29.830 28.575 30.000 ;
        RECT 28.865 29.830 30.865 30.000 ;
        RECT 31.655 29.310 31.825 39.070 ;
        RECT 32.615 38.380 34.615 38.550 ;
        RECT 34.905 38.380 36.905 38.550 ;
        RECT 37.195 38.380 39.195 38.550 ;
        RECT 39.485 38.380 41.485 38.550 ;
        RECT 32.385 30.170 32.555 38.210 ;
        RECT 34.675 30.170 34.845 38.210 ;
        RECT 36.965 30.170 37.135 38.210 ;
        RECT 39.255 30.170 39.425 38.210 ;
        RECT 41.545 30.170 41.715 38.210 ;
        RECT 32.615 29.830 34.615 30.000 ;
        RECT 34.905 29.830 36.905 30.000 ;
        RECT 37.195 29.830 39.195 30.000 ;
        RECT 39.485 29.830 41.485 30.000 ;
        RECT 42.275 29.310 42.445 39.070 ;
        RECT 43.235 38.380 45.235 38.550 ;
        RECT 45.525 38.380 47.525 38.550 ;
        RECT 47.815 38.380 49.815 38.550 ;
        RECT 50.105 38.380 52.105 38.550 ;
        RECT 43.005 30.170 43.175 38.210 ;
        RECT 45.295 30.170 45.465 38.210 ;
        RECT 47.585 30.170 47.755 38.210 ;
        RECT 49.875 30.170 50.045 38.210 ;
        RECT 52.165 30.170 52.335 38.210 ;
        RECT 43.235 29.830 45.235 30.000 ;
        RECT 45.525 29.830 47.525 30.000 ;
        RECT 47.815 29.830 49.815 30.000 ;
        RECT 50.105 29.830 52.105 30.000 ;
        RECT 52.895 29.310 53.065 39.070 ;
        RECT 53.855 38.380 55.855 38.550 ;
        RECT 56.145 38.380 58.145 38.550 ;
        RECT 58.435 38.380 60.435 38.550 ;
        RECT 60.725 38.380 62.725 38.550 ;
        RECT 53.625 30.170 53.795 38.210 ;
        RECT 55.915 30.170 56.085 38.210 ;
        RECT 58.205 30.170 58.375 38.210 ;
        RECT 60.495 30.170 60.665 38.210 ;
        RECT 62.785 30.170 62.955 38.210 ;
        RECT 53.855 29.830 55.855 30.000 ;
        RECT 56.145 29.830 58.145 30.000 ;
        RECT 58.435 29.830 60.435 30.000 ;
        RECT 60.725 29.830 62.725 30.000 ;
        RECT 63.515 29.310 63.685 39.070 ;
        RECT 64.475 38.380 66.475 38.550 ;
        RECT 66.765 38.380 68.765 38.550 ;
        RECT 69.055 38.380 71.055 38.550 ;
        RECT 71.345 38.380 73.345 38.550 ;
        RECT 64.245 30.170 64.415 38.210 ;
        RECT 66.535 30.170 66.705 38.210 ;
        RECT 68.825 30.170 68.995 38.210 ;
        RECT 71.115 30.170 71.285 38.210 ;
        RECT 73.405 30.170 73.575 38.210 ;
        RECT 64.475 29.830 66.475 30.000 ;
        RECT 66.765 29.830 68.765 30.000 ;
        RECT 69.055 29.830 71.055 30.000 ;
        RECT 71.345 29.830 73.345 30.000 ;
        RECT 74.135 29.310 74.665 39.070 ;
        RECT 10.055 29.140 74.665 29.310 ;
        RECT 10.055 19.380 10.585 29.140 ;
        RECT 11.375 28.450 13.375 28.620 ;
        RECT 13.665 28.450 15.665 28.620 ;
        RECT 15.955 28.450 17.955 28.620 ;
        RECT 18.245 28.450 20.245 28.620 ;
        RECT 11.145 20.240 11.315 28.280 ;
        RECT 13.435 20.240 13.605 28.280 ;
        RECT 15.725 20.240 15.895 28.280 ;
        RECT 18.015 20.240 18.185 28.280 ;
        RECT 20.305 20.240 20.475 28.280 ;
        RECT 11.375 19.900 13.375 20.070 ;
        RECT 13.665 19.900 15.665 20.070 ;
        RECT 15.955 19.900 17.955 20.070 ;
        RECT 18.245 19.900 20.245 20.070 ;
        RECT 21.035 19.380 21.205 29.140 ;
        RECT 21.995 28.450 23.995 28.620 ;
        RECT 24.285 28.450 26.285 28.620 ;
        RECT 26.575 28.450 28.575 28.620 ;
        RECT 28.865 28.450 30.865 28.620 ;
        RECT 21.765 20.240 21.935 28.280 ;
        RECT 24.055 20.240 24.225 28.280 ;
        RECT 26.345 20.240 26.515 28.280 ;
        RECT 28.635 20.240 28.805 28.280 ;
        RECT 30.925 20.240 31.095 28.280 ;
        RECT 21.995 19.900 23.995 20.070 ;
        RECT 24.285 19.900 26.285 20.070 ;
        RECT 26.575 19.900 28.575 20.070 ;
        RECT 28.865 19.900 30.865 20.070 ;
        RECT 31.655 19.380 31.825 29.140 ;
        RECT 32.615 28.450 34.615 28.620 ;
        RECT 34.905 28.450 36.905 28.620 ;
        RECT 37.195 28.450 39.195 28.620 ;
        RECT 39.485 28.450 41.485 28.620 ;
        RECT 32.385 20.240 32.555 28.280 ;
        RECT 34.675 20.240 34.845 28.280 ;
        RECT 36.965 20.240 37.135 28.280 ;
        RECT 39.255 20.240 39.425 28.280 ;
        RECT 41.545 20.240 41.715 28.280 ;
        RECT 32.615 19.900 34.615 20.070 ;
        RECT 34.905 19.900 36.905 20.070 ;
        RECT 37.195 19.900 39.195 20.070 ;
        RECT 39.485 19.900 41.485 20.070 ;
        RECT 42.275 19.380 42.445 29.140 ;
        RECT 43.235 28.450 45.235 28.620 ;
        RECT 45.525 28.450 47.525 28.620 ;
        RECT 47.815 28.450 49.815 28.620 ;
        RECT 50.105 28.450 52.105 28.620 ;
        RECT 43.005 20.240 43.175 28.280 ;
        RECT 45.295 20.240 45.465 28.280 ;
        RECT 47.585 20.240 47.755 28.280 ;
        RECT 49.875 20.240 50.045 28.280 ;
        RECT 52.165 20.240 52.335 28.280 ;
        RECT 43.235 19.900 45.235 20.070 ;
        RECT 45.525 19.900 47.525 20.070 ;
        RECT 47.815 19.900 49.815 20.070 ;
        RECT 50.105 19.900 52.105 20.070 ;
        RECT 52.895 19.380 53.065 29.140 ;
        RECT 53.855 28.450 55.855 28.620 ;
        RECT 56.145 28.450 58.145 28.620 ;
        RECT 58.435 28.450 60.435 28.620 ;
        RECT 60.725 28.450 62.725 28.620 ;
        RECT 53.625 20.240 53.795 28.280 ;
        RECT 55.915 20.240 56.085 28.280 ;
        RECT 58.205 20.240 58.375 28.280 ;
        RECT 60.495 20.240 60.665 28.280 ;
        RECT 62.785 20.240 62.955 28.280 ;
        RECT 53.855 19.900 55.855 20.070 ;
        RECT 56.145 19.900 58.145 20.070 ;
        RECT 58.435 19.900 60.435 20.070 ;
        RECT 60.725 19.900 62.725 20.070 ;
        RECT 63.515 19.380 63.685 29.140 ;
        RECT 64.475 28.450 66.475 28.620 ;
        RECT 66.765 28.450 68.765 28.620 ;
        RECT 69.055 28.450 71.055 28.620 ;
        RECT 71.345 28.450 73.345 28.620 ;
        RECT 64.245 20.240 64.415 28.280 ;
        RECT 66.535 20.240 66.705 28.280 ;
        RECT 68.825 20.240 68.995 28.280 ;
        RECT 71.115 20.240 71.285 28.280 ;
        RECT 73.405 20.240 73.575 28.280 ;
        RECT 64.475 19.900 66.475 20.070 ;
        RECT 66.765 19.900 68.765 20.070 ;
        RECT 69.055 19.900 71.055 20.070 ;
        RECT 71.345 19.900 73.345 20.070 ;
        RECT 74.135 19.380 74.665 29.140 ;
        RECT 10.055 19.210 74.665 19.380 ;
        RECT 10.055 9.450 10.585 19.210 ;
        RECT 11.375 18.520 13.375 18.690 ;
        RECT 13.665 18.520 15.665 18.690 ;
        RECT 15.955 18.520 17.955 18.690 ;
        RECT 18.245 18.520 20.245 18.690 ;
        RECT 11.145 10.310 11.315 18.350 ;
        RECT 13.435 10.310 13.605 18.350 ;
        RECT 15.725 10.310 15.895 18.350 ;
        RECT 18.015 10.310 18.185 18.350 ;
        RECT 20.305 10.310 20.475 18.350 ;
        RECT 11.375 9.970 13.375 10.140 ;
        RECT 13.665 9.970 15.665 10.140 ;
        RECT 15.955 9.970 17.955 10.140 ;
        RECT 18.245 9.970 20.245 10.140 ;
        RECT 21.035 9.450 21.205 19.210 ;
        RECT 21.995 18.520 23.995 18.690 ;
        RECT 24.285 18.520 26.285 18.690 ;
        RECT 26.575 18.520 28.575 18.690 ;
        RECT 28.865 18.520 30.865 18.690 ;
        RECT 21.765 10.310 21.935 18.350 ;
        RECT 24.055 10.310 24.225 18.350 ;
        RECT 26.345 10.310 26.515 18.350 ;
        RECT 28.635 10.310 28.805 18.350 ;
        RECT 30.925 10.310 31.095 18.350 ;
        RECT 21.995 9.970 23.995 10.140 ;
        RECT 24.285 9.970 26.285 10.140 ;
        RECT 26.575 9.970 28.575 10.140 ;
        RECT 28.865 9.970 30.865 10.140 ;
        RECT 31.655 9.450 31.825 19.210 ;
        RECT 32.615 18.520 34.615 18.690 ;
        RECT 34.905 18.520 36.905 18.690 ;
        RECT 37.195 18.520 39.195 18.690 ;
        RECT 39.485 18.520 41.485 18.690 ;
        RECT 32.385 10.310 32.555 18.350 ;
        RECT 34.675 10.310 34.845 18.350 ;
        RECT 36.965 10.310 37.135 18.350 ;
        RECT 39.255 10.310 39.425 18.350 ;
        RECT 41.545 10.310 41.715 18.350 ;
        RECT 32.615 9.970 34.615 10.140 ;
        RECT 34.905 9.970 36.905 10.140 ;
        RECT 37.195 9.970 39.195 10.140 ;
        RECT 39.485 9.970 41.485 10.140 ;
        RECT 42.275 9.450 42.445 19.210 ;
        RECT 43.235 18.520 45.235 18.690 ;
        RECT 45.525 18.520 47.525 18.690 ;
        RECT 47.815 18.520 49.815 18.690 ;
        RECT 50.105 18.520 52.105 18.690 ;
        RECT 43.005 10.310 43.175 18.350 ;
        RECT 45.295 10.310 45.465 18.350 ;
        RECT 47.585 10.310 47.755 18.350 ;
        RECT 49.875 10.310 50.045 18.350 ;
        RECT 52.165 10.310 52.335 18.350 ;
        RECT 43.235 9.970 45.235 10.140 ;
        RECT 45.525 9.970 47.525 10.140 ;
        RECT 47.815 9.970 49.815 10.140 ;
        RECT 50.105 9.970 52.105 10.140 ;
        RECT 52.895 9.450 53.065 19.210 ;
        RECT 53.855 18.520 55.855 18.690 ;
        RECT 56.145 18.520 58.145 18.690 ;
        RECT 58.435 18.520 60.435 18.690 ;
        RECT 60.725 18.520 62.725 18.690 ;
        RECT 53.625 10.310 53.795 18.350 ;
        RECT 55.915 10.310 56.085 18.350 ;
        RECT 58.205 10.310 58.375 18.350 ;
        RECT 60.495 10.310 60.665 18.350 ;
        RECT 62.785 10.310 62.955 18.350 ;
        RECT 53.855 9.970 55.855 10.140 ;
        RECT 56.145 9.970 58.145 10.140 ;
        RECT 58.435 9.970 60.435 10.140 ;
        RECT 60.725 9.970 62.725 10.140 ;
        RECT 63.515 9.450 63.685 19.210 ;
        RECT 64.475 18.520 66.475 18.690 ;
        RECT 66.765 18.520 68.765 18.690 ;
        RECT 69.055 18.520 71.055 18.690 ;
        RECT 71.345 18.520 73.345 18.690 ;
        RECT 64.245 10.310 64.415 18.350 ;
        RECT 66.535 10.310 66.705 18.350 ;
        RECT 68.825 10.310 68.995 18.350 ;
        RECT 71.115 10.310 71.285 18.350 ;
        RECT 73.405 10.310 73.575 18.350 ;
        RECT 64.475 9.970 66.475 10.140 ;
        RECT 66.765 9.970 68.765 10.140 ;
        RECT 69.055 9.970 71.055 10.140 ;
        RECT 71.345 9.970 73.345 10.140 ;
        RECT 74.135 9.450 74.665 19.210 ;
        RECT 10.055 8.920 74.665 9.450 ;
        RECT 79.695 39.070 128.905 39.600 ;
        RECT 79.695 29.310 80.225 39.070 ;
        RECT 80.785 38.210 85.535 39.070 ;
        RECT 80.785 30.170 80.955 38.210 ;
        RECT 83.075 30.170 83.245 38.210 ;
        RECT 85.365 30.170 85.535 38.210 ;
        RECT 81.015 29.830 83.015 30.000 ;
        RECT 83.305 29.830 85.305 30.000 ;
        RECT 86.095 29.310 86.265 39.070 ;
        RECT 87.055 38.380 89.055 38.550 ;
        RECT 89.345 38.380 91.345 38.550 ;
        RECT 86.825 30.170 86.995 38.210 ;
        RECT 89.115 30.170 89.285 38.210 ;
        RECT 91.405 30.170 91.575 38.210 ;
        RECT 87.055 29.830 89.055 30.000 ;
        RECT 89.345 29.830 91.345 30.000 ;
        RECT 92.135 29.310 92.305 39.070 ;
        RECT 93.095 38.380 95.095 38.550 ;
        RECT 95.385 38.380 97.385 38.550 ;
        RECT 92.865 30.170 93.035 38.210 ;
        RECT 95.155 30.170 95.325 38.210 ;
        RECT 97.445 30.170 97.615 38.210 ;
        RECT 93.095 29.830 95.095 30.000 ;
        RECT 95.385 29.830 97.385 30.000 ;
        RECT 98.175 29.310 98.345 39.070 ;
        RECT 99.135 38.380 101.135 38.550 ;
        RECT 101.425 38.380 103.425 38.550 ;
        RECT 98.905 30.170 99.075 38.210 ;
        RECT 101.195 30.170 101.365 38.210 ;
        RECT 103.485 30.170 103.655 38.210 ;
        RECT 99.135 29.830 101.135 30.000 ;
        RECT 101.425 29.830 103.425 30.000 ;
        RECT 104.215 29.310 104.385 39.070 ;
        RECT 105.175 38.380 107.175 38.550 ;
        RECT 107.465 38.380 109.465 38.550 ;
        RECT 104.945 30.170 105.115 38.210 ;
        RECT 107.235 30.170 107.405 38.210 ;
        RECT 109.525 30.170 109.695 38.210 ;
        RECT 105.175 29.830 107.175 30.000 ;
        RECT 107.465 29.830 109.465 30.000 ;
        RECT 110.255 29.310 110.425 39.070 ;
        RECT 111.215 38.380 113.215 38.550 ;
        RECT 113.505 38.380 115.505 38.550 ;
        RECT 110.985 30.170 111.155 38.210 ;
        RECT 113.275 30.170 113.445 38.210 ;
        RECT 115.565 30.170 115.735 38.210 ;
        RECT 111.215 29.830 113.215 30.000 ;
        RECT 113.505 29.830 115.505 30.000 ;
        RECT 116.295 29.310 116.465 39.070 ;
        RECT 117.255 38.380 119.255 38.550 ;
        RECT 119.545 38.380 121.545 38.550 ;
        RECT 117.025 30.170 117.195 38.210 ;
        RECT 119.315 30.170 119.485 38.210 ;
        RECT 121.605 30.170 121.775 38.210 ;
        RECT 117.255 29.830 119.255 30.000 ;
        RECT 119.545 29.830 121.545 30.000 ;
        RECT 122.335 29.310 122.505 39.070 ;
        RECT 123.065 38.210 127.815 39.070 ;
        RECT 123.065 30.170 123.235 38.210 ;
        RECT 125.355 30.170 125.525 38.210 ;
        RECT 127.645 30.170 127.815 38.210 ;
        RECT 123.295 29.830 125.295 30.000 ;
        RECT 125.585 29.830 127.585 30.000 ;
        RECT 128.375 29.310 128.905 39.070 ;
        RECT 79.695 29.140 128.905 29.310 ;
        RECT 79.695 19.380 80.225 29.140 ;
        RECT 81.015 28.450 83.015 28.620 ;
        RECT 83.305 28.450 85.305 28.620 ;
        RECT 80.785 20.240 80.955 28.280 ;
        RECT 83.075 20.240 83.245 28.280 ;
        RECT 85.365 20.240 85.535 28.280 ;
        RECT 80.785 19.380 85.535 20.240 ;
        RECT 86.095 19.380 86.265 29.140 ;
        RECT 87.055 28.450 89.055 28.620 ;
        RECT 89.345 28.450 91.345 28.620 ;
        RECT 86.825 20.240 86.995 28.280 ;
        RECT 89.115 20.240 89.285 28.280 ;
        RECT 91.405 20.240 91.575 28.280 ;
        RECT 87.055 19.900 89.055 20.070 ;
        RECT 89.345 19.900 91.345 20.070 ;
        RECT 92.135 19.380 92.305 29.140 ;
        RECT 93.095 28.450 95.095 28.620 ;
        RECT 95.385 28.450 97.385 28.620 ;
        RECT 92.865 20.240 93.035 28.280 ;
        RECT 95.155 20.240 95.325 28.280 ;
        RECT 97.445 20.240 97.615 28.280 ;
        RECT 93.095 19.900 95.095 20.070 ;
        RECT 95.385 19.900 97.385 20.070 ;
        RECT 98.175 19.380 98.345 29.140 ;
        RECT 99.135 28.450 101.135 28.620 ;
        RECT 101.425 28.450 103.425 28.620 ;
        RECT 98.905 20.240 99.075 28.280 ;
        RECT 101.195 20.240 101.365 28.280 ;
        RECT 103.485 20.240 103.655 28.280 ;
        RECT 99.135 19.900 101.135 20.070 ;
        RECT 101.425 19.900 103.425 20.070 ;
        RECT 104.215 19.380 104.385 29.140 ;
        RECT 105.175 28.450 107.175 28.620 ;
        RECT 107.465 28.450 109.465 28.620 ;
        RECT 104.945 20.240 105.115 28.280 ;
        RECT 107.235 20.240 107.405 28.280 ;
        RECT 109.525 20.240 109.695 28.280 ;
        RECT 105.175 19.900 107.175 20.070 ;
        RECT 107.465 19.900 109.465 20.070 ;
        RECT 110.255 19.380 110.425 29.140 ;
        RECT 111.215 28.450 113.215 28.620 ;
        RECT 113.505 28.450 115.505 28.620 ;
        RECT 110.985 20.240 111.155 28.280 ;
        RECT 113.275 20.240 113.445 28.280 ;
        RECT 115.565 20.240 115.735 28.280 ;
        RECT 111.215 19.900 113.215 20.070 ;
        RECT 113.505 19.900 115.505 20.070 ;
        RECT 116.295 19.380 116.465 29.140 ;
        RECT 117.255 28.450 119.255 28.620 ;
        RECT 119.545 28.450 121.545 28.620 ;
        RECT 117.025 20.240 117.195 28.280 ;
        RECT 119.315 20.240 119.485 28.280 ;
        RECT 121.605 20.240 121.775 28.280 ;
        RECT 117.255 19.900 119.255 20.070 ;
        RECT 119.545 19.900 121.545 20.070 ;
        RECT 122.335 19.380 122.505 29.140 ;
        RECT 123.295 28.450 125.295 28.620 ;
        RECT 125.585 28.450 127.585 28.620 ;
        RECT 123.065 20.240 123.235 28.280 ;
        RECT 125.355 20.240 125.525 28.280 ;
        RECT 127.645 20.240 127.815 28.280 ;
        RECT 123.065 19.380 127.815 20.240 ;
        RECT 128.375 19.380 128.905 29.140 ;
        RECT 79.695 19.210 128.905 19.380 ;
        RECT 79.695 9.450 80.225 19.210 ;
        RECT 81.015 18.520 83.015 18.690 ;
        RECT 83.305 18.520 85.305 18.690 ;
        RECT 80.785 10.310 80.955 18.350 ;
        RECT 83.075 10.310 83.245 18.350 ;
        RECT 85.365 10.310 85.535 18.350 ;
        RECT 80.785 9.450 85.535 10.310 ;
        RECT 86.095 9.450 86.265 19.210 ;
        RECT 87.055 18.520 89.055 18.690 ;
        RECT 89.345 18.520 91.345 18.690 ;
        RECT 86.825 10.310 86.995 18.350 ;
        RECT 89.115 10.310 89.285 18.350 ;
        RECT 91.405 10.310 91.575 18.350 ;
        RECT 86.825 9.450 91.575 10.310 ;
        RECT 92.135 9.450 92.305 19.210 ;
        RECT 93.095 18.520 95.095 18.690 ;
        RECT 95.385 18.520 97.385 18.690 ;
        RECT 92.865 10.310 93.035 18.350 ;
        RECT 95.155 10.310 95.325 18.350 ;
        RECT 97.445 10.310 97.615 18.350 ;
        RECT 92.865 9.450 97.615 10.310 ;
        RECT 98.175 9.450 98.345 19.210 ;
        RECT 99.135 18.520 101.135 18.690 ;
        RECT 101.425 18.520 103.425 18.690 ;
        RECT 98.905 10.310 99.075 18.350 ;
        RECT 101.195 10.310 101.365 18.350 ;
        RECT 103.485 10.310 103.655 18.350 ;
        RECT 98.905 9.450 103.655 10.310 ;
        RECT 104.215 9.450 104.385 19.210 ;
        RECT 105.175 18.520 107.175 18.690 ;
        RECT 107.465 18.520 109.465 18.690 ;
        RECT 104.945 10.310 105.115 18.350 ;
        RECT 107.235 10.310 107.405 18.350 ;
        RECT 109.525 10.310 109.695 18.350 ;
        RECT 104.945 9.450 109.695 10.310 ;
        RECT 110.255 9.450 110.425 19.210 ;
        RECT 111.215 18.520 113.215 18.690 ;
        RECT 113.505 18.520 115.505 18.690 ;
        RECT 110.985 10.310 111.155 18.350 ;
        RECT 113.275 10.310 113.445 18.350 ;
        RECT 115.565 10.310 115.735 18.350 ;
        RECT 110.985 9.450 115.735 10.310 ;
        RECT 116.295 9.450 116.465 19.210 ;
        RECT 117.255 18.520 119.255 18.690 ;
        RECT 119.545 18.520 121.545 18.690 ;
        RECT 117.025 10.310 117.195 18.350 ;
        RECT 119.315 10.310 119.485 18.350 ;
        RECT 121.605 10.310 121.775 18.350 ;
        RECT 117.025 9.450 121.775 10.310 ;
        RECT 122.335 9.450 122.505 19.210 ;
        RECT 123.295 18.520 125.295 18.690 ;
        RECT 125.585 18.520 127.585 18.690 ;
        RECT 123.065 10.310 123.235 18.350 ;
        RECT 125.355 10.310 125.525 18.350 ;
        RECT 127.645 10.310 127.815 18.350 ;
        RECT 123.065 9.450 127.815 10.310 ;
        RECT 128.375 9.450 128.905 19.210 ;
        RECT 135.150 18.895 135.680 104.785 ;
        RECT 136.265 103.615 138.425 104.305 ;
        RECT 136.265 102.445 138.425 103.135 ;
        RECT 136.265 101.275 138.425 101.965 ;
        RECT 136.265 100.105 138.425 100.795 ;
        RECT 136.265 98.935 138.425 99.625 ;
        RECT 136.265 97.765 138.425 98.455 ;
        RECT 136.265 96.595 138.425 97.285 ;
        RECT 136.265 95.425 138.425 96.115 ;
        RECT 136.265 94.255 138.425 94.945 ;
        RECT 136.265 93.085 138.425 93.775 ;
        RECT 136.265 91.915 138.425 92.605 ;
        RECT 136.265 90.745 138.425 91.435 ;
        RECT 136.265 89.575 138.425 90.265 ;
        RECT 136.265 88.405 138.425 89.095 ;
        RECT 136.265 87.235 138.425 87.925 ;
        RECT 136.265 86.065 138.425 86.755 ;
        RECT 136.265 84.895 138.425 85.585 ;
        RECT 136.265 83.725 138.425 84.415 ;
        RECT 136.265 82.555 138.425 83.245 ;
        RECT 136.265 81.385 138.425 82.075 ;
        RECT 136.265 80.215 138.425 80.905 ;
        RECT 136.265 79.045 138.425 79.735 ;
        RECT 136.265 77.875 138.425 78.565 ;
        RECT 136.265 76.705 138.425 77.395 ;
        RECT 136.265 75.535 138.425 76.225 ;
        RECT 136.265 74.365 138.425 75.055 ;
        RECT 136.265 73.195 138.425 73.885 ;
        RECT 136.265 72.025 138.425 72.715 ;
        RECT 136.265 70.855 138.425 71.545 ;
        RECT 136.265 69.685 138.425 70.375 ;
        RECT 136.265 68.515 138.425 69.205 ;
        RECT 136.265 67.345 138.425 68.035 ;
        RECT 136.265 66.175 138.425 66.865 ;
        RECT 136.265 65.005 138.425 65.695 ;
        RECT 136.265 63.835 138.425 64.525 ;
        RECT 136.265 62.665 138.425 63.355 ;
        RECT 136.265 61.495 138.425 62.185 ;
        RECT 136.265 60.325 138.425 61.015 ;
        RECT 136.265 59.155 138.425 59.845 ;
        RECT 136.265 57.985 138.425 58.675 ;
        RECT 136.265 56.815 138.425 57.505 ;
        RECT 136.265 55.645 138.425 56.335 ;
        RECT 136.265 54.475 138.425 55.165 ;
        RECT 136.265 53.305 138.425 53.995 ;
        RECT 136.265 52.135 138.425 52.825 ;
        RECT 136.265 50.965 138.425 51.655 ;
        RECT 136.265 49.795 138.425 50.485 ;
        RECT 136.265 48.625 138.425 49.315 ;
        RECT 136.265 47.455 138.425 48.145 ;
        RECT 136.265 46.285 138.425 46.975 ;
        RECT 136.265 45.115 138.425 45.805 ;
        RECT 136.265 43.945 138.425 44.635 ;
        RECT 136.265 42.775 138.425 43.465 ;
        RECT 136.265 41.605 138.425 42.295 ;
        RECT 136.265 40.435 138.425 41.125 ;
        RECT 136.265 39.265 138.425 39.955 ;
        RECT 136.265 38.095 138.425 38.785 ;
        RECT 136.265 36.925 138.425 37.615 ;
        RECT 136.265 35.755 138.425 36.445 ;
        RECT 136.265 34.585 138.425 35.275 ;
        RECT 136.265 33.415 138.425 34.105 ;
        RECT 136.265 32.245 138.425 32.935 ;
        RECT 136.265 31.075 138.425 31.765 ;
        RECT 136.265 29.905 138.425 30.595 ;
        RECT 136.265 28.735 138.425 29.425 ;
        RECT 136.265 27.565 138.425 28.255 ;
        RECT 136.265 26.395 138.425 27.085 ;
        RECT 136.265 25.225 138.425 25.915 ;
        RECT 136.265 24.055 138.425 24.745 ;
        RECT 136.265 22.885 138.425 23.575 ;
        RECT 136.265 21.715 138.425 22.405 ;
        RECT 136.265 20.545 138.425 21.235 ;
        RECT 136.265 19.375 138.425 20.065 ;
        RECT 139.150 18.895 145.540 104.785 ;
        RECT 146.265 103.615 148.425 104.305 ;
        RECT 146.265 102.445 148.425 103.135 ;
        RECT 146.265 101.275 148.425 101.965 ;
        RECT 146.265 100.105 148.425 100.795 ;
        RECT 146.265 98.935 148.425 99.625 ;
        RECT 146.265 97.765 148.425 98.455 ;
        RECT 146.265 96.595 148.425 97.285 ;
        RECT 146.265 95.425 148.425 96.115 ;
        RECT 146.265 94.255 148.425 94.945 ;
        RECT 146.265 93.085 148.425 93.775 ;
        RECT 146.265 91.915 148.425 92.605 ;
        RECT 146.265 90.745 148.425 91.435 ;
        RECT 146.265 89.575 148.425 90.265 ;
        RECT 146.265 88.405 148.425 89.095 ;
        RECT 146.265 87.235 148.425 87.925 ;
        RECT 146.265 86.065 148.425 86.755 ;
        RECT 146.265 84.895 148.425 85.585 ;
        RECT 146.265 83.725 148.425 84.415 ;
        RECT 146.265 82.555 148.425 83.245 ;
        RECT 146.265 81.385 148.425 82.075 ;
        RECT 146.265 80.215 148.425 80.905 ;
        RECT 146.265 79.045 148.425 79.735 ;
        RECT 146.265 77.875 148.425 78.565 ;
        RECT 146.265 76.705 148.425 77.395 ;
        RECT 146.265 75.535 148.425 76.225 ;
        RECT 146.265 74.365 148.425 75.055 ;
        RECT 146.265 73.195 148.425 73.885 ;
        RECT 146.265 72.025 148.425 72.715 ;
        RECT 146.265 70.855 148.425 71.545 ;
        RECT 146.265 69.685 148.425 70.375 ;
        RECT 146.265 68.515 148.425 69.205 ;
        RECT 146.265 67.345 148.425 68.035 ;
        RECT 146.265 66.175 148.425 66.865 ;
        RECT 146.265 65.005 148.425 65.695 ;
        RECT 146.265 63.835 148.425 64.525 ;
        RECT 146.265 62.665 148.425 63.355 ;
        RECT 146.265 61.495 148.425 62.185 ;
        RECT 146.265 60.325 148.425 61.015 ;
        RECT 146.265 59.155 148.425 59.845 ;
        RECT 146.265 57.985 148.425 58.675 ;
        RECT 146.265 56.815 148.425 57.505 ;
        RECT 146.265 55.645 148.425 56.335 ;
        RECT 146.265 54.475 148.425 55.165 ;
        RECT 146.265 53.305 148.425 53.995 ;
        RECT 146.265 52.135 148.425 52.825 ;
        RECT 146.265 50.965 148.425 51.655 ;
        RECT 146.265 49.795 148.425 50.485 ;
        RECT 146.265 48.625 148.425 49.315 ;
        RECT 146.265 47.455 148.425 48.145 ;
        RECT 146.265 46.285 148.425 46.975 ;
        RECT 146.265 45.115 148.425 45.805 ;
        RECT 146.265 43.945 148.425 44.635 ;
        RECT 146.265 42.775 148.425 43.465 ;
        RECT 146.265 41.605 148.425 42.295 ;
        RECT 146.265 40.435 148.425 41.125 ;
        RECT 146.265 39.265 148.425 39.955 ;
        RECT 146.265 38.095 148.425 38.785 ;
        RECT 146.265 36.925 148.425 37.615 ;
        RECT 146.265 35.755 148.425 36.445 ;
        RECT 146.265 34.585 148.425 35.275 ;
        RECT 146.265 33.415 148.425 34.105 ;
        RECT 146.265 32.245 148.425 32.935 ;
        RECT 146.265 31.075 148.425 31.765 ;
        RECT 146.265 29.905 148.425 30.595 ;
        RECT 146.265 28.735 148.425 29.425 ;
        RECT 146.265 27.565 148.425 28.255 ;
        RECT 146.265 26.395 148.425 27.085 ;
        RECT 146.265 25.225 148.425 25.915 ;
        RECT 146.265 24.055 148.425 24.745 ;
        RECT 146.265 22.885 148.425 23.575 ;
        RECT 146.265 21.715 148.425 22.405 ;
        RECT 146.265 20.545 148.425 21.235 ;
        RECT 146.265 19.375 148.425 20.065 ;
        RECT 149.010 18.895 149.540 104.785 ;
        RECT 135.150 13.490 149.540 18.895 ;
        RECT 79.695 8.920 128.905 9.450 ;
        RECT 155.300 4.700 155.700 180.620 ;
        RECT 4.300 4.300 155.700 4.700 ;
      LAYER met1 ;
        RECT 4.100 216.515 102.825 222.630 ;
        RECT 106.340 220.315 153.245 220.715 ;
        RECT 106.340 217.515 108.920 220.315 ;
        RECT 109.605 219.705 110.565 219.935 ;
        RECT 110.895 219.705 111.855 220.055 ;
        RECT 109.325 219.255 109.555 219.500 ;
        RECT 110.615 219.255 110.845 219.500 ;
        RECT 111.905 219.255 112.135 219.500 ;
        RECT 109.290 217.755 109.590 219.255 ;
        RECT 110.580 217.755 110.880 219.255 ;
        RECT 111.870 217.755 112.170 219.255 ;
        RECT 4.100 212.490 63.455 216.515 ;
        RECT 64.175 215.825 80.135 216.055 ;
        RECT 81.805 215.825 97.765 216.055 ;
        RECT 63.895 214.620 64.125 215.620 ;
        RECT 80.185 214.620 81.755 215.620 ;
        RECT 97.815 214.620 98.045 215.620 ;
        RECT 64.175 214.185 80.135 214.415 ;
        RECT 81.805 214.185 97.765 214.415 ;
        RECT 77.595 213.035 78.595 213.270 ;
        RECT 83.345 213.035 84.345 213.270 ;
        RECT 64.175 212.805 80.135 213.035 ;
        RECT 81.805 212.805 97.765 213.035 ;
        RECT 4.100 211.660 56.570 212.490 ;
        RECT 4.100 191.850 9.525 211.660 ;
        RECT 10.245 210.970 18.205 211.200 ;
        RECT 18.535 210.970 26.495 211.200 ;
        RECT 28.165 210.970 36.125 211.200 ;
        RECT 36.455 210.970 44.415 211.200 ;
        RECT 9.965 210.465 10.195 210.765 ;
        RECT 9.925 209.065 10.225 210.465 ;
        RECT 9.965 202.765 10.195 209.065 ;
        RECT 18.255 207.465 18.485 210.765 ;
        RECT 18.215 206.065 18.515 207.465 ;
        RECT 18.255 202.765 18.485 206.065 ;
        RECT 26.545 204.465 26.775 210.765 ;
        RECT 27.885 204.465 28.115 210.765 ;
        RECT 36.175 207.465 36.405 210.765 ;
        RECT 44.465 210.465 44.695 210.765 ;
        RECT 44.425 209.065 44.725 210.465 ;
        RECT 45.135 210.150 56.570 211.660 ;
        RECT 36.165 206.065 36.465 207.465 ;
        RECT 26.505 203.065 26.805 204.465 ;
        RECT 27.845 203.065 28.145 204.465 ;
        RECT 26.505 202.560 28.145 203.065 ;
        RECT 36.175 202.765 36.405 206.065 ;
        RECT 44.465 202.765 44.695 209.065 ;
        RECT 45.135 207.460 50.745 210.150 ;
        RECT 54.835 209.565 56.570 210.150 ;
        RECT 51.315 207.460 51.905 209.565 ;
        RECT 52.485 207.460 54.245 209.565 ;
        RECT 54.825 207.460 56.570 209.565 ;
        RECT 10.245 202.330 18.205 202.560 ;
        RECT 18.535 202.330 36.125 202.560 ;
        RECT 36.455 202.330 44.415 202.560 ;
        RECT 10.245 201.180 44.415 202.330 ;
        RECT 10.245 200.950 18.205 201.180 ;
        RECT 18.535 200.950 36.125 201.180 ;
        RECT 36.455 200.950 44.415 201.180 ;
        RECT 9.965 194.445 10.195 200.745 ;
        RECT 18.255 197.445 18.485 200.745 ;
        RECT 26.505 200.445 28.145 200.950 ;
        RECT 26.505 199.045 26.805 200.445 ;
        RECT 27.845 199.045 28.145 200.445 ;
        RECT 18.215 196.045 18.515 197.445 ;
        RECT 9.925 193.045 10.225 194.445 ;
        RECT 9.965 192.745 10.195 193.045 ;
        RECT 18.255 192.745 18.485 196.045 ;
        RECT 26.545 192.745 26.775 199.045 ;
        RECT 27.885 192.745 28.115 199.045 ;
        RECT 36.175 197.445 36.405 200.745 ;
        RECT 36.165 196.045 36.465 197.445 ;
        RECT 36.175 192.745 36.405 196.045 ;
        RECT 44.465 194.445 44.695 200.745 ;
        RECT 44.425 193.045 44.725 194.445 ;
        RECT 44.465 192.745 44.695 193.045 ;
        RECT 10.245 192.310 18.205 192.540 ;
        RECT 18.535 192.310 26.495 192.540 ;
        RECT 28.165 192.310 36.125 192.540 ;
        RECT 36.455 192.310 44.415 192.540 ;
        RECT 45.135 191.850 49.450 207.460 ;
        RECT 4.100 190.670 49.450 191.850 ;
        RECT 4.100 180.880 9.525 190.670 ;
        RECT 9.965 189.980 12.205 190.210 ;
        RECT 12.535 189.980 14.495 190.210 ;
        RECT 9.965 184.050 10.195 189.980 ;
        RECT 12.535 189.775 13.090 189.980 ;
        RECT 12.255 189.350 13.090 189.775 ;
        RECT 9.930 182.650 10.230 184.050 ;
        RECT 9.965 181.570 10.195 182.650 ;
        RECT 12.255 181.775 12.485 189.350 ;
        RECT 14.545 188.900 14.775 189.775 ;
        RECT 14.510 187.500 14.810 188.900 ;
        RECT 14.545 181.775 14.775 187.500 ;
        RECT 9.965 181.340 12.205 181.570 ;
        RECT 12.535 181.340 14.495 181.570 ;
        RECT 15.215 180.880 16.545 190.670 ;
        RECT 45.135 190.570 49.450 190.670 ;
        RECT 56.110 190.570 56.570 207.460 ;
        RECT 17.265 189.980 19.225 190.210 ;
        RECT 19.555 189.980 21.515 190.210 ;
        RECT 21.845 189.980 23.805 190.210 ;
        RECT 24.135 189.980 26.095 190.210 ;
        RECT 26.425 189.980 28.385 190.210 ;
        RECT 28.715 189.980 30.675 190.210 ;
        RECT 31.005 189.980 32.965 190.210 ;
        RECT 33.295 189.980 35.255 190.210 ;
        RECT 35.585 189.980 37.545 190.210 ;
        RECT 37.875 189.980 39.835 190.210 ;
        RECT 40.165 189.980 42.125 190.210 ;
        RECT 42.455 189.980 44.415 190.210 ;
        RECT 16.985 189.645 17.215 189.775 ;
        RECT 16.950 188.245 17.250 189.645 ;
        RECT 16.985 181.775 17.215 188.245 ;
        RECT 19.275 186.555 19.505 189.775 ;
        RECT 21.565 189.645 21.795 189.775 ;
        RECT 21.530 188.245 21.830 189.645 ;
        RECT 19.240 184.995 19.540 186.555 ;
        RECT 19.275 181.775 19.505 184.995 ;
        RECT 21.565 181.775 21.795 188.245 ;
        RECT 23.855 186.555 24.085 189.775 ;
        RECT 26.145 189.645 26.375 189.775 ;
        RECT 26.110 188.245 26.410 189.645 ;
        RECT 23.820 184.995 24.120 186.555 ;
        RECT 23.855 181.775 24.085 184.995 ;
        RECT 26.145 181.775 26.375 188.245 ;
        RECT 28.435 186.555 28.665 189.775 ;
        RECT 30.725 189.645 30.955 189.775 ;
        RECT 30.690 188.245 30.990 189.645 ;
        RECT 28.400 184.995 28.700 186.555 ;
        RECT 28.435 181.775 28.665 184.995 ;
        RECT 30.725 181.775 30.955 188.245 ;
        RECT 33.015 186.555 33.245 189.775 ;
        RECT 35.305 189.645 35.535 189.775 ;
        RECT 35.270 188.245 35.570 189.645 ;
        RECT 32.980 184.995 33.280 186.555 ;
        RECT 33.015 181.775 33.245 184.995 ;
        RECT 35.305 181.775 35.535 188.245 ;
        RECT 37.595 186.555 37.825 189.775 ;
        RECT 39.885 189.645 40.115 189.775 ;
        RECT 39.850 188.245 40.150 189.645 ;
        RECT 37.560 184.995 37.860 186.555 ;
        RECT 37.595 181.775 37.825 184.995 ;
        RECT 39.885 181.775 40.115 188.245 ;
        RECT 42.175 186.555 42.405 189.775 ;
        RECT 44.465 189.645 44.695 189.775 ;
        RECT 44.430 188.245 44.730 189.645 ;
        RECT 42.140 184.995 42.440 186.555 ;
        RECT 42.175 181.775 42.405 184.995 ;
        RECT 44.465 181.775 44.695 188.245 ;
        RECT 45.135 187.880 50.745 190.570 ;
        RECT 51.315 188.465 53.075 190.570 ;
        RECT 53.655 188.465 54.245 190.570 ;
        RECT 54.825 188.465 56.570 190.570 ;
        RECT 54.835 187.880 56.570 188.465 ;
        RECT 45.135 187.650 56.570 187.880 ;
        RECT 17.465 181.570 19.025 181.605 ;
        RECT 19.755 181.570 21.315 181.605 ;
        RECT 22.045 181.570 23.605 181.605 ;
        RECT 24.335 181.570 25.895 181.605 ;
        RECT 26.625 181.570 28.185 181.605 ;
        RECT 28.915 181.570 30.475 181.605 ;
        RECT 31.205 181.570 32.765 181.605 ;
        RECT 33.495 181.570 35.055 181.605 ;
        RECT 35.785 181.570 37.345 181.605 ;
        RECT 38.075 181.570 39.635 181.605 ;
        RECT 40.365 181.570 41.925 181.605 ;
        RECT 42.655 181.570 44.215 181.605 ;
        RECT 17.265 181.340 44.415 181.570 ;
        RECT 17.465 181.305 19.025 181.340 ;
        RECT 19.755 181.305 21.315 181.340 ;
        RECT 22.045 181.305 23.605 181.340 ;
        RECT 24.335 181.305 25.895 181.340 ;
        RECT 26.625 181.305 28.185 181.340 ;
        RECT 28.915 181.305 30.475 181.340 ;
        RECT 31.205 181.305 32.765 181.340 ;
        RECT 33.495 181.305 35.055 181.340 ;
        RECT 35.785 181.305 37.345 181.340 ;
        RECT 38.075 181.305 39.635 181.340 ;
        RECT 40.365 181.305 41.925 181.340 ;
        RECT 42.655 181.305 44.215 181.340 ;
        RECT 45.135 180.880 46.085 187.650 ;
        RECT 4.100 180.050 46.085 180.880 ;
        RECT 4.100 127.485 4.900 180.050 ;
        RECT 5.910 178.420 53.180 179.250 ;
        RECT 5.910 168.720 9.530 178.420 ;
        RECT 17.400 177.960 18.800 178.130 ;
        RECT 19.690 177.960 21.090 178.130 ;
        RECT 26.560 177.960 27.960 178.130 ;
        RECT 28.850 177.960 30.250 178.130 ;
        RECT 35.720 177.960 37.120 178.130 ;
        RECT 38.010 177.960 39.410 178.130 ;
        RECT 44.880 177.960 46.280 178.130 ;
        RECT 47.170 177.960 48.570 178.130 ;
        RECT 49.460 177.960 50.860 178.130 ;
        RECT 10.250 177.730 12.210 177.960 ;
        RECT 12.540 177.730 14.500 177.960 ;
        RECT 14.830 177.730 16.790 177.960 ;
        RECT 17.120 177.730 19.080 177.960 ;
        RECT 19.410 177.730 21.370 177.960 ;
        RECT 21.700 177.730 23.660 177.960 ;
        RECT 23.990 177.730 25.950 177.960 ;
        RECT 26.280 177.730 28.240 177.960 ;
        RECT 28.570 177.730 30.530 177.960 ;
        RECT 30.860 177.730 32.820 177.960 ;
        RECT 33.150 177.730 35.110 177.960 ;
        RECT 35.440 177.730 37.400 177.960 ;
        RECT 37.730 177.730 39.690 177.960 ;
        RECT 40.020 177.730 41.980 177.960 ;
        RECT 42.310 177.730 44.270 177.960 ;
        RECT 44.600 177.730 46.560 177.960 ;
        RECT 46.890 177.730 48.850 177.960 ;
        RECT 49.180 177.730 51.140 177.960 ;
        RECT 9.970 174.270 10.200 177.570 ;
        RECT 12.260 174.270 12.490 177.570 ;
        RECT 14.550 176.670 14.780 177.570 ;
        RECT 14.465 175.270 14.865 176.670 ;
        RECT 9.885 172.870 10.285 174.270 ;
        RECT 12.175 172.870 12.575 174.270 ;
        RECT 9.970 169.570 10.200 172.870 ;
        RECT 12.260 169.570 12.490 172.870 ;
        RECT 14.550 169.570 14.780 175.270 ;
        RECT 16.840 174.270 17.070 177.570 ;
        RECT 16.755 172.870 17.155 174.270 ;
        RECT 16.840 169.570 17.070 172.870 ;
        RECT 19.130 171.870 19.360 177.570 ;
        RECT 21.420 174.270 21.650 177.570 ;
        RECT 23.710 176.670 23.940 177.570 ;
        RECT 23.625 175.270 24.025 176.670 ;
        RECT 21.335 172.870 21.735 174.270 ;
        RECT 19.045 170.470 19.445 171.870 ;
        RECT 19.130 169.570 19.360 170.470 ;
        RECT 21.420 169.570 21.650 172.870 ;
        RECT 23.710 169.570 23.940 175.270 ;
        RECT 26.000 174.270 26.230 177.570 ;
        RECT 25.915 172.870 26.315 174.270 ;
        RECT 26.000 169.570 26.230 172.870 ;
        RECT 28.290 171.870 28.520 177.570 ;
        RECT 30.580 174.270 30.810 177.570 ;
        RECT 32.870 176.670 33.100 177.570 ;
        RECT 32.785 175.270 33.185 176.670 ;
        RECT 30.495 172.870 30.895 174.270 ;
        RECT 28.205 170.470 28.605 171.870 ;
        RECT 28.290 169.570 28.520 170.470 ;
        RECT 30.580 169.570 30.810 172.870 ;
        RECT 32.870 169.570 33.100 175.270 ;
        RECT 35.160 174.270 35.390 177.570 ;
        RECT 35.075 172.870 35.475 174.270 ;
        RECT 35.160 169.570 35.390 172.870 ;
        RECT 37.450 171.870 37.680 177.570 ;
        RECT 39.740 174.270 39.970 177.570 ;
        RECT 42.030 176.670 42.260 177.570 ;
        RECT 41.945 175.270 42.345 176.670 ;
        RECT 39.655 172.870 40.055 174.270 ;
        RECT 37.365 170.470 37.765 171.870 ;
        RECT 37.450 169.570 37.680 170.470 ;
        RECT 39.740 169.570 39.970 172.870 ;
        RECT 42.030 169.570 42.260 175.270 ;
        RECT 44.320 174.270 44.550 177.570 ;
        RECT 44.235 172.870 44.635 174.270 ;
        RECT 44.320 169.570 44.550 172.870 ;
        RECT 46.610 171.870 46.840 177.570 ;
        RECT 48.900 174.270 49.130 177.570 ;
        RECT 51.190 174.270 51.420 177.570 ;
        RECT 48.815 172.870 49.215 174.270 ;
        RECT 51.105 172.870 51.505 174.270 ;
        RECT 46.525 170.470 46.925 171.870 ;
        RECT 46.610 169.570 46.840 170.470 ;
        RECT 48.900 169.570 49.130 172.870 ;
        RECT 51.190 169.570 51.420 172.870 ;
        RECT 10.250 169.180 12.210 169.410 ;
        RECT 12.540 169.180 14.500 169.410 ;
        RECT 14.830 169.180 16.790 169.410 ;
        RECT 17.120 169.180 19.080 169.410 ;
        RECT 19.410 169.180 21.370 169.410 ;
        RECT 21.700 169.180 23.660 169.410 ;
        RECT 23.990 169.180 25.950 169.410 ;
        RECT 26.280 169.180 28.240 169.410 ;
        RECT 28.570 169.180 30.530 169.410 ;
        RECT 30.860 169.180 32.820 169.410 ;
        RECT 33.150 169.180 35.110 169.410 ;
        RECT 35.440 169.180 37.400 169.410 ;
        RECT 37.730 169.180 39.690 169.410 ;
        RECT 40.020 169.180 41.980 169.410 ;
        RECT 42.310 169.180 44.270 169.410 ;
        RECT 44.600 169.180 46.560 169.410 ;
        RECT 46.890 169.180 48.850 169.410 ;
        RECT 49.180 169.180 51.140 169.410 ;
        RECT 10.530 169.010 11.930 169.180 ;
        RECT 12.820 169.010 14.220 169.180 ;
        RECT 15.110 169.010 16.510 169.180 ;
        RECT 21.980 169.010 23.380 169.180 ;
        RECT 24.270 169.010 25.670 169.180 ;
        RECT 31.140 169.010 32.540 169.180 ;
        RECT 33.430 169.010 34.830 169.180 ;
        RECT 40.300 169.010 41.700 169.180 ;
        RECT 42.590 169.010 43.990 169.180 ;
        RECT 51.860 168.720 53.180 178.420 ;
        RECT 5.910 167.830 53.180 168.720 ;
        RECT 5.910 148.290 9.530 167.830 ;
        RECT 10.310 167.140 12.270 167.370 ;
        RECT 12.600 167.140 14.560 167.370 ;
        RECT 16.350 167.140 18.310 167.370 ;
        RECT 18.640 167.140 20.600 167.370 ;
        RECT 22.390 167.140 24.350 167.370 ;
        RECT 24.680 167.140 26.640 167.370 ;
        RECT 28.430 167.140 30.390 167.370 ;
        RECT 30.720 167.140 32.680 167.370 ;
        RECT 34.470 167.140 36.430 167.370 ;
        RECT 36.760 167.140 38.720 167.370 ;
        RECT 40.510 167.140 42.470 167.370 ;
        RECT 42.800 167.140 44.760 167.370 ;
        RECT 46.550 167.140 48.510 167.370 ;
        RECT 48.840 167.140 50.800 167.370 ;
        RECT 10.030 161.265 10.260 166.980 ;
        RECT 12.320 161.265 12.550 166.980 ;
        RECT 14.610 161.265 14.840 166.980 ;
        RECT 16.070 161.265 16.300 166.980 ;
        RECT 18.360 166.565 18.590 166.980 ;
        RECT 18.325 165.865 18.625 166.565 ;
        RECT 9.995 159.865 10.295 161.265 ;
        RECT 12.285 159.865 12.585 161.265 ;
        RECT 14.575 159.865 14.875 161.265 ;
        RECT 16.035 159.865 16.335 161.265 ;
        RECT 10.030 158.820 10.260 159.865 ;
        RECT 12.320 158.820 12.550 159.865 ;
        RECT 14.610 158.820 14.840 159.865 ;
        RECT 16.070 158.980 16.300 159.865 ;
        RECT 18.360 158.980 18.590 165.865 ;
        RECT 20.650 161.265 20.880 166.980 ;
        RECT 22.110 161.265 22.340 166.980 ;
        RECT 24.400 166.565 24.630 166.980 ;
        RECT 24.365 165.865 24.665 166.565 ;
        RECT 20.615 159.865 20.915 161.265 ;
        RECT 22.075 159.865 22.375 161.265 ;
        RECT 20.650 158.980 20.880 159.865 ;
        RECT 22.110 158.980 22.340 159.865 ;
        RECT 24.400 158.980 24.630 165.865 ;
        RECT 26.690 161.265 26.920 166.980 ;
        RECT 28.150 161.265 28.380 166.980 ;
        RECT 30.440 162.965 30.670 166.980 ;
        RECT 30.405 162.265 30.705 162.965 ;
        RECT 26.655 159.865 26.955 161.265 ;
        RECT 28.115 159.865 28.415 161.265 ;
        RECT 26.690 158.980 26.920 159.865 ;
        RECT 28.150 158.980 28.380 159.865 ;
        RECT 30.440 158.980 30.670 162.265 ;
        RECT 32.730 161.265 32.960 166.980 ;
        RECT 34.190 161.265 34.420 166.980 ;
        RECT 36.480 166.565 36.710 166.980 ;
        RECT 36.445 165.865 36.745 166.565 ;
        RECT 32.695 159.865 32.995 161.265 ;
        RECT 34.155 159.865 34.455 161.265 ;
        RECT 32.730 158.980 32.960 159.865 ;
        RECT 34.190 158.980 34.420 159.865 ;
        RECT 36.480 158.980 36.710 165.865 ;
        RECT 38.770 161.265 39.000 166.980 ;
        RECT 40.230 161.265 40.460 166.980 ;
        RECT 42.520 166.565 42.750 166.980 ;
        RECT 42.485 165.865 42.785 166.565 ;
        RECT 38.735 159.865 39.035 161.265 ;
        RECT 40.195 159.865 40.495 161.265 ;
        RECT 38.770 158.980 39.000 159.865 ;
        RECT 40.230 158.980 40.460 159.865 ;
        RECT 42.520 158.980 42.750 165.865 ;
        RECT 44.810 161.265 45.040 166.980 ;
        RECT 46.270 161.265 46.500 166.980 ;
        RECT 48.560 161.265 48.790 166.980 ;
        RECT 50.850 161.265 51.080 166.980 ;
        RECT 44.775 159.865 45.075 161.265 ;
        RECT 46.235 159.865 46.535 161.265 ;
        RECT 48.525 159.865 48.825 161.265 ;
        RECT 50.815 159.865 51.115 161.265 ;
        RECT 44.810 158.980 45.040 159.865 ;
        RECT 46.270 158.820 46.500 159.865 ;
        RECT 48.560 158.820 48.790 159.865 ;
        RECT 50.850 158.820 51.080 159.865 ;
        RECT 10.030 158.590 14.840 158.820 ;
        RECT 10.030 157.210 14.840 157.440 ;
        RECT 16.350 157.210 44.760 158.820 ;
        RECT 46.270 158.590 51.080 158.820 ;
        RECT 46.270 157.210 51.080 157.440 ;
        RECT 10.030 156.165 10.260 157.210 ;
        RECT 12.320 156.165 12.550 157.210 ;
        RECT 14.610 156.165 14.840 157.210 ;
        RECT 16.070 156.165 16.300 157.050 ;
        RECT 9.995 154.765 10.295 156.165 ;
        RECT 12.285 154.765 12.585 156.165 ;
        RECT 14.575 154.765 14.875 156.165 ;
        RECT 16.035 154.765 16.335 156.165 ;
        RECT 10.030 149.050 10.260 154.765 ;
        RECT 12.320 149.050 12.550 154.765 ;
        RECT 14.610 149.050 14.840 154.765 ;
        RECT 16.070 149.050 16.300 154.765 ;
        RECT 18.360 150.165 18.590 157.050 ;
        RECT 20.650 156.165 20.880 157.050 ;
        RECT 22.110 156.165 22.340 157.050 ;
        RECT 20.615 154.765 20.915 156.165 ;
        RECT 22.075 154.765 22.375 156.165 ;
        RECT 18.325 149.465 18.625 150.165 ;
        RECT 18.360 149.050 18.590 149.465 ;
        RECT 20.650 149.050 20.880 154.765 ;
        RECT 22.110 149.050 22.340 154.765 ;
        RECT 24.400 151.965 24.630 157.050 ;
        RECT 26.690 156.165 26.920 157.050 ;
        RECT 28.150 156.165 28.380 157.050 ;
        RECT 26.655 154.765 26.955 156.165 ;
        RECT 28.115 154.765 28.415 156.165 ;
        RECT 24.365 151.265 24.665 151.965 ;
        RECT 24.400 149.050 24.630 151.265 ;
        RECT 26.690 149.050 26.920 154.765 ;
        RECT 28.150 149.050 28.380 154.765 ;
        RECT 30.440 149.050 30.670 157.210 ;
        RECT 32.730 156.165 32.960 157.050 ;
        RECT 32.695 154.765 32.995 156.165 ;
        RECT 32.730 149.050 32.960 154.765 ;
        RECT 34.190 149.050 34.420 157.210 ;
        RECT 36.480 149.050 36.710 157.210 ;
        RECT 38.770 149.050 39.000 157.210 ;
        RECT 40.230 156.165 40.460 157.050 ;
        RECT 40.195 154.765 40.495 156.165 ;
        RECT 40.230 149.050 40.460 154.765 ;
        RECT 42.520 150.165 42.750 157.050 ;
        RECT 44.810 156.165 45.040 157.050 ;
        RECT 46.270 156.165 46.500 157.210 ;
        RECT 48.560 156.165 48.790 157.210 ;
        RECT 50.850 156.165 51.080 157.210 ;
        RECT 44.775 154.765 45.075 156.165 ;
        RECT 46.235 154.765 46.535 156.165 ;
        RECT 48.525 154.765 48.825 156.165 ;
        RECT 50.815 154.765 51.115 156.165 ;
        RECT 42.485 149.465 42.785 150.165 ;
        RECT 42.520 149.050 42.750 149.465 ;
        RECT 44.810 149.050 45.040 154.765 ;
        RECT 46.270 149.050 46.500 154.765 ;
        RECT 48.560 149.050 48.790 154.765 ;
        RECT 50.850 149.050 51.080 154.765 ;
        RECT 10.310 148.660 12.270 148.890 ;
        RECT 12.600 148.660 14.560 148.890 ;
        RECT 16.350 148.660 18.310 148.890 ;
        RECT 18.640 148.660 20.600 148.890 ;
        RECT 22.390 148.660 24.350 148.890 ;
        RECT 24.680 148.660 26.640 148.890 ;
        RECT 28.430 148.660 30.390 148.890 ;
        RECT 30.720 148.660 32.680 148.890 ;
        RECT 34.470 148.660 36.430 148.890 ;
        RECT 36.760 148.660 38.720 148.890 ;
        RECT 40.510 148.660 42.470 148.890 ;
        RECT 42.800 148.660 44.760 148.890 ;
        RECT 46.550 148.660 48.510 148.890 ;
        RECT 48.840 148.660 50.800 148.890 ;
        RECT 51.580 148.290 53.180 167.830 ;
        RECT 5.910 143.745 53.180 148.290 ;
        RECT 62.865 171.445 63.455 212.490 ;
        RECT 63.895 211.600 64.595 212.600 ;
        RECT 77.595 212.570 78.595 212.805 ;
        RECT 77.595 211.395 78.595 211.630 ;
        RECT 80.185 211.600 81.755 212.600 ;
        RECT 83.345 212.570 84.345 212.805 ;
        RECT 83.345 211.395 84.345 211.630 ;
        RECT 97.345 211.600 98.045 212.600 ;
        RECT 64.175 211.165 80.135 211.395 ;
        RECT 81.805 211.165 97.765 211.395 ;
        RECT 77.595 210.930 78.595 211.165 ;
        RECT 83.345 210.930 84.345 211.165 ;
        RECT 77.595 210.015 78.595 210.250 ;
        RECT 83.345 210.015 84.345 210.250 ;
        RECT 64.175 209.785 80.135 210.015 ;
        RECT 81.805 209.785 97.765 210.015 ;
        RECT 63.895 208.580 64.595 209.580 ;
        RECT 77.595 209.550 78.595 209.785 ;
        RECT 77.595 208.375 78.595 208.610 ;
        RECT 80.185 208.580 81.755 209.580 ;
        RECT 83.345 209.550 84.345 209.785 ;
        RECT 83.345 208.375 84.345 208.610 ;
        RECT 97.345 208.580 98.045 209.580 ;
        RECT 64.175 208.145 80.135 208.375 ;
        RECT 81.805 208.145 97.765 208.375 ;
        RECT 77.595 207.910 78.595 208.145 ;
        RECT 83.345 207.910 84.345 208.145 ;
        RECT 77.595 206.995 78.595 207.230 ;
        RECT 83.345 206.995 84.345 207.230 ;
        RECT 64.175 206.765 80.135 206.995 ;
        RECT 81.805 206.765 97.765 206.995 ;
        RECT 63.895 205.560 64.595 206.560 ;
        RECT 77.595 206.530 78.595 206.765 ;
        RECT 77.595 205.355 78.595 205.590 ;
        RECT 80.185 205.560 81.755 206.560 ;
        RECT 83.345 206.530 84.345 206.765 ;
        RECT 83.345 205.355 84.345 205.590 ;
        RECT 97.345 205.560 98.045 206.560 ;
        RECT 64.175 205.125 80.135 205.355 ;
        RECT 81.805 205.125 97.765 205.355 ;
        RECT 77.595 204.890 78.595 205.125 ;
        RECT 83.345 204.890 84.345 205.125 ;
        RECT 77.595 203.975 78.595 204.210 ;
        RECT 83.345 203.975 84.345 204.210 ;
        RECT 64.175 203.745 80.135 203.975 ;
        RECT 81.805 203.745 97.765 203.975 ;
        RECT 63.895 202.540 75.695 203.540 ;
        RECT 77.595 203.510 78.595 203.745 ;
        RECT 77.595 202.335 78.595 202.570 ;
        RECT 80.185 202.540 81.755 203.540 ;
        RECT 83.345 203.510 84.345 203.745 ;
        RECT 83.345 202.335 84.345 202.570 ;
        RECT 86.245 202.540 98.045 203.540 ;
        RECT 64.175 202.105 80.135 202.335 ;
        RECT 81.805 202.105 97.765 202.335 ;
        RECT 77.595 201.870 78.595 202.105 ;
        RECT 83.345 201.870 84.345 202.105 ;
        RECT 77.595 200.955 78.595 201.190 ;
        RECT 83.345 200.955 84.345 201.190 ;
        RECT 64.175 200.725 80.135 200.955 ;
        RECT 81.805 200.725 97.765 200.955 ;
        RECT 63.895 199.520 70.195 200.520 ;
        RECT 77.595 200.490 78.595 200.725 ;
        RECT 77.595 199.315 78.595 199.550 ;
        RECT 80.185 199.520 81.755 200.520 ;
        RECT 83.345 200.490 84.345 200.725 ;
        RECT 83.345 199.315 84.345 199.550 ;
        RECT 91.745 199.520 98.045 200.520 ;
        RECT 64.175 199.085 80.135 199.315 ;
        RECT 81.805 199.085 97.765 199.315 ;
        RECT 77.595 198.850 78.595 199.085 ;
        RECT 83.345 198.850 84.345 199.085 ;
        RECT 77.595 197.935 78.595 198.170 ;
        RECT 83.345 197.935 84.345 198.170 ;
        RECT 64.175 197.705 80.135 197.935 ;
        RECT 81.805 197.705 97.765 197.935 ;
        RECT 63.895 196.500 67.445 197.500 ;
        RECT 77.595 197.470 78.595 197.705 ;
        RECT 77.595 196.295 78.595 196.530 ;
        RECT 80.185 196.500 81.755 197.500 ;
        RECT 83.345 197.470 84.345 197.705 ;
        RECT 83.345 196.295 84.345 196.530 ;
        RECT 94.495 196.500 98.045 197.500 ;
        RECT 64.175 196.065 80.135 196.295 ;
        RECT 81.805 196.065 97.765 196.295 ;
        RECT 77.595 195.830 78.595 196.065 ;
        RECT 83.345 195.830 84.345 196.065 ;
        RECT 77.595 194.915 78.595 195.150 ;
        RECT 83.345 194.915 84.345 195.150 ;
        RECT 64.175 194.685 80.135 194.915 ;
        RECT 81.805 194.685 97.765 194.915 ;
        RECT 63.895 193.480 72.945 194.480 ;
        RECT 77.595 194.450 78.595 194.685 ;
        RECT 77.595 193.275 78.595 193.510 ;
        RECT 80.185 193.480 81.755 194.480 ;
        RECT 83.345 194.450 84.345 194.685 ;
        RECT 83.345 193.275 84.345 193.510 ;
        RECT 88.995 193.480 98.045 194.480 ;
        RECT 64.175 193.045 80.135 193.275 ;
        RECT 81.805 193.045 97.765 193.275 ;
        RECT 77.595 192.810 78.595 193.045 ;
        RECT 83.345 192.810 84.345 193.045 ;
        RECT 77.595 191.895 78.595 192.130 ;
        RECT 83.345 191.895 84.345 192.130 ;
        RECT 64.175 191.665 80.135 191.895 ;
        RECT 81.805 191.665 97.765 191.895 ;
        RECT 63.895 190.460 67.445 191.460 ;
        RECT 77.595 191.430 78.595 191.665 ;
        RECT 77.595 190.255 78.595 190.490 ;
        RECT 80.185 190.460 81.755 191.460 ;
        RECT 83.345 191.430 84.345 191.665 ;
        RECT 83.345 190.255 84.345 190.490 ;
        RECT 94.495 190.460 98.045 191.460 ;
        RECT 64.175 190.025 80.135 190.255 ;
        RECT 81.805 190.025 97.765 190.255 ;
        RECT 77.595 189.790 78.595 190.025 ;
        RECT 83.345 189.790 84.345 190.025 ;
        RECT 77.595 188.875 78.595 189.110 ;
        RECT 83.345 188.875 84.345 189.110 ;
        RECT 64.175 188.645 80.135 188.875 ;
        RECT 81.805 188.645 97.765 188.875 ;
        RECT 63.895 187.440 70.195 188.440 ;
        RECT 77.595 188.410 78.595 188.645 ;
        RECT 77.595 187.235 78.595 187.470 ;
        RECT 80.185 187.440 81.755 188.440 ;
        RECT 83.345 188.410 84.345 188.645 ;
        RECT 83.345 187.235 84.345 187.470 ;
        RECT 91.745 187.440 98.045 188.440 ;
        RECT 64.175 187.005 80.135 187.235 ;
        RECT 81.805 187.005 97.765 187.235 ;
        RECT 77.595 186.770 78.595 187.005 ;
        RECT 83.345 186.770 84.345 187.005 ;
        RECT 77.595 185.855 78.595 186.090 ;
        RECT 83.345 185.855 84.345 186.090 ;
        RECT 64.175 185.625 80.135 185.855 ;
        RECT 81.805 185.625 97.765 185.855 ;
        RECT 63.895 184.420 75.695 185.420 ;
        RECT 77.595 185.390 78.595 185.625 ;
        RECT 77.595 184.215 78.595 184.450 ;
        RECT 80.185 184.420 81.755 185.420 ;
        RECT 83.345 185.390 84.345 185.625 ;
        RECT 83.345 184.215 84.345 184.450 ;
        RECT 86.245 184.420 98.045 185.420 ;
        RECT 64.175 183.985 80.135 184.215 ;
        RECT 81.805 183.985 97.765 184.215 ;
        RECT 77.595 183.750 78.595 183.985 ;
        RECT 83.345 183.750 84.345 183.985 ;
        RECT 77.595 182.835 78.595 183.070 ;
        RECT 83.345 182.835 84.345 183.070 ;
        RECT 64.175 182.605 80.135 182.835 ;
        RECT 81.805 182.605 97.765 182.835 ;
        RECT 98.485 182.710 102.825 216.515 ;
        RECT 108.520 216.690 108.920 217.515 ;
        RECT 109.325 217.500 109.555 217.755 ;
        RECT 110.615 217.500 110.845 217.755 ;
        RECT 111.905 217.500 112.135 217.755 ;
        RECT 109.605 216.945 110.565 217.295 ;
        RECT 110.895 217.065 111.855 217.295 ;
        RECT 112.545 216.690 112.950 220.315 ;
        RECT 113.635 219.705 114.595 219.935 ;
        RECT 114.925 219.705 115.885 220.055 ;
        RECT 113.355 219.255 113.585 219.500 ;
        RECT 114.645 219.255 114.875 219.500 ;
        RECT 115.935 219.255 116.165 219.500 ;
        RECT 113.320 217.755 113.620 219.255 ;
        RECT 114.610 217.755 114.910 219.255 ;
        RECT 115.900 217.755 116.200 219.255 ;
        RECT 113.355 217.500 113.585 217.755 ;
        RECT 114.645 217.500 114.875 217.755 ;
        RECT 115.935 217.500 116.165 217.755 ;
        RECT 113.635 216.945 114.595 217.295 ;
        RECT 114.925 217.065 115.885 217.295 ;
        RECT 116.575 216.690 116.980 220.315 ;
        RECT 117.665 219.705 118.625 219.935 ;
        RECT 118.955 219.705 119.915 220.055 ;
        RECT 117.385 219.255 117.615 219.500 ;
        RECT 118.675 219.255 118.905 219.500 ;
        RECT 119.965 219.255 120.195 219.500 ;
        RECT 117.350 217.755 117.650 219.255 ;
        RECT 118.640 217.755 118.940 219.255 ;
        RECT 119.930 217.755 120.230 219.255 ;
        RECT 117.385 217.500 117.615 217.755 ;
        RECT 118.675 217.500 118.905 217.755 ;
        RECT 119.965 217.500 120.195 217.755 ;
        RECT 117.665 216.945 118.625 217.295 ;
        RECT 118.955 217.065 119.915 217.295 ;
        RECT 120.605 216.690 121.010 220.315 ;
        RECT 121.695 219.705 122.655 219.935 ;
        RECT 122.985 219.705 123.945 220.055 ;
        RECT 121.415 219.255 121.645 219.500 ;
        RECT 122.705 219.255 122.935 219.500 ;
        RECT 123.995 219.255 124.225 219.500 ;
        RECT 121.380 217.755 121.680 219.255 ;
        RECT 122.670 217.755 122.970 219.255 ;
        RECT 123.960 217.755 124.260 219.255 ;
        RECT 121.415 217.500 121.645 217.755 ;
        RECT 122.705 217.500 122.935 217.755 ;
        RECT 123.995 217.500 124.225 217.755 ;
        RECT 121.695 216.945 122.655 217.295 ;
        RECT 122.985 217.065 123.945 217.295 ;
        RECT 124.635 216.690 125.040 220.315 ;
        RECT 125.725 219.705 126.685 219.935 ;
        RECT 127.015 219.705 127.975 220.055 ;
        RECT 125.445 219.255 125.675 219.500 ;
        RECT 126.735 219.255 126.965 219.500 ;
        RECT 128.025 219.255 128.255 219.500 ;
        RECT 125.410 217.755 125.710 219.255 ;
        RECT 126.700 217.755 127.000 219.255 ;
        RECT 127.990 217.755 128.290 219.255 ;
        RECT 125.445 217.500 125.675 217.755 ;
        RECT 126.735 217.500 126.965 217.755 ;
        RECT 128.025 217.500 128.255 217.755 ;
        RECT 125.725 216.945 126.685 217.295 ;
        RECT 127.015 217.065 127.975 217.295 ;
        RECT 128.665 216.690 129.070 220.315 ;
        RECT 129.755 219.705 130.715 219.935 ;
        RECT 131.045 219.705 132.005 220.055 ;
        RECT 129.475 219.255 129.705 219.500 ;
        RECT 130.765 219.255 130.995 219.500 ;
        RECT 132.055 219.255 132.285 219.500 ;
        RECT 129.440 217.755 129.740 219.255 ;
        RECT 130.730 217.755 131.030 219.255 ;
        RECT 132.020 217.755 132.320 219.255 ;
        RECT 129.475 217.500 129.705 217.755 ;
        RECT 130.765 217.500 130.995 217.755 ;
        RECT 132.055 217.500 132.285 217.755 ;
        RECT 129.755 216.945 130.715 217.295 ;
        RECT 131.045 217.065 132.005 217.295 ;
        RECT 132.695 216.690 133.100 220.315 ;
        RECT 133.785 219.705 134.745 219.935 ;
        RECT 135.075 219.705 136.035 220.055 ;
        RECT 133.505 219.255 133.735 219.500 ;
        RECT 134.795 219.255 135.025 219.500 ;
        RECT 136.085 219.255 136.315 219.500 ;
        RECT 133.470 217.755 133.770 219.255 ;
        RECT 134.760 217.755 135.060 219.255 ;
        RECT 136.050 217.755 136.350 219.255 ;
        RECT 133.505 217.500 133.735 217.755 ;
        RECT 134.795 217.500 135.025 217.755 ;
        RECT 136.085 217.500 136.315 217.755 ;
        RECT 133.785 216.945 134.745 217.295 ;
        RECT 135.075 217.065 136.035 217.295 ;
        RECT 136.725 216.690 137.130 220.315 ;
        RECT 137.815 219.705 138.775 219.935 ;
        RECT 139.105 219.705 140.065 220.055 ;
        RECT 137.535 219.255 137.765 219.500 ;
        RECT 138.825 219.255 139.055 219.500 ;
        RECT 140.115 219.255 140.345 219.500 ;
        RECT 137.500 217.755 137.800 219.255 ;
        RECT 138.790 217.755 139.090 219.255 ;
        RECT 140.080 217.755 140.380 219.255 ;
        RECT 137.535 217.500 137.765 217.755 ;
        RECT 138.825 217.500 139.055 217.755 ;
        RECT 140.115 217.500 140.345 217.755 ;
        RECT 137.815 216.945 138.775 217.295 ;
        RECT 139.105 217.065 140.065 217.295 ;
        RECT 140.755 216.690 141.160 220.315 ;
        RECT 141.845 219.705 142.805 219.935 ;
        RECT 143.135 219.705 144.095 220.055 ;
        RECT 141.565 219.255 141.795 219.500 ;
        RECT 142.855 219.255 143.085 219.500 ;
        RECT 144.145 219.255 144.375 219.500 ;
        RECT 141.530 217.755 141.830 219.255 ;
        RECT 142.820 217.755 143.120 219.255 ;
        RECT 144.110 217.755 144.410 219.255 ;
        RECT 141.565 217.500 141.795 217.755 ;
        RECT 142.855 217.500 143.085 217.755 ;
        RECT 144.145 217.500 144.375 217.755 ;
        RECT 141.845 216.945 142.805 217.295 ;
        RECT 143.135 217.065 144.095 217.295 ;
        RECT 144.785 216.690 145.190 220.315 ;
        RECT 145.875 219.705 146.835 219.935 ;
        RECT 147.165 219.705 148.125 220.055 ;
        RECT 145.595 219.255 145.825 219.500 ;
        RECT 146.885 219.255 147.115 219.500 ;
        RECT 148.175 219.255 148.405 219.500 ;
        RECT 145.560 217.755 145.860 219.255 ;
        RECT 146.850 217.755 147.150 219.255 ;
        RECT 148.140 217.755 148.440 219.255 ;
        RECT 145.595 217.500 145.825 217.755 ;
        RECT 146.885 217.500 147.115 217.755 ;
        RECT 148.175 217.500 148.405 217.755 ;
        RECT 145.875 216.945 146.835 217.295 ;
        RECT 147.165 217.065 148.125 217.295 ;
        RECT 148.815 216.690 149.220 220.315 ;
        RECT 149.905 219.705 150.865 219.935 ;
        RECT 151.195 219.705 152.155 220.055 ;
        RECT 149.625 219.255 149.855 219.500 ;
        RECT 150.915 219.255 151.145 219.500 ;
        RECT 152.205 219.255 152.435 219.500 ;
        RECT 149.590 217.755 149.890 219.255 ;
        RECT 150.880 217.755 151.180 219.255 ;
        RECT 152.170 217.755 152.470 219.255 ;
        RECT 149.625 217.500 149.855 217.755 ;
        RECT 150.915 217.500 151.145 217.755 ;
        RECT 152.205 217.500 152.435 217.755 ;
        RECT 149.905 216.945 150.865 217.295 ;
        RECT 151.195 217.065 152.155 217.295 ;
        RECT 152.845 216.690 153.245 220.315 ;
        RECT 108.520 216.290 153.245 216.690 ;
        RECT 106.415 213.340 153.245 213.740 ;
        RECT 106.415 210.540 108.915 213.340 ;
        RECT 109.605 212.735 110.565 212.965 ;
        RECT 110.895 212.735 111.855 212.965 ;
        RECT 108.515 203.720 108.915 210.540 ;
        RECT 109.325 205.495 109.555 212.530 ;
        RECT 110.615 211.190 110.845 212.530 ;
        RECT 110.580 209.690 110.880 211.190 ;
        RECT 109.290 204.795 109.590 205.495 ;
        RECT 109.325 204.530 109.555 204.795 ;
        RECT 110.615 204.530 110.845 209.690 ;
        RECT 111.905 206.705 112.135 212.530 ;
        RECT 111.870 206.005 112.170 206.705 ;
        RECT 111.905 204.530 112.135 206.005 ;
        RECT 109.605 203.995 110.565 204.325 ;
        RECT 110.895 203.995 111.855 204.325 ;
        RECT 112.545 203.720 112.945 213.340 ;
        RECT 113.635 212.735 114.595 212.965 ;
        RECT 114.925 212.735 115.885 212.965 ;
        RECT 113.355 205.495 113.585 212.530 ;
        RECT 114.645 211.190 114.875 212.530 ;
        RECT 114.610 209.690 114.910 211.190 ;
        RECT 113.320 204.795 113.620 205.495 ;
        RECT 113.355 204.530 113.585 204.795 ;
        RECT 114.645 204.530 114.875 209.690 ;
        RECT 115.935 206.705 116.165 212.530 ;
        RECT 115.900 206.005 116.200 206.705 ;
        RECT 115.935 204.530 116.165 206.005 ;
        RECT 113.635 203.995 114.595 204.325 ;
        RECT 114.925 203.995 115.885 204.325 ;
        RECT 116.575 203.720 116.975 213.340 ;
        RECT 117.665 212.735 118.625 212.965 ;
        RECT 118.955 212.735 119.915 212.965 ;
        RECT 117.385 205.495 117.615 212.530 ;
        RECT 118.675 211.190 118.905 212.530 ;
        RECT 118.640 209.690 118.940 211.190 ;
        RECT 117.350 204.795 117.650 205.495 ;
        RECT 117.385 204.530 117.615 204.795 ;
        RECT 118.675 204.530 118.905 209.690 ;
        RECT 119.965 206.705 120.195 212.530 ;
        RECT 119.930 206.005 120.230 206.705 ;
        RECT 119.965 204.530 120.195 206.005 ;
        RECT 117.665 203.995 118.625 204.325 ;
        RECT 118.955 203.995 119.915 204.325 ;
        RECT 120.605 203.720 121.005 213.340 ;
        RECT 121.695 212.735 122.655 212.965 ;
        RECT 122.985 212.735 123.945 212.965 ;
        RECT 121.415 205.495 121.645 212.530 ;
        RECT 122.705 211.190 122.935 212.530 ;
        RECT 122.670 209.690 122.970 211.190 ;
        RECT 121.380 204.795 121.680 205.495 ;
        RECT 121.415 204.530 121.645 204.795 ;
        RECT 122.705 204.530 122.935 209.690 ;
        RECT 123.995 206.705 124.225 212.530 ;
        RECT 123.960 206.005 124.260 206.705 ;
        RECT 123.995 204.530 124.225 206.005 ;
        RECT 121.695 203.995 122.655 204.325 ;
        RECT 122.985 203.995 123.945 204.325 ;
        RECT 124.635 203.720 125.035 213.340 ;
        RECT 125.725 212.735 126.685 212.965 ;
        RECT 127.015 212.735 127.975 212.965 ;
        RECT 125.445 205.495 125.675 212.530 ;
        RECT 126.735 211.190 126.965 212.530 ;
        RECT 126.700 209.690 127.000 211.190 ;
        RECT 125.410 204.795 125.710 205.495 ;
        RECT 125.445 204.530 125.675 204.795 ;
        RECT 126.735 204.530 126.965 209.690 ;
        RECT 128.025 206.705 128.255 212.530 ;
        RECT 127.990 206.005 128.290 206.705 ;
        RECT 128.025 204.530 128.255 206.005 ;
        RECT 125.725 203.995 126.685 204.325 ;
        RECT 127.015 203.995 127.975 204.325 ;
        RECT 128.665 203.720 129.065 213.340 ;
        RECT 129.755 212.735 130.715 212.965 ;
        RECT 131.045 212.735 132.005 212.965 ;
        RECT 129.475 205.495 129.705 212.530 ;
        RECT 130.765 211.190 130.995 212.530 ;
        RECT 130.730 209.690 131.030 211.190 ;
        RECT 129.440 204.795 129.740 205.495 ;
        RECT 129.475 204.530 129.705 204.795 ;
        RECT 130.765 204.530 130.995 209.690 ;
        RECT 132.055 206.705 132.285 212.530 ;
        RECT 132.020 206.005 132.320 206.705 ;
        RECT 132.055 204.530 132.285 206.005 ;
        RECT 129.755 203.995 130.715 204.325 ;
        RECT 131.045 203.995 132.005 204.325 ;
        RECT 132.695 203.720 133.095 213.340 ;
        RECT 133.785 212.735 134.745 212.965 ;
        RECT 135.075 212.735 136.035 212.965 ;
        RECT 133.505 205.495 133.735 212.530 ;
        RECT 134.795 211.190 135.025 212.530 ;
        RECT 134.760 209.690 135.060 211.190 ;
        RECT 133.470 204.795 133.770 205.495 ;
        RECT 133.505 204.530 133.735 204.795 ;
        RECT 134.795 204.530 135.025 209.690 ;
        RECT 136.085 206.705 136.315 212.530 ;
        RECT 136.050 206.005 136.350 206.705 ;
        RECT 136.085 204.530 136.315 206.005 ;
        RECT 133.785 203.995 134.745 204.325 ;
        RECT 135.075 203.995 136.035 204.325 ;
        RECT 136.725 203.720 137.125 213.340 ;
        RECT 137.815 212.735 138.775 212.965 ;
        RECT 139.105 212.735 140.065 212.965 ;
        RECT 137.535 205.495 137.765 212.530 ;
        RECT 138.825 211.190 139.055 212.530 ;
        RECT 138.790 209.690 139.090 211.190 ;
        RECT 137.500 204.795 137.800 205.495 ;
        RECT 137.535 204.530 137.765 204.795 ;
        RECT 138.825 204.530 139.055 209.690 ;
        RECT 140.115 206.705 140.345 212.530 ;
        RECT 140.080 206.005 140.380 206.705 ;
        RECT 140.115 204.530 140.345 206.005 ;
        RECT 137.815 203.995 138.775 204.325 ;
        RECT 139.105 203.995 140.065 204.325 ;
        RECT 140.755 203.720 141.155 213.340 ;
        RECT 141.845 212.735 142.805 212.965 ;
        RECT 143.135 212.735 144.095 212.965 ;
        RECT 141.565 205.495 141.795 212.530 ;
        RECT 142.855 211.190 143.085 212.530 ;
        RECT 142.820 209.690 143.120 211.190 ;
        RECT 141.530 204.795 141.830 205.495 ;
        RECT 141.565 204.530 141.795 204.795 ;
        RECT 142.855 204.530 143.085 209.690 ;
        RECT 144.145 206.705 144.375 212.530 ;
        RECT 144.110 206.005 144.410 206.705 ;
        RECT 144.145 204.530 144.375 206.005 ;
        RECT 141.845 203.995 142.805 204.325 ;
        RECT 143.135 203.995 144.095 204.325 ;
        RECT 144.785 203.720 145.185 213.340 ;
        RECT 145.875 212.735 146.835 212.965 ;
        RECT 147.165 212.735 148.125 212.965 ;
        RECT 145.595 205.495 145.825 212.530 ;
        RECT 146.885 211.190 147.115 212.530 ;
        RECT 146.850 209.690 147.150 211.190 ;
        RECT 145.560 204.795 145.860 205.495 ;
        RECT 145.595 204.530 145.825 204.795 ;
        RECT 146.885 204.530 147.115 209.690 ;
        RECT 148.175 206.705 148.405 212.530 ;
        RECT 148.140 206.005 148.440 206.705 ;
        RECT 148.175 204.530 148.405 206.005 ;
        RECT 145.875 203.995 146.835 204.325 ;
        RECT 147.165 203.995 148.125 204.325 ;
        RECT 148.815 203.720 149.215 213.340 ;
        RECT 149.905 212.735 150.865 212.965 ;
        RECT 151.195 212.735 152.155 212.965 ;
        RECT 149.625 205.495 149.855 212.530 ;
        RECT 150.915 211.190 151.145 212.530 ;
        RECT 150.880 209.690 151.180 211.190 ;
        RECT 149.590 204.795 149.890 205.495 ;
        RECT 149.625 204.530 149.855 204.795 ;
        RECT 150.915 204.530 151.145 209.690 ;
        RECT 152.205 206.705 152.435 212.530 ;
        RECT 152.170 206.005 152.470 206.705 ;
        RECT 152.205 204.530 152.435 206.005 ;
        RECT 149.905 203.995 150.865 204.325 ;
        RECT 151.195 203.995 152.155 204.325 ;
        RECT 152.845 203.720 153.245 213.340 ;
        RECT 108.515 203.320 153.245 203.720 ;
        RECT 108.515 200.625 153.245 201.025 ;
        RECT 108.515 195.095 108.915 200.625 ;
        RECT 109.735 200.250 110.435 200.320 ;
        RECT 111.025 200.250 111.725 200.320 ;
        RECT 109.605 200.020 110.565 200.250 ;
        RECT 110.895 200.020 111.855 200.250 ;
        RECT 109.325 199.635 109.555 199.860 ;
        RECT 109.290 198.935 109.590 199.635 ;
        RECT 110.615 198.955 110.845 199.860 ;
        RECT 111.905 199.635 112.135 199.860 ;
        RECT 109.325 195.860 109.555 198.935 ;
        RECT 110.580 196.855 110.880 198.955 ;
        RECT 111.870 198.935 112.170 199.635 ;
        RECT 110.615 195.860 110.845 196.855 ;
        RECT 111.905 195.860 112.135 198.935 ;
        RECT 109.605 195.470 110.565 195.700 ;
        RECT 110.895 195.470 111.855 195.700 ;
        RECT 112.545 195.095 112.945 200.625 ;
        RECT 113.765 200.250 114.465 200.320 ;
        RECT 115.055 200.250 115.755 200.320 ;
        RECT 113.635 200.020 114.595 200.250 ;
        RECT 114.925 200.020 115.885 200.250 ;
        RECT 113.355 199.635 113.585 199.860 ;
        RECT 113.320 198.935 113.620 199.635 ;
        RECT 114.645 198.955 114.875 199.860 ;
        RECT 115.935 199.635 116.165 199.860 ;
        RECT 113.355 195.860 113.585 198.935 ;
        RECT 114.610 196.855 114.910 198.955 ;
        RECT 115.900 198.935 116.200 199.635 ;
        RECT 114.645 195.860 114.875 196.855 ;
        RECT 115.935 195.860 116.165 198.935 ;
        RECT 113.635 195.470 114.595 195.700 ;
        RECT 114.925 195.470 115.885 195.700 ;
        RECT 116.575 195.095 116.975 200.625 ;
        RECT 117.795 200.250 118.495 200.320 ;
        RECT 119.085 200.250 119.785 200.320 ;
        RECT 117.665 200.020 118.625 200.250 ;
        RECT 118.955 200.020 119.915 200.250 ;
        RECT 117.385 199.635 117.615 199.860 ;
        RECT 117.350 198.935 117.650 199.635 ;
        RECT 118.675 198.955 118.905 199.860 ;
        RECT 119.965 199.635 120.195 199.860 ;
        RECT 117.385 195.860 117.615 198.935 ;
        RECT 118.640 196.855 118.940 198.955 ;
        RECT 119.930 198.935 120.230 199.635 ;
        RECT 118.675 195.860 118.905 196.855 ;
        RECT 119.965 195.860 120.195 198.935 ;
        RECT 117.665 195.470 118.625 195.700 ;
        RECT 118.955 195.470 119.915 195.700 ;
        RECT 120.605 195.095 121.005 200.625 ;
        RECT 121.825 200.250 122.525 200.320 ;
        RECT 123.115 200.250 123.815 200.320 ;
        RECT 121.695 200.020 122.655 200.250 ;
        RECT 122.985 200.020 123.945 200.250 ;
        RECT 121.415 199.635 121.645 199.860 ;
        RECT 121.380 198.935 121.680 199.635 ;
        RECT 122.705 198.955 122.935 199.860 ;
        RECT 123.995 199.635 124.225 199.860 ;
        RECT 121.415 195.860 121.645 198.935 ;
        RECT 122.670 196.855 122.970 198.955 ;
        RECT 123.960 198.935 124.260 199.635 ;
        RECT 122.705 195.860 122.935 196.855 ;
        RECT 123.995 195.860 124.225 198.935 ;
        RECT 121.695 195.470 122.655 195.700 ;
        RECT 122.985 195.470 123.945 195.700 ;
        RECT 124.635 195.095 125.035 200.625 ;
        RECT 125.855 200.250 126.555 200.320 ;
        RECT 127.145 200.250 127.845 200.320 ;
        RECT 125.725 200.020 126.685 200.250 ;
        RECT 127.015 200.020 127.975 200.250 ;
        RECT 125.445 199.635 125.675 199.860 ;
        RECT 125.410 198.935 125.710 199.635 ;
        RECT 126.735 198.955 126.965 199.860 ;
        RECT 128.025 199.635 128.255 199.860 ;
        RECT 125.445 195.860 125.675 198.935 ;
        RECT 126.700 196.855 127.000 198.955 ;
        RECT 127.990 198.935 128.290 199.635 ;
        RECT 126.735 195.860 126.965 196.855 ;
        RECT 128.025 195.860 128.255 198.935 ;
        RECT 125.725 195.470 126.685 195.700 ;
        RECT 127.015 195.470 127.975 195.700 ;
        RECT 128.665 195.095 129.065 200.625 ;
        RECT 129.885 200.250 130.585 200.320 ;
        RECT 131.175 200.250 131.875 200.320 ;
        RECT 129.755 200.020 130.715 200.250 ;
        RECT 131.045 200.020 132.005 200.250 ;
        RECT 129.475 199.635 129.705 199.860 ;
        RECT 129.440 198.935 129.740 199.635 ;
        RECT 130.765 198.955 130.995 199.860 ;
        RECT 132.055 199.635 132.285 199.860 ;
        RECT 129.475 195.860 129.705 198.935 ;
        RECT 130.730 196.855 131.030 198.955 ;
        RECT 132.020 198.935 132.320 199.635 ;
        RECT 130.765 195.860 130.995 196.855 ;
        RECT 132.055 195.860 132.285 198.935 ;
        RECT 129.755 195.470 130.715 195.700 ;
        RECT 131.045 195.470 132.005 195.700 ;
        RECT 132.695 195.095 133.095 200.625 ;
        RECT 133.915 200.250 134.615 200.320 ;
        RECT 135.205 200.250 135.905 200.320 ;
        RECT 133.785 200.020 134.745 200.250 ;
        RECT 135.075 200.020 136.035 200.250 ;
        RECT 133.505 199.635 133.735 199.860 ;
        RECT 133.470 198.935 133.770 199.635 ;
        RECT 134.795 198.955 135.025 199.860 ;
        RECT 136.085 199.635 136.315 199.860 ;
        RECT 133.505 195.860 133.735 198.935 ;
        RECT 134.760 196.855 135.060 198.955 ;
        RECT 136.050 198.935 136.350 199.635 ;
        RECT 134.795 195.860 135.025 196.855 ;
        RECT 136.085 195.860 136.315 198.935 ;
        RECT 133.785 195.470 134.745 195.700 ;
        RECT 135.075 195.470 136.035 195.700 ;
        RECT 136.725 195.095 137.125 200.625 ;
        RECT 137.945 200.250 138.645 200.320 ;
        RECT 139.235 200.250 139.935 200.320 ;
        RECT 137.815 200.020 138.775 200.250 ;
        RECT 139.105 200.020 140.065 200.250 ;
        RECT 137.535 199.635 137.765 199.860 ;
        RECT 137.500 198.935 137.800 199.635 ;
        RECT 138.825 198.955 139.055 199.860 ;
        RECT 140.115 199.635 140.345 199.860 ;
        RECT 137.535 195.860 137.765 198.935 ;
        RECT 138.790 196.855 139.090 198.955 ;
        RECT 140.080 198.935 140.380 199.635 ;
        RECT 138.825 195.860 139.055 196.855 ;
        RECT 140.115 195.860 140.345 198.935 ;
        RECT 137.815 195.470 138.775 195.700 ;
        RECT 139.105 195.470 140.065 195.700 ;
        RECT 140.755 195.095 141.155 200.625 ;
        RECT 141.975 200.250 142.675 200.320 ;
        RECT 143.265 200.250 143.965 200.320 ;
        RECT 141.845 200.020 142.805 200.250 ;
        RECT 143.135 200.020 144.095 200.250 ;
        RECT 141.565 199.635 141.795 199.860 ;
        RECT 141.530 198.935 141.830 199.635 ;
        RECT 142.855 198.955 143.085 199.860 ;
        RECT 144.145 199.635 144.375 199.860 ;
        RECT 141.565 195.860 141.795 198.935 ;
        RECT 142.820 196.855 143.120 198.955 ;
        RECT 144.110 198.935 144.410 199.635 ;
        RECT 142.855 195.860 143.085 196.855 ;
        RECT 144.145 195.860 144.375 198.935 ;
        RECT 141.845 195.470 142.805 195.700 ;
        RECT 143.135 195.470 144.095 195.700 ;
        RECT 144.785 195.095 145.185 200.625 ;
        RECT 146.005 200.250 146.705 200.320 ;
        RECT 147.295 200.250 147.995 200.320 ;
        RECT 145.875 200.020 146.835 200.250 ;
        RECT 147.165 200.020 148.125 200.250 ;
        RECT 145.595 199.635 145.825 199.860 ;
        RECT 145.560 198.935 145.860 199.635 ;
        RECT 146.885 198.955 147.115 199.860 ;
        RECT 148.175 199.635 148.405 199.860 ;
        RECT 145.595 195.860 145.825 198.935 ;
        RECT 146.850 196.855 147.150 198.955 ;
        RECT 148.140 198.935 148.440 199.635 ;
        RECT 146.885 195.860 147.115 196.855 ;
        RECT 148.175 195.860 148.405 198.935 ;
        RECT 145.875 195.470 146.835 195.700 ;
        RECT 147.165 195.470 148.125 195.700 ;
        RECT 148.815 195.095 149.215 200.625 ;
        RECT 150.035 200.250 150.735 200.320 ;
        RECT 151.325 200.250 152.025 200.320 ;
        RECT 149.905 200.020 150.865 200.250 ;
        RECT 151.195 200.020 152.155 200.250 ;
        RECT 149.625 199.635 149.855 199.860 ;
        RECT 149.590 198.935 149.890 199.635 ;
        RECT 150.915 198.955 151.145 199.860 ;
        RECT 152.205 199.635 152.435 199.860 ;
        RECT 149.625 195.860 149.855 198.935 ;
        RECT 150.880 196.855 151.180 198.955 ;
        RECT 152.170 198.935 152.470 199.635 ;
        RECT 150.915 195.860 151.145 196.855 ;
        RECT 152.205 195.860 152.435 198.935 ;
        RECT 149.905 195.470 150.865 195.700 ;
        RECT 151.195 195.470 152.155 195.700 ;
        RECT 152.845 195.095 153.245 200.625 ;
        RECT 108.515 194.695 153.245 195.095 ;
        RECT 108.515 185.165 108.915 194.695 ;
        RECT 109.605 194.320 110.305 194.390 ;
        RECT 111.155 194.320 111.855 194.390 ;
        RECT 109.605 194.090 110.565 194.320 ;
        RECT 110.895 194.090 111.855 194.320 ;
        RECT 109.325 192.835 109.555 193.930 ;
        RECT 109.290 191.335 109.590 192.835 ;
        RECT 109.325 185.930 109.555 191.335 ;
        RECT 110.615 189.090 110.845 193.930 ;
        RECT 111.905 192.835 112.135 193.930 ;
        RECT 111.870 191.335 112.170 192.835 ;
        RECT 110.580 187.590 110.880 189.090 ;
        RECT 110.615 185.930 110.845 187.590 ;
        RECT 111.905 185.930 112.135 191.335 ;
        RECT 109.605 185.540 110.565 185.770 ;
        RECT 110.895 185.540 111.855 185.770 ;
        RECT 112.545 185.165 112.945 194.695 ;
        RECT 113.635 194.320 114.335 194.390 ;
        RECT 115.185 194.320 115.885 194.390 ;
        RECT 113.635 194.090 114.595 194.320 ;
        RECT 114.925 194.090 115.885 194.320 ;
        RECT 113.355 192.835 113.585 193.930 ;
        RECT 113.320 191.335 113.620 192.835 ;
        RECT 113.355 185.930 113.585 191.335 ;
        RECT 114.645 189.090 114.875 193.930 ;
        RECT 115.935 192.835 116.165 193.930 ;
        RECT 115.900 191.335 116.200 192.835 ;
        RECT 114.610 187.590 114.910 189.090 ;
        RECT 114.645 185.930 114.875 187.590 ;
        RECT 115.935 185.930 116.165 191.335 ;
        RECT 113.635 185.540 114.595 185.770 ;
        RECT 114.925 185.540 115.885 185.770 ;
        RECT 116.575 185.165 116.975 194.695 ;
        RECT 117.665 194.320 118.365 194.390 ;
        RECT 119.215 194.320 119.915 194.390 ;
        RECT 117.665 194.090 118.625 194.320 ;
        RECT 118.955 194.090 119.915 194.320 ;
        RECT 117.385 192.835 117.615 193.930 ;
        RECT 117.350 191.335 117.650 192.835 ;
        RECT 117.385 185.930 117.615 191.335 ;
        RECT 118.675 189.090 118.905 193.930 ;
        RECT 119.965 192.835 120.195 193.930 ;
        RECT 119.930 191.335 120.230 192.835 ;
        RECT 118.640 187.590 118.940 189.090 ;
        RECT 118.675 185.930 118.905 187.590 ;
        RECT 119.965 185.930 120.195 191.335 ;
        RECT 117.665 185.540 118.625 185.770 ;
        RECT 118.955 185.540 119.915 185.770 ;
        RECT 120.605 185.165 121.005 194.695 ;
        RECT 121.695 194.320 122.395 194.390 ;
        RECT 123.245 194.320 123.945 194.390 ;
        RECT 121.695 194.090 122.655 194.320 ;
        RECT 122.985 194.090 123.945 194.320 ;
        RECT 121.415 192.835 121.645 193.930 ;
        RECT 121.380 191.335 121.680 192.835 ;
        RECT 121.415 185.930 121.645 191.335 ;
        RECT 122.705 189.090 122.935 193.930 ;
        RECT 123.995 192.835 124.225 193.930 ;
        RECT 123.960 191.335 124.260 192.835 ;
        RECT 122.670 187.590 122.970 189.090 ;
        RECT 122.705 185.930 122.935 187.590 ;
        RECT 123.995 185.930 124.225 191.335 ;
        RECT 121.695 185.540 122.655 185.770 ;
        RECT 122.985 185.540 123.945 185.770 ;
        RECT 124.635 185.165 125.035 194.695 ;
        RECT 125.725 194.320 126.425 194.390 ;
        RECT 127.275 194.320 127.975 194.390 ;
        RECT 125.725 194.090 126.685 194.320 ;
        RECT 127.015 194.090 127.975 194.320 ;
        RECT 125.445 192.835 125.675 193.930 ;
        RECT 125.410 191.335 125.710 192.835 ;
        RECT 125.445 185.930 125.675 191.335 ;
        RECT 126.735 189.090 126.965 193.930 ;
        RECT 128.025 192.835 128.255 193.930 ;
        RECT 127.990 191.335 128.290 192.835 ;
        RECT 126.700 187.590 127.000 189.090 ;
        RECT 126.735 185.930 126.965 187.590 ;
        RECT 128.025 185.930 128.255 191.335 ;
        RECT 125.725 185.540 126.685 185.770 ;
        RECT 127.015 185.540 127.975 185.770 ;
        RECT 128.665 185.165 129.065 194.695 ;
        RECT 129.755 194.320 130.455 194.390 ;
        RECT 131.305 194.320 132.005 194.390 ;
        RECT 129.755 194.090 130.715 194.320 ;
        RECT 131.045 194.090 132.005 194.320 ;
        RECT 129.475 192.835 129.705 193.930 ;
        RECT 129.440 191.335 129.740 192.835 ;
        RECT 129.475 185.930 129.705 191.335 ;
        RECT 130.765 189.090 130.995 193.930 ;
        RECT 132.055 192.835 132.285 193.930 ;
        RECT 132.020 191.335 132.320 192.835 ;
        RECT 130.730 187.590 131.030 189.090 ;
        RECT 130.765 185.930 130.995 187.590 ;
        RECT 132.055 185.930 132.285 191.335 ;
        RECT 129.755 185.540 130.715 185.770 ;
        RECT 131.045 185.540 132.005 185.770 ;
        RECT 132.695 185.165 133.095 194.695 ;
        RECT 133.785 194.320 134.485 194.390 ;
        RECT 135.335 194.320 136.035 194.390 ;
        RECT 133.785 194.090 134.745 194.320 ;
        RECT 135.075 194.090 136.035 194.320 ;
        RECT 133.505 192.835 133.735 193.930 ;
        RECT 133.470 191.335 133.770 192.835 ;
        RECT 133.505 185.930 133.735 191.335 ;
        RECT 134.795 189.090 135.025 193.930 ;
        RECT 136.085 192.835 136.315 193.930 ;
        RECT 136.050 191.335 136.350 192.835 ;
        RECT 134.760 187.590 135.060 189.090 ;
        RECT 134.795 185.930 135.025 187.590 ;
        RECT 136.085 185.930 136.315 191.335 ;
        RECT 133.785 185.540 134.745 185.770 ;
        RECT 135.075 185.540 136.035 185.770 ;
        RECT 136.725 185.165 137.125 194.695 ;
        RECT 137.815 194.320 138.515 194.390 ;
        RECT 139.365 194.320 140.065 194.390 ;
        RECT 137.815 194.090 138.775 194.320 ;
        RECT 139.105 194.090 140.065 194.320 ;
        RECT 137.535 192.835 137.765 193.930 ;
        RECT 137.500 191.335 137.800 192.835 ;
        RECT 137.535 185.930 137.765 191.335 ;
        RECT 138.825 189.090 139.055 193.930 ;
        RECT 140.115 192.835 140.345 193.930 ;
        RECT 140.080 191.335 140.380 192.835 ;
        RECT 138.790 187.590 139.090 189.090 ;
        RECT 138.825 185.930 139.055 187.590 ;
        RECT 140.115 185.930 140.345 191.335 ;
        RECT 137.815 185.540 138.775 185.770 ;
        RECT 139.105 185.540 140.065 185.770 ;
        RECT 140.755 185.165 141.155 194.695 ;
        RECT 141.845 194.320 142.545 194.390 ;
        RECT 143.395 194.320 144.095 194.390 ;
        RECT 141.845 194.090 142.805 194.320 ;
        RECT 143.135 194.090 144.095 194.320 ;
        RECT 141.565 192.835 141.795 193.930 ;
        RECT 141.530 191.335 141.830 192.835 ;
        RECT 141.565 185.930 141.795 191.335 ;
        RECT 142.855 189.090 143.085 193.930 ;
        RECT 144.145 192.835 144.375 193.930 ;
        RECT 144.110 191.335 144.410 192.835 ;
        RECT 142.820 187.590 143.120 189.090 ;
        RECT 142.855 185.930 143.085 187.590 ;
        RECT 144.145 185.930 144.375 191.335 ;
        RECT 141.845 185.540 142.805 185.770 ;
        RECT 143.135 185.540 144.095 185.770 ;
        RECT 144.785 185.165 145.185 194.695 ;
        RECT 145.875 194.320 146.575 194.390 ;
        RECT 147.425 194.320 148.125 194.390 ;
        RECT 145.875 194.090 146.835 194.320 ;
        RECT 147.165 194.090 148.125 194.320 ;
        RECT 145.595 192.835 145.825 193.930 ;
        RECT 145.560 191.335 145.860 192.835 ;
        RECT 145.595 185.930 145.825 191.335 ;
        RECT 146.885 189.090 147.115 193.930 ;
        RECT 148.175 192.835 148.405 193.930 ;
        RECT 148.140 191.335 148.440 192.835 ;
        RECT 146.850 187.590 147.150 189.090 ;
        RECT 146.885 185.930 147.115 187.590 ;
        RECT 148.175 185.930 148.405 191.335 ;
        RECT 145.875 185.540 146.835 185.770 ;
        RECT 147.165 185.540 148.125 185.770 ;
        RECT 148.815 185.165 149.215 194.695 ;
        RECT 149.905 194.320 150.605 194.390 ;
        RECT 151.455 194.320 152.155 194.390 ;
        RECT 149.905 194.090 150.865 194.320 ;
        RECT 151.195 194.090 152.155 194.320 ;
        RECT 149.625 192.835 149.855 193.930 ;
        RECT 149.590 191.335 149.890 192.835 ;
        RECT 149.625 185.930 149.855 191.335 ;
        RECT 150.915 189.090 151.145 193.930 ;
        RECT 152.205 192.835 152.435 193.930 ;
        RECT 152.170 191.335 152.470 192.835 ;
        RECT 150.880 187.590 151.180 189.090 ;
        RECT 150.915 185.930 151.145 187.590 ;
        RECT 152.205 185.930 152.435 191.335 ;
        RECT 152.845 187.965 153.245 194.695 ;
        RECT 149.905 185.540 150.865 185.770 ;
        RECT 151.195 185.540 152.155 185.770 ;
        RECT 152.845 185.165 155.165 187.965 ;
        RECT 108.515 184.765 155.165 185.165 ;
        RECT 63.895 181.400 64.595 182.400 ;
        RECT 77.595 182.370 78.595 182.605 ;
        RECT 77.595 181.195 78.595 181.430 ;
        RECT 80.185 181.400 81.755 182.400 ;
        RECT 83.345 182.370 84.345 182.605 ;
        RECT 83.345 181.195 84.345 181.430 ;
        RECT 97.345 181.400 98.045 182.400 ;
        RECT 64.175 180.965 80.135 181.195 ;
        RECT 81.805 180.965 97.765 181.195 ;
        RECT 77.595 180.730 78.595 180.965 ;
        RECT 83.345 180.730 84.345 180.965 ;
        RECT 98.485 180.110 155.900 182.710 ;
        RECT 77.595 179.815 78.595 180.050 ;
        RECT 83.345 179.815 84.345 180.050 ;
        RECT 64.175 179.585 80.135 179.815 ;
        RECT 81.805 179.585 97.765 179.815 ;
        RECT 63.895 178.380 64.595 179.380 ;
        RECT 77.595 179.350 78.595 179.585 ;
        RECT 77.595 178.175 78.595 178.410 ;
        RECT 80.185 178.380 81.755 179.380 ;
        RECT 83.345 179.350 84.345 179.585 ;
        RECT 83.345 178.175 84.345 178.410 ;
        RECT 97.345 178.380 98.045 179.380 ;
        RECT 64.175 177.945 80.135 178.175 ;
        RECT 81.805 177.945 97.765 178.175 ;
        RECT 77.595 177.710 78.595 177.945 ;
        RECT 83.345 177.710 84.345 177.945 ;
        RECT 77.595 176.795 78.595 177.030 ;
        RECT 83.345 176.795 84.345 177.030 ;
        RECT 64.175 176.565 80.135 176.795 ;
        RECT 81.805 176.565 97.765 176.795 ;
        RECT 63.895 175.360 64.595 176.360 ;
        RECT 77.595 176.330 78.595 176.565 ;
        RECT 77.595 175.155 78.595 175.390 ;
        RECT 80.185 175.360 81.755 176.360 ;
        RECT 83.345 176.330 84.345 176.565 ;
        RECT 83.345 175.155 84.345 175.390 ;
        RECT 97.345 175.360 98.045 176.360 ;
        RECT 64.175 174.925 80.135 175.155 ;
        RECT 81.805 174.925 97.765 175.155 ;
        RECT 77.595 174.690 78.595 174.925 ;
        RECT 83.345 174.690 84.345 174.925 ;
        RECT 64.175 173.545 80.135 173.775 ;
        RECT 81.805 173.545 97.765 173.775 ;
        RECT 63.895 172.340 64.125 173.340 ;
        RECT 80.185 172.340 81.755 173.340 ;
        RECT 97.815 172.340 98.045 173.340 ;
        RECT 64.175 171.905 80.135 172.135 ;
        RECT 81.805 171.905 97.765 172.135 ;
        RECT 98.485 171.445 100.480 180.110 ;
        RECT 62.865 160.555 100.480 171.445 ;
        RECT 5.910 143.155 58.705 143.745 ;
        RECT 5.910 140.725 23.785 143.155 ;
        RECT 24.505 143.045 25.505 143.155 ;
        RECT 24.255 142.435 57.645 142.665 ;
        RECT 24.255 141.275 24.485 142.435 ;
        RECT 28.015 141.965 29.015 142.435 ;
        RECT 32.545 141.275 32.775 142.435 ;
        RECT 36.305 141.965 37.305 142.435 ;
        RECT 40.835 141.275 41.065 142.435 ;
        RECT 44.595 141.965 45.595 142.435 ;
        RECT 49.125 141.275 49.355 142.435 ;
        RECT 52.885 141.965 53.885 142.435 ;
        RECT 57.415 141.275 57.645 142.435 ;
        RECT 24.535 140.885 32.495 141.115 ;
        RECT 32.825 140.885 40.785 141.115 ;
        RECT 41.115 140.885 49.075 141.115 ;
        RECT 49.405 140.885 57.365 141.115 ;
        RECT 5.910 139.725 24.955 140.725 ;
        RECT 32.545 139.725 32.775 140.725 ;
        RECT 40.835 139.725 41.065 140.725 ;
        RECT 49.125 139.725 49.355 140.725 ;
        RECT 56.545 139.725 57.645 140.725 ;
        RECT 5.910 139.175 23.785 139.725 ;
        RECT 24.535 139.335 32.495 139.565 ;
        RECT 32.825 139.335 40.785 139.565 ;
        RECT 41.115 139.335 49.075 139.565 ;
        RECT 49.405 139.335 57.365 139.565 ;
        RECT 5.910 138.175 24.955 139.175 ;
        RECT 32.545 138.175 32.775 139.175 ;
        RECT 40.835 138.175 41.065 139.175 ;
        RECT 49.125 138.175 49.355 139.175 ;
        RECT 53.035 138.175 57.645 139.175 ;
        RECT 5.910 137.925 23.785 138.175 ;
        RECT 5.910 137.075 9.990 137.925 ;
        RECT 11.145 137.465 11.845 137.535 ;
        RECT 14.080 137.465 14.780 137.535 ;
        RECT 15.370 137.465 16.070 137.535 ;
        RECT 18.305 137.465 19.005 137.535 ;
        RECT 11.015 137.235 11.975 137.465 ;
        RECT 13.950 137.235 14.910 137.465 ;
        RECT 15.240 137.235 16.200 137.465 ;
        RECT 18.175 137.235 19.135 137.465 ;
        RECT 5.910 136.075 10.965 137.075 ;
        RECT 12.025 136.925 12.255 137.075 ;
        RECT 11.990 136.225 12.290 136.925 ;
        RECT 12.025 136.075 12.255 136.225 ;
        RECT 5.910 135.225 9.990 136.075 ;
        RECT 13.670 135.825 13.900 137.075 ;
        RECT 14.960 136.925 15.190 137.075 ;
        RECT 16.250 136.925 16.480 137.075 ;
        RECT 14.925 136.225 15.225 136.925 ;
        RECT 16.215 136.225 16.515 136.925 ;
        RECT 14.960 136.075 15.190 136.225 ;
        RECT 16.250 136.075 16.480 136.225 ;
        RECT 13.435 135.525 14.135 135.825 ;
        RECT 17.895 135.225 18.125 137.075 ;
        RECT 19.185 136.775 19.415 137.075 ;
        RECT 19.150 136.075 19.450 136.775 ;
        RECT 20.160 135.745 23.785 137.925 ;
        RECT 24.535 137.785 32.495 138.015 ;
        RECT 32.825 137.785 40.785 138.015 ;
        RECT 41.115 137.785 49.075 138.015 ;
        RECT 49.405 137.785 57.365 138.015 ;
        RECT 24.255 136.465 24.485 137.625 ;
        RECT 28.015 136.465 29.015 136.935 ;
        RECT 32.545 136.465 32.775 137.625 ;
        RECT 36.305 136.465 37.305 136.935 ;
        RECT 40.835 136.465 41.065 137.625 ;
        RECT 44.595 136.465 45.595 136.935 ;
        RECT 49.125 136.465 49.355 137.625 ;
        RECT 52.885 136.465 53.885 136.935 ;
        RECT 57.415 136.465 57.645 137.625 ;
        RECT 24.255 136.235 57.645 136.465 ;
        RECT 24.505 135.745 25.505 135.855 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 20.160 135.225 58.705 135.745 ;
        RECT 5.910 132.225 58.705 135.225 ;
        RECT 62.865 139.455 69.970 160.555 ;
        RECT 71.220 157.040 89.820 159.315 ;
        RECT 71.220 142.990 73.495 157.040 ;
        RECT 76.385 157.030 77.215 157.040 ;
        RECT 80.105 157.030 80.935 157.040 ;
        RECT 83.825 157.030 84.655 157.040 ;
        RECT 74.940 154.420 86.100 155.595 ;
        RECT 74.940 153.050 76.115 154.420 ;
        RECT 76.385 153.310 77.215 154.140 ;
        RECT 77.485 153.050 79.835 154.420 ;
        RECT 80.105 153.310 80.935 154.140 ;
        RECT 81.205 153.050 83.555 154.420 ;
        RECT 83.825 153.310 84.655 154.140 ;
        RECT 84.925 153.050 86.100 154.420 ;
        RECT 74.940 150.700 86.100 153.050 ;
        RECT 74.940 149.330 76.115 150.700 ;
        RECT 76.385 149.590 77.215 150.420 ;
        RECT 77.485 149.330 79.835 150.700 ;
        RECT 80.105 149.590 80.935 150.420 ;
        RECT 81.205 149.330 83.555 150.700 ;
        RECT 83.825 149.590 84.655 150.420 ;
        RECT 84.925 149.330 86.100 150.700 ;
        RECT 74.940 146.980 86.100 149.330 ;
        RECT 74.940 145.610 76.115 146.980 ;
        RECT 76.385 145.870 77.215 146.700 ;
        RECT 77.485 145.610 79.835 146.980 ;
        RECT 80.105 145.870 80.935 146.700 ;
        RECT 81.205 145.610 83.555 146.980 ;
        RECT 83.825 145.870 84.655 146.700 ;
        RECT 84.925 145.610 86.100 146.980 ;
        RECT 74.940 144.435 86.100 145.610 ;
        RECT 87.545 142.990 89.820 157.040 ;
        RECT 71.220 140.715 89.820 142.990 ;
        RECT 91.070 139.455 100.480 160.555 ;
        RECT 101.935 176.325 152.755 178.210 ;
        RECT 101.935 174.870 114.420 176.325 ;
        RECT 115.200 175.635 118.030 176.165 ;
        RECT 119.820 175.635 122.650 176.165 ;
        RECT 124.440 175.635 127.270 176.165 ;
        RECT 129.060 175.635 131.890 176.165 ;
        RECT 133.680 175.635 136.510 176.165 ;
        RECT 138.300 175.635 141.130 176.165 ;
        RECT 142.920 175.635 145.750 176.165 ;
        RECT 147.540 175.635 150.370 176.165 ;
        RECT 114.920 174.870 115.150 175.475 ;
        RECT 101.935 172.215 115.185 174.870 ;
        RECT 101.935 162.685 103.025 172.215 ;
        RECT 103.715 171.610 104.675 171.840 ;
        RECT 105.005 171.610 105.965 171.840 ;
        RECT 103.435 170.840 103.665 171.450 ;
        RECT 103.400 168.540 103.700 170.840 ;
        RECT 103.435 163.450 103.665 168.540 ;
        RECT 104.725 167.140 104.955 171.450 ;
        RECT 106.015 170.840 106.245 171.450 ;
        RECT 105.980 168.540 106.280 170.840 ;
        RECT 104.690 164.840 104.990 167.140 ;
        RECT 104.725 163.450 104.955 164.840 ;
        RECT 106.015 163.450 106.245 168.540 ;
        RECT 103.715 163.060 104.675 163.290 ;
        RECT 105.005 163.060 105.965 163.290 ;
        RECT 103.715 162.990 104.415 163.060 ;
        RECT 105.265 162.990 105.965 163.060 ;
        RECT 106.655 162.685 107.055 172.215 ;
        RECT 110.685 172.070 115.185 172.215 ;
        RECT 107.745 171.610 108.705 171.840 ;
        RECT 109.035 171.610 109.995 171.840 ;
        RECT 107.465 170.840 107.695 171.450 ;
        RECT 107.430 168.540 107.730 170.840 ;
        RECT 107.465 163.450 107.695 168.540 ;
        RECT 108.755 167.140 108.985 171.450 ;
        RECT 110.045 170.840 110.275 171.450 ;
        RECT 110.010 168.540 110.310 170.840 ;
        RECT 108.720 164.840 109.020 167.140 ;
        RECT 108.755 163.450 108.985 164.840 ;
        RECT 110.045 163.450 110.275 168.540 ;
        RECT 110.685 166.625 114.420 172.070 ;
        RECT 114.920 167.475 115.150 172.070 ;
        RECT 115.710 170.895 115.940 175.475 ;
        RECT 116.500 174.870 116.730 175.475 ;
        RECT 116.465 172.070 116.765 174.870 ;
        RECT 115.675 168.095 115.975 170.895 ;
        RECT 115.710 167.475 115.940 168.095 ;
        RECT 116.500 167.475 116.730 172.070 ;
        RECT 117.290 170.895 117.520 175.475 ;
        RECT 118.080 174.870 118.310 175.475 ;
        RECT 119.540 174.870 119.770 175.475 ;
        RECT 118.045 172.070 118.345 174.870 ;
        RECT 119.505 172.070 119.805 174.870 ;
        RECT 117.255 168.095 117.555 170.895 ;
        RECT 117.290 167.475 117.520 168.095 ;
        RECT 118.080 167.475 118.310 172.070 ;
        RECT 119.540 167.475 119.770 172.070 ;
        RECT 120.330 170.895 120.560 175.475 ;
        RECT 121.120 174.870 121.350 175.475 ;
        RECT 121.085 172.070 121.385 174.870 ;
        RECT 120.295 168.095 120.595 170.895 ;
        RECT 120.330 167.475 120.560 168.095 ;
        RECT 121.120 167.475 121.350 172.070 ;
        RECT 121.910 170.895 122.140 175.475 ;
        RECT 122.700 174.870 122.930 175.475 ;
        RECT 124.160 174.870 124.390 175.475 ;
        RECT 122.665 172.070 122.965 174.870 ;
        RECT 124.125 172.070 124.425 174.870 ;
        RECT 121.875 168.095 122.175 170.895 ;
        RECT 121.910 167.475 122.140 168.095 ;
        RECT 122.700 167.475 122.930 172.070 ;
        RECT 124.160 167.475 124.390 172.070 ;
        RECT 124.950 170.895 125.180 175.475 ;
        RECT 125.740 174.870 125.970 175.475 ;
        RECT 125.705 172.070 126.005 174.870 ;
        RECT 124.915 168.095 125.215 170.895 ;
        RECT 124.950 167.475 125.180 168.095 ;
        RECT 125.740 167.475 125.970 172.070 ;
        RECT 126.530 170.895 126.760 175.475 ;
        RECT 127.320 174.870 127.550 175.475 ;
        RECT 128.780 174.870 129.010 175.475 ;
        RECT 127.285 172.070 127.585 174.870 ;
        RECT 128.745 172.070 129.045 174.870 ;
        RECT 126.495 168.095 126.795 170.895 ;
        RECT 126.530 167.475 126.760 168.095 ;
        RECT 127.320 167.475 127.550 172.070 ;
        RECT 128.780 167.475 129.010 172.070 ;
        RECT 129.570 170.895 129.800 175.475 ;
        RECT 130.360 174.870 130.590 175.475 ;
        RECT 130.325 172.070 130.625 174.870 ;
        RECT 129.535 168.095 129.835 170.895 ;
        RECT 129.570 167.475 129.800 168.095 ;
        RECT 130.360 167.475 130.590 172.070 ;
        RECT 131.150 170.895 131.380 175.475 ;
        RECT 131.940 174.870 132.170 175.475 ;
        RECT 133.400 174.870 133.630 175.475 ;
        RECT 131.905 172.070 132.205 174.870 ;
        RECT 133.365 172.070 133.665 174.870 ;
        RECT 131.115 168.095 131.415 170.895 ;
        RECT 131.150 167.475 131.380 168.095 ;
        RECT 131.940 167.475 132.170 172.070 ;
        RECT 133.400 167.475 133.630 172.070 ;
        RECT 134.190 170.895 134.420 175.475 ;
        RECT 134.980 174.870 135.210 175.475 ;
        RECT 134.945 172.070 135.245 174.870 ;
        RECT 134.155 168.095 134.455 170.895 ;
        RECT 134.190 167.475 134.420 168.095 ;
        RECT 134.980 167.475 135.210 172.070 ;
        RECT 135.770 170.895 136.000 175.475 ;
        RECT 136.560 174.870 136.790 175.475 ;
        RECT 138.020 174.870 138.250 175.475 ;
        RECT 136.525 172.070 136.825 174.870 ;
        RECT 137.985 172.070 138.285 174.870 ;
        RECT 135.735 168.095 136.035 170.895 ;
        RECT 135.770 167.475 136.000 168.095 ;
        RECT 136.560 167.475 136.790 172.070 ;
        RECT 138.020 167.475 138.250 172.070 ;
        RECT 138.810 170.895 139.040 175.475 ;
        RECT 139.600 174.870 139.830 175.475 ;
        RECT 139.565 172.070 139.865 174.870 ;
        RECT 138.775 168.095 139.075 170.895 ;
        RECT 138.810 167.475 139.040 168.095 ;
        RECT 139.600 167.475 139.830 172.070 ;
        RECT 140.390 170.895 140.620 175.475 ;
        RECT 141.180 174.870 141.410 175.475 ;
        RECT 142.640 174.870 142.870 175.475 ;
        RECT 141.145 172.070 141.445 174.870 ;
        RECT 142.605 172.070 142.905 174.870 ;
        RECT 140.355 168.095 140.655 170.895 ;
        RECT 140.390 167.475 140.620 168.095 ;
        RECT 141.180 167.475 141.410 172.070 ;
        RECT 142.640 167.475 142.870 172.070 ;
        RECT 143.430 170.895 143.660 175.475 ;
        RECT 144.220 174.870 144.450 175.475 ;
        RECT 144.185 172.070 144.485 174.870 ;
        RECT 143.395 168.095 143.695 170.895 ;
        RECT 143.430 167.475 143.660 168.095 ;
        RECT 144.220 167.475 144.450 172.070 ;
        RECT 145.010 170.895 145.240 175.475 ;
        RECT 145.800 174.870 146.030 175.475 ;
        RECT 147.260 174.870 147.490 175.475 ;
        RECT 145.765 172.070 146.065 174.870 ;
        RECT 147.225 172.070 147.525 174.870 ;
        RECT 144.975 168.095 145.275 170.895 ;
        RECT 145.010 167.475 145.240 168.095 ;
        RECT 145.800 167.475 146.030 172.070 ;
        RECT 147.260 167.475 147.490 172.070 ;
        RECT 148.050 170.895 148.280 175.475 ;
        RECT 148.840 174.870 149.070 175.475 ;
        RECT 148.805 172.070 149.105 174.870 ;
        RECT 148.015 168.095 148.315 170.895 ;
        RECT 148.050 167.475 148.280 168.095 ;
        RECT 148.840 167.475 149.070 172.070 ;
        RECT 149.630 170.895 149.860 175.475 ;
        RECT 150.420 174.870 150.650 175.475 ;
        RECT 150.385 172.070 150.685 174.870 ;
        RECT 149.595 168.095 149.895 170.895 ;
        RECT 149.630 167.475 149.860 168.095 ;
        RECT 150.420 167.475 150.650 172.070 ;
        RECT 115.200 167.085 115.660 167.315 ;
        RECT 115.990 167.085 116.450 167.315 ;
        RECT 116.780 167.085 117.240 167.315 ;
        RECT 117.570 167.085 118.030 167.315 ;
        RECT 119.820 167.085 120.280 167.315 ;
        RECT 120.610 167.085 121.070 167.315 ;
        RECT 121.400 167.085 121.860 167.315 ;
        RECT 122.190 167.085 122.650 167.315 ;
        RECT 124.440 167.085 124.900 167.315 ;
        RECT 125.230 167.085 125.690 167.315 ;
        RECT 126.020 167.085 126.480 167.315 ;
        RECT 126.810 167.085 127.270 167.315 ;
        RECT 129.060 167.085 129.520 167.315 ;
        RECT 129.850 167.085 130.310 167.315 ;
        RECT 130.640 167.085 131.100 167.315 ;
        RECT 131.430 167.085 131.890 167.315 ;
        RECT 133.680 167.085 134.140 167.315 ;
        RECT 134.470 167.085 134.930 167.315 ;
        RECT 135.260 167.085 135.720 167.315 ;
        RECT 136.050 167.085 136.510 167.315 ;
        RECT 138.300 167.085 138.760 167.315 ;
        RECT 139.090 167.085 139.550 167.315 ;
        RECT 139.880 167.085 140.340 167.315 ;
        RECT 140.670 167.085 141.130 167.315 ;
        RECT 142.920 167.085 143.380 167.315 ;
        RECT 143.710 167.085 144.170 167.315 ;
        RECT 144.500 167.085 144.960 167.315 ;
        RECT 145.290 167.085 145.750 167.315 ;
        RECT 147.540 167.085 148.000 167.315 ;
        RECT 148.330 167.085 148.790 167.315 ;
        RECT 149.120 167.085 149.580 167.315 ;
        RECT 149.910 167.085 150.370 167.315 ;
        RECT 151.150 166.625 152.755 176.325 ;
        RECT 110.685 166.035 152.755 166.625 ;
        RECT 107.745 163.060 108.705 163.290 ;
        RECT 109.035 163.060 109.995 163.290 ;
        RECT 107.745 162.990 108.445 163.060 ;
        RECT 109.295 162.990 109.995 163.060 ;
        RECT 110.685 162.685 114.420 166.035 ;
        RECT 134.745 165.030 135.445 165.080 ;
        RECT 146.905 165.030 147.605 165.080 ;
        RECT 134.745 164.430 147.605 165.030 ;
        RECT 134.745 164.380 135.445 164.430 ;
        RECT 146.905 164.380 147.605 164.430 ;
        RECT 133.735 163.740 134.435 163.790 ;
        RECT 143.985 163.740 144.685 163.790 ;
        RECT 133.735 163.140 144.685 163.740 ;
        RECT 133.735 163.090 134.435 163.140 ;
        RECT 143.985 163.090 144.685 163.140 ;
        RECT 101.935 162.285 114.420 162.685 ;
        RECT 101.935 158.755 103.025 162.285 ;
        RECT 103.435 160.445 103.665 161.520 ;
        RECT 103.400 159.745 103.700 160.445 ;
        RECT 103.435 159.520 103.665 159.745 ;
        RECT 104.725 159.520 104.955 162.285 ;
        RECT 106.015 160.445 106.245 161.520 ;
        RECT 105.980 159.745 106.280 160.445 ;
        RECT 106.015 159.520 106.245 159.745 ;
        RECT 103.715 159.130 104.675 159.360 ;
        RECT 105.005 159.130 105.965 159.360 ;
        RECT 103.845 159.060 104.545 159.130 ;
        RECT 105.135 159.060 105.835 159.130 ;
        RECT 106.655 158.755 107.055 162.285 ;
        RECT 107.465 160.445 107.695 161.520 ;
        RECT 107.430 159.745 107.730 160.445 ;
        RECT 107.465 159.520 107.695 159.745 ;
        RECT 108.755 159.520 108.985 162.285 ;
        RECT 110.045 160.445 110.275 161.520 ;
        RECT 110.010 159.745 110.310 160.445 ;
        RECT 110.045 159.520 110.275 159.745 ;
        RECT 107.745 159.130 108.705 159.360 ;
        RECT 109.035 159.130 109.995 159.360 ;
        RECT 107.875 159.060 108.575 159.130 ;
        RECT 109.165 159.060 109.865 159.130 ;
        RECT 110.685 158.755 114.420 162.285 ;
        RECT 136.825 162.330 137.525 162.400 ;
        RECT 143.985 162.330 144.685 162.400 ;
        RECT 136.825 161.730 144.685 162.330 ;
        RECT 136.825 161.700 137.525 161.730 ;
        RECT 143.985 161.700 144.685 161.730 ;
        RECT 134.745 160.160 135.445 160.210 ;
        RECT 145.575 160.160 146.275 160.210 ;
        RECT 134.745 159.560 146.275 160.160 ;
        RECT 134.745 159.510 135.445 159.560 ;
        RECT 145.575 159.510 146.275 159.560 ;
        RECT 101.935 157.850 114.420 158.755 ;
        RECT 141.665 159.150 142.365 159.200 ;
        RECT 148.605 159.150 149.305 159.200 ;
        RECT 141.665 158.550 149.305 159.150 ;
        RECT 141.665 158.500 142.365 158.550 ;
        RECT 148.605 158.500 149.305 158.550 ;
        RECT 153.960 158.060 155.900 180.110 ;
        RECT 115.985 156.185 155.900 158.060 ;
        RECT 115.985 156.060 116.575 156.185 ;
        RECT 102.625 155.660 116.575 156.060 ;
        RECT 102.625 152.040 103.025 155.660 ;
        RECT 103.715 155.055 104.675 155.385 ;
        RECT 105.005 155.055 105.965 155.385 ;
        RECT 103.435 153.515 103.665 154.850 ;
        RECT 103.400 152.815 103.700 153.515 ;
        RECT 104.725 152.040 104.955 154.850 ;
        RECT 106.015 154.585 106.245 154.850 ;
        RECT 105.980 153.885 106.280 154.585 ;
        RECT 106.015 152.850 106.245 153.885 ;
        RECT 106.655 152.040 107.055 155.660 ;
        RECT 107.745 155.055 108.705 155.385 ;
        RECT 109.035 155.055 109.995 155.385 ;
        RECT 107.465 153.515 107.695 154.850 ;
        RECT 107.430 152.815 107.730 153.515 ;
        RECT 108.755 152.040 108.985 154.850 ;
        RECT 110.045 154.585 110.275 154.850 ;
        RECT 110.010 153.885 110.310 154.585 ;
        RECT 110.045 152.850 110.275 153.885 ;
        RECT 110.685 152.040 116.575 155.660 ;
        RECT 102.625 151.550 116.575 152.040 ;
        RECT 102.625 142.020 103.025 151.550 ;
        RECT 103.715 151.035 104.675 151.365 ;
        RECT 105.005 151.035 105.965 151.365 ;
        RECT 103.435 145.785 103.665 150.830 ;
        RECT 104.725 149.485 104.955 150.830 ;
        RECT 104.690 147.185 104.990 149.485 ;
        RECT 103.400 143.485 103.700 145.785 ;
        RECT 103.435 142.830 103.665 143.485 ;
        RECT 104.725 142.830 104.955 147.185 ;
        RECT 106.015 145.785 106.245 150.830 ;
        RECT 105.980 143.485 106.280 145.785 ;
        RECT 106.015 142.830 106.245 143.485 ;
        RECT 103.715 142.395 104.675 142.625 ;
        RECT 105.005 142.395 105.965 142.625 ;
        RECT 106.655 142.020 107.055 151.550 ;
        RECT 107.745 151.035 108.705 151.365 ;
        RECT 109.035 151.035 109.995 151.365 ;
        RECT 107.465 145.785 107.695 150.830 ;
        RECT 108.755 149.485 108.985 150.830 ;
        RECT 108.720 147.185 109.020 149.485 ;
        RECT 107.430 143.485 107.730 145.785 ;
        RECT 107.465 142.830 107.695 143.485 ;
        RECT 108.755 142.830 108.985 147.185 ;
        RECT 110.045 145.785 110.275 150.830 ;
        RECT 110.010 143.485 110.310 145.785 ;
        RECT 110.045 142.830 110.275 143.485 ;
        RECT 107.745 142.395 108.705 142.625 ;
        RECT 109.035 142.395 109.995 142.625 ;
        RECT 110.685 142.020 116.575 151.550 ;
        RECT 117.160 142.145 119.265 155.605 ;
        RECT 122.405 146.245 124.510 155.605 ;
        RECT 125.090 146.825 127.195 155.605 ;
        RECT 130.335 146.825 132.440 155.605 ;
        RECT 133.020 154.960 135.125 155.660 ;
        RECT 133.020 152.675 135.125 154.435 ;
        RECT 138.265 153.845 140.370 155.605 ;
        RECT 133.020 151.450 135.125 152.150 ;
        RECT 138.265 151.505 140.370 153.265 ;
        RECT 140.950 152.675 143.055 156.185 ;
        RECT 146.195 152.675 148.300 156.185 ;
        RECT 140.950 151.460 143.055 152.160 ;
        RECT 133.020 150.280 135.125 150.980 ;
        RECT 133.020 149.110 135.125 149.810 ;
        RECT 138.265 149.165 140.370 150.925 ;
        RECT 140.950 149.165 143.055 150.925 ;
        RECT 146.195 150.335 148.300 152.095 ;
        RECT 133.020 146.825 135.125 148.585 ;
        RECT 138.265 146.825 140.370 148.585 ;
        RECT 140.950 146.825 143.055 148.585 ;
        RECT 146.195 147.995 148.300 149.755 ;
        RECT 122.405 142.145 127.195 146.245 ;
        RECT 130.335 142.145 132.440 146.245 ;
        RECT 133.020 142.145 135.125 146.245 ;
        RECT 138.265 142.145 140.370 146.245 ;
        RECT 140.950 144.485 143.055 146.245 ;
        RECT 146.195 145.655 148.300 147.415 ;
        RECT 140.950 143.290 143.055 143.990 ;
        RECT 146.195 143.315 148.300 145.075 ;
        RECT 140.950 142.040 143.055 142.740 ;
        RECT 146.195 142.080 148.300 142.780 ;
        RECT 102.625 141.620 116.575 142.020 ;
        RECT 62.865 130.990 100.480 139.455 ;
        RECT 111.085 141.565 116.575 141.620 ;
        RECT 148.885 141.565 155.900 156.185 ;
        RECT 111.085 137.690 155.900 141.565 ;
        RECT 111.085 130.990 135.120 137.690 ;
        RECT 62.865 127.485 135.120 130.990 ;
        RECT 138.080 134.100 145.960 137.690 ;
        RECT 138.080 130.310 138.670 134.100 ;
        RECT 139.615 133.640 140.315 133.760 ;
        RECT 140.905 133.640 141.605 133.760 ;
        RECT 139.485 133.410 140.445 133.640 ;
        RECT 140.775 133.410 141.735 133.640 ;
        RECT 139.205 132.990 139.435 133.205 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 139.205 131.205 139.435 131.390 ;
        RECT 140.495 130.310 140.725 133.205 ;
        RECT 141.785 132.990 142.015 133.205 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 143.315 132.640 143.545 133.205 ;
        RECT 143.280 131.940 143.580 132.640 ;
        RECT 141.785 131.205 142.015 131.390 ;
        RECT 143.315 131.205 143.545 131.940 ;
        RECT 144.605 131.205 144.835 134.100 ;
        RECT 143.595 130.770 144.555 131.000 ;
        RECT 143.725 130.700 144.425 130.770 ;
        RECT 145.370 130.310 145.960 134.100 ;
        RECT 138.080 129.720 145.960 130.310 ;
        RECT 4.100 124.285 135.120 127.485 ;
        RECT 4.100 44.835 4.900 124.285 ;
        RECT 8.665 123.695 70.175 124.285 ;
        RECT 8.665 122.800 10.615 123.695 ;
        RECT 11.335 123.005 13.295 123.235 ;
        RECT 13.625 123.005 15.585 123.235 ;
        RECT 17.255 123.005 19.215 123.305 ;
        RECT 19.545 123.005 21.505 123.305 ;
        RECT 23.175 123.005 25.135 123.305 ;
        RECT 25.465 123.005 27.425 123.305 ;
        RECT 29.095 123.005 31.055 123.305 ;
        RECT 31.385 123.005 33.345 123.305 ;
        RECT 35.015 123.005 36.975 123.305 ;
        RECT 37.305 123.005 39.265 123.305 ;
        RECT 40.935 123.005 42.895 123.305 ;
        RECT 43.225 123.005 45.185 123.305 ;
        RECT 46.855 123.005 48.815 123.305 ;
        RECT 49.145 123.005 51.105 123.305 ;
        RECT 52.775 123.005 54.735 123.305 ;
        RECT 55.065 123.005 57.025 123.305 ;
        RECT 58.695 123.005 60.655 123.305 ;
        RECT 60.985 123.005 62.945 123.305 ;
        RECT 64.615 123.005 66.575 123.235 ;
        RECT 66.905 123.005 68.865 123.235 ;
        RECT 69.585 122.800 70.175 123.695 ;
        RECT 8.665 117.050 11.285 122.800 ;
        RECT 13.345 117.050 13.575 122.800 ;
        RECT 15.635 117.050 15.865 122.800 ;
        RECT 16.975 117.050 17.205 122.800 ;
        RECT 19.265 122.050 19.495 122.800 ;
        RECT 19.030 120.550 19.730 122.050 ;
        RECT 8.665 115.550 11.520 117.050 ;
        RECT 13.110 115.550 13.810 117.050 ;
        RECT 15.400 115.550 16.100 117.050 ;
        RECT 16.740 115.550 17.440 117.050 ;
        RECT 8.665 114.595 11.285 115.550 ;
        RECT 13.345 114.595 13.575 115.550 ;
        RECT 15.635 114.595 15.865 115.550 ;
        RECT 16.975 114.800 17.205 115.550 ;
        RECT 19.265 114.800 19.495 120.550 ;
        RECT 21.555 117.050 21.785 122.800 ;
        RECT 22.895 117.050 23.125 122.800 ;
        RECT 25.185 119.550 25.415 122.800 ;
        RECT 24.950 118.050 25.650 119.550 ;
        RECT 21.320 115.550 22.020 117.050 ;
        RECT 22.660 115.550 23.360 117.050 ;
        RECT 21.555 114.800 21.785 115.550 ;
        RECT 22.895 114.800 23.125 115.550 ;
        RECT 25.185 114.800 25.415 118.050 ;
        RECT 27.475 117.050 27.705 122.800 ;
        RECT 28.815 117.050 29.045 122.800 ;
        RECT 27.240 115.550 27.940 117.050 ;
        RECT 28.580 115.550 29.280 117.050 ;
        RECT 27.475 114.800 27.705 115.550 ;
        RECT 28.815 114.800 29.045 115.550 ;
        RECT 31.105 114.595 31.335 122.800 ;
        RECT 33.395 117.050 33.625 122.800 ;
        RECT 34.735 117.050 34.965 122.800 ;
        RECT 37.025 122.050 37.255 122.800 ;
        RECT 36.790 120.550 37.490 122.050 ;
        RECT 33.160 115.550 33.860 117.050 ;
        RECT 34.500 115.550 35.200 117.050 ;
        RECT 33.395 114.800 33.625 115.550 ;
        RECT 34.735 114.800 34.965 115.550 ;
        RECT 37.025 114.800 37.255 120.550 ;
        RECT 39.315 117.050 39.545 122.800 ;
        RECT 40.655 117.050 40.885 122.800 ;
        RECT 42.945 122.050 43.175 122.800 ;
        RECT 42.710 120.550 43.410 122.050 ;
        RECT 39.080 115.550 39.780 117.050 ;
        RECT 40.420 115.550 41.120 117.050 ;
        RECT 39.315 114.800 39.545 115.550 ;
        RECT 40.655 114.800 40.885 115.550 ;
        RECT 42.945 114.800 43.175 120.550 ;
        RECT 45.235 117.050 45.465 122.800 ;
        RECT 46.575 117.050 46.805 122.800 ;
        RECT 45.000 115.550 45.700 117.050 ;
        RECT 46.340 115.550 47.040 117.050 ;
        RECT 45.235 114.800 45.465 115.550 ;
        RECT 46.575 114.800 46.805 115.550 ;
        RECT 48.865 114.595 49.095 122.800 ;
        RECT 51.155 117.050 51.385 122.800 ;
        RECT 52.495 117.050 52.725 122.800 ;
        RECT 54.785 119.550 55.015 122.800 ;
        RECT 54.550 118.050 55.250 119.550 ;
        RECT 50.920 115.550 51.620 117.050 ;
        RECT 52.260 115.550 52.960 117.050 ;
        RECT 51.155 114.800 51.385 115.550 ;
        RECT 52.495 114.800 52.725 115.550 ;
        RECT 54.785 114.800 55.015 118.050 ;
        RECT 57.075 117.050 57.305 122.800 ;
        RECT 58.415 117.050 58.645 122.800 ;
        RECT 60.705 122.050 60.935 122.800 ;
        RECT 60.470 120.550 61.170 122.050 ;
        RECT 56.840 115.550 57.540 117.050 ;
        RECT 58.180 115.550 58.880 117.050 ;
        RECT 57.075 114.800 57.305 115.550 ;
        RECT 58.415 114.800 58.645 115.550 ;
        RECT 60.705 114.800 60.935 120.550 ;
        RECT 62.995 117.050 63.225 122.800 ;
        RECT 64.335 117.050 64.565 122.800 ;
        RECT 66.625 117.050 66.855 122.800 ;
        RECT 68.915 117.050 70.175 122.800 ;
        RECT 62.760 115.550 63.460 117.050 ;
        RECT 64.100 115.550 64.800 117.050 ;
        RECT 66.390 115.550 67.090 117.050 ;
        RECT 68.680 115.550 70.175 117.050 ;
        RECT 62.995 114.800 63.225 115.550 ;
        RECT 64.335 114.595 64.565 115.550 ;
        RECT 66.625 114.595 66.855 115.550 ;
        RECT 68.915 114.595 70.175 115.550 ;
        RECT 8.665 114.365 15.865 114.595 ;
        RECT 8.665 113.215 10.615 114.365 ;
        RECT 17.255 114.295 19.215 114.595 ;
        RECT 19.545 114.295 21.505 114.595 ;
        RECT 23.175 114.295 25.135 114.595 ;
        RECT 25.465 114.295 27.425 114.595 ;
        RECT 29.095 114.365 33.345 114.595 ;
        RECT 29.095 114.295 31.055 114.365 ;
        RECT 31.385 114.295 33.345 114.365 ;
        RECT 35.015 114.295 36.975 114.595 ;
        RECT 37.305 114.295 39.265 114.595 ;
        RECT 40.935 114.295 42.895 114.595 ;
        RECT 43.225 114.295 45.185 114.595 ;
        RECT 46.855 114.365 51.105 114.595 ;
        RECT 46.855 114.295 48.815 114.365 ;
        RECT 49.145 114.295 51.105 114.365 ;
        RECT 52.775 114.295 54.735 114.595 ;
        RECT 55.065 114.295 57.025 114.595 ;
        RECT 58.695 114.295 60.655 114.595 ;
        RECT 60.985 114.295 62.945 114.595 ;
        RECT 64.335 114.365 70.175 114.595 ;
        RECT 8.665 112.985 15.865 113.215 ;
        RECT 17.255 112.985 19.215 113.285 ;
        RECT 19.545 112.985 21.505 113.285 ;
        RECT 23.175 112.985 25.135 113.285 ;
        RECT 25.465 112.985 27.425 113.285 ;
        RECT 29.095 113.215 31.055 113.285 ;
        RECT 31.385 113.215 33.345 113.285 ;
        RECT 29.095 112.985 33.345 113.215 ;
        RECT 35.015 112.985 36.975 113.285 ;
        RECT 37.305 112.985 39.265 113.285 ;
        RECT 40.935 112.985 42.895 113.285 ;
        RECT 43.225 112.985 45.185 113.285 ;
        RECT 46.855 113.215 48.815 113.285 ;
        RECT 49.145 113.215 51.105 113.285 ;
        RECT 46.855 112.985 51.105 113.215 ;
        RECT 52.775 112.985 54.735 113.285 ;
        RECT 55.065 112.985 57.025 113.285 ;
        RECT 58.695 112.985 60.655 113.285 ;
        RECT 60.985 112.985 62.945 113.285 ;
        RECT 69.585 113.215 70.175 114.365 ;
        RECT 64.335 112.985 70.175 113.215 ;
        RECT 8.665 112.030 11.285 112.985 ;
        RECT 13.345 112.030 13.575 112.985 ;
        RECT 15.635 112.030 15.865 112.985 ;
        RECT 16.975 112.030 17.205 112.780 ;
        RECT 8.665 110.530 11.520 112.030 ;
        RECT 13.110 110.530 13.810 112.030 ;
        RECT 15.400 110.530 16.100 112.030 ;
        RECT 16.740 110.530 17.440 112.030 ;
        RECT 8.665 104.780 11.285 110.530 ;
        RECT 13.345 104.780 13.575 110.530 ;
        RECT 15.635 104.780 15.865 110.530 ;
        RECT 16.975 104.780 17.205 110.530 ;
        RECT 19.265 107.030 19.495 112.780 ;
        RECT 21.555 112.030 21.785 112.780 ;
        RECT 22.895 112.030 23.125 112.780 ;
        RECT 21.320 110.530 22.020 112.030 ;
        RECT 22.660 110.530 23.360 112.030 ;
        RECT 19.030 105.530 19.730 107.030 ;
        RECT 19.265 104.780 19.495 105.530 ;
        RECT 21.555 104.780 21.785 110.530 ;
        RECT 22.895 104.780 23.125 110.530 ;
        RECT 25.185 109.530 25.415 112.780 ;
        RECT 27.475 112.030 27.705 112.780 ;
        RECT 28.815 112.030 29.045 112.780 ;
        RECT 27.240 110.530 27.940 112.030 ;
        RECT 28.580 110.530 29.280 112.030 ;
        RECT 24.950 108.030 25.650 109.530 ;
        RECT 25.185 104.780 25.415 108.030 ;
        RECT 27.475 104.780 27.705 110.530 ;
        RECT 28.815 104.780 29.045 110.530 ;
        RECT 31.105 104.780 31.335 112.985 ;
        RECT 33.395 112.030 33.625 112.780 ;
        RECT 34.735 112.030 34.965 112.780 ;
        RECT 33.160 110.530 33.860 112.030 ;
        RECT 34.500 110.530 35.200 112.030 ;
        RECT 33.395 104.780 33.625 110.530 ;
        RECT 34.735 104.780 34.965 110.530 ;
        RECT 37.025 107.030 37.255 112.780 ;
        RECT 39.315 112.030 39.545 112.780 ;
        RECT 40.655 112.030 40.885 112.780 ;
        RECT 39.080 110.530 39.780 112.030 ;
        RECT 40.420 110.530 41.120 112.030 ;
        RECT 36.790 105.530 37.490 107.030 ;
        RECT 37.025 104.780 37.255 105.530 ;
        RECT 39.315 104.780 39.545 110.530 ;
        RECT 40.655 104.780 40.885 110.530 ;
        RECT 42.945 107.030 43.175 112.780 ;
        RECT 45.235 112.030 45.465 112.780 ;
        RECT 46.575 112.030 46.805 112.780 ;
        RECT 45.000 110.530 45.700 112.030 ;
        RECT 46.340 110.530 47.040 112.030 ;
        RECT 42.710 105.530 43.410 107.030 ;
        RECT 42.945 104.780 43.175 105.530 ;
        RECT 45.235 104.780 45.465 110.530 ;
        RECT 46.575 104.780 46.805 110.530 ;
        RECT 48.865 104.780 49.095 112.985 ;
        RECT 51.155 112.030 51.385 112.780 ;
        RECT 52.495 112.030 52.725 112.780 ;
        RECT 50.920 110.530 51.620 112.030 ;
        RECT 52.260 110.530 52.960 112.030 ;
        RECT 51.155 104.780 51.385 110.530 ;
        RECT 52.495 104.780 52.725 110.530 ;
        RECT 54.785 109.530 55.015 112.780 ;
        RECT 57.075 112.030 57.305 112.780 ;
        RECT 58.415 112.030 58.645 112.780 ;
        RECT 56.840 110.530 57.540 112.030 ;
        RECT 58.180 110.530 58.880 112.030 ;
        RECT 54.550 108.030 55.250 109.530 ;
        RECT 54.785 104.780 55.015 108.030 ;
        RECT 57.075 104.780 57.305 110.530 ;
        RECT 58.415 104.780 58.645 110.530 ;
        RECT 60.705 107.030 60.935 112.780 ;
        RECT 62.995 112.030 63.225 112.780 ;
        RECT 64.335 112.030 64.565 112.985 ;
        RECT 66.625 112.030 66.855 112.985 ;
        RECT 68.915 112.030 70.175 112.985 ;
        RECT 62.760 110.530 63.460 112.030 ;
        RECT 64.100 110.530 64.800 112.030 ;
        RECT 66.390 110.530 67.090 112.030 ;
        RECT 68.680 110.530 70.175 112.030 ;
        RECT 60.470 105.530 61.170 107.030 ;
        RECT 60.705 104.780 60.935 105.530 ;
        RECT 62.995 104.780 63.225 110.530 ;
        RECT 64.335 104.780 64.565 110.530 ;
        RECT 66.625 104.780 66.855 110.530 ;
        RECT 68.915 104.780 70.175 110.530 ;
        RECT 8.665 103.885 10.615 104.780 ;
        RECT 11.335 104.345 13.295 104.575 ;
        RECT 13.625 104.345 15.585 104.575 ;
        RECT 17.255 104.275 19.215 104.575 ;
        RECT 19.545 104.275 21.505 104.575 ;
        RECT 23.175 104.275 25.135 104.575 ;
        RECT 25.465 104.275 27.425 104.575 ;
        RECT 29.095 104.275 31.055 104.575 ;
        RECT 31.385 104.275 33.345 104.575 ;
        RECT 35.015 104.275 36.975 104.575 ;
        RECT 37.305 104.275 39.265 104.575 ;
        RECT 40.935 104.275 42.895 104.575 ;
        RECT 43.225 104.275 45.185 104.575 ;
        RECT 46.855 104.275 48.815 104.575 ;
        RECT 49.145 104.275 51.105 104.575 ;
        RECT 52.775 104.275 54.735 104.575 ;
        RECT 55.065 104.275 57.025 104.575 ;
        RECT 58.695 104.275 60.655 104.575 ;
        RECT 60.985 104.275 62.945 104.575 ;
        RECT 64.615 104.345 66.575 104.575 ;
        RECT 66.905 104.345 68.865 104.575 ;
        RECT 69.585 103.885 70.175 104.780 ;
        RECT 8.665 102.705 70.175 103.885 ;
        RECT 71.775 123.695 114.165 124.285 ;
        RECT 71.775 103.885 72.365 123.695 ;
        RECT 72.805 122.800 77.615 123.695 ;
        RECT 79.005 123.005 80.965 123.305 ;
        RECT 81.295 123.005 83.255 123.305 ;
        RECT 84.925 123.005 86.885 123.305 ;
        RECT 87.215 123.005 89.175 123.305 ;
        RECT 90.845 123.005 95.095 123.305 ;
        RECT 96.765 123.005 98.725 123.305 ;
        RECT 99.055 123.005 101.015 123.305 ;
        RECT 102.685 123.005 104.645 123.305 ;
        RECT 104.975 123.005 106.935 123.305 ;
        RECT 72.805 114.800 73.035 122.800 ;
        RECT 75.095 114.800 75.325 122.800 ;
        RECT 77.385 114.800 77.615 122.800 ;
        RECT 78.725 120.650 78.955 122.800 ;
        RECT 78.490 119.950 79.190 120.650 ;
        RECT 78.725 114.800 78.955 119.950 ;
        RECT 81.015 119.150 81.245 122.800 ;
        RECT 83.305 120.650 83.535 122.800 ;
        RECT 83.070 119.950 83.770 120.650 ;
        RECT 80.780 118.450 81.480 119.150 ;
        RECT 81.015 114.800 81.245 118.450 ;
        RECT 83.305 114.800 83.535 119.950 ;
        RECT 84.645 116.150 84.875 122.800 ;
        RECT 86.935 117.650 87.165 122.800 ;
        RECT 86.700 116.950 87.400 117.650 ;
        RECT 84.410 115.450 85.110 116.150 ;
        RECT 84.645 114.800 84.875 115.450 ;
        RECT 86.935 114.800 87.165 116.950 ;
        RECT 89.225 116.150 89.455 122.800 ;
        RECT 90.565 122.150 90.795 122.800 ;
        RECT 90.330 121.450 91.030 122.150 ;
        RECT 88.990 115.450 89.690 116.150 ;
        RECT 89.225 114.800 89.455 115.450 ;
        RECT 90.565 114.800 90.795 121.450 ;
        RECT 92.855 114.800 93.085 123.005 ;
        RECT 108.325 122.800 113.135 123.695 ;
        RECT 95.145 122.150 95.375 122.800 ;
        RECT 94.910 121.450 95.610 122.150 ;
        RECT 95.145 114.800 95.375 121.450 ;
        RECT 96.485 116.150 96.715 122.800 ;
        RECT 98.775 117.650 99.005 122.800 ;
        RECT 98.540 116.950 99.240 117.650 ;
        RECT 96.250 115.450 96.950 116.150 ;
        RECT 96.485 114.800 96.715 115.450 ;
        RECT 98.775 114.800 99.005 116.950 ;
        RECT 101.065 116.150 101.295 122.800 ;
        RECT 102.405 120.650 102.635 122.800 ;
        RECT 102.170 119.950 102.870 120.650 ;
        RECT 100.830 115.450 101.530 116.150 ;
        RECT 101.065 114.800 101.295 115.450 ;
        RECT 102.405 114.800 102.635 119.950 ;
        RECT 104.695 119.150 104.925 122.800 ;
        RECT 106.985 120.650 107.215 122.800 ;
        RECT 106.750 119.950 107.450 120.650 ;
        RECT 104.460 118.450 105.160 119.150 ;
        RECT 104.695 114.800 104.925 118.450 ;
        RECT 106.985 114.800 107.215 119.950 ;
        RECT 108.325 114.800 108.555 122.800 ;
        RECT 110.615 114.800 110.845 122.800 ;
        RECT 112.905 114.800 113.135 122.800 ;
        RECT 73.085 114.365 75.045 114.595 ;
        RECT 75.375 114.365 77.335 114.595 ;
        RECT 79.005 114.295 80.965 114.595 ;
        RECT 81.295 114.295 83.255 114.595 ;
        RECT 84.925 114.295 86.885 114.595 ;
        RECT 87.215 114.295 89.175 114.595 ;
        RECT 90.845 114.295 92.805 114.595 ;
        RECT 93.135 114.295 95.095 114.595 ;
        RECT 96.765 114.295 98.725 114.595 ;
        RECT 99.055 114.295 101.015 114.595 ;
        RECT 102.685 114.295 104.645 114.595 ;
        RECT 104.975 114.295 106.935 114.595 ;
        RECT 108.605 114.365 110.565 114.595 ;
        RECT 110.895 114.365 112.855 114.595 ;
        RECT 73.085 112.985 75.045 113.215 ;
        RECT 75.375 112.985 77.335 113.215 ;
        RECT 79.005 112.985 80.965 113.285 ;
        RECT 81.295 112.985 83.255 113.285 ;
        RECT 84.925 112.985 86.885 113.285 ;
        RECT 87.215 112.985 89.175 113.285 ;
        RECT 90.845 112.985 92.805 113.285 ;
        RECT 93.135 112.985 95.095 113.285 ;
        RECT 96.765 112.985 98.725 113.285 ;
        RECT 99.055 112.985 101.015 113.285 ;
        RECT 102.685 112.985 104.645 113.285 ;
        RECT 104.975 112.985 106.935 113.285 ;
        RECT 108.605 112.985 110.565 113.215 ;
        RECT 110.895 112.985 112.855 113.215 ;
        RECT 72.805 104.780 73.035 112.780 ;
        RECT 75.095 104.780 75.325 112.780 ;
        RECT 77.385 104.780 77.615 112.780 ;
        RECT 78.725 107.630 78.955 112.780 ;
        RECT 81.015 109.130 81.245 112.780 ;
        RECT 80.780 108.430 81.480 109.130 ;
        RECT 78.490 106.930 79.190 107.630 ;
        RECT 78.725 104.780 78.955 106.930 ;
        RECT 81.015 104.780 81.245 108.430 ;
        RECT 83.305 107.630 83.535 112.780 ;
        RECT 84.645 112.130 84.875 112.780 ;
        RECT 84.410 111.430 85.110 112.130 ;
        RECT 83.070 106.930 83.770 107.630 ;
        RECT 83.305 104.780 83.535 106.930 ;
        RECT 84.645 104.780 84.875 111.430 ;
        RECT 86.935 110.630 87.165 112.780 ;
        RECT 89.225 112.130 89.455 112.780 ;
        RECT 88.990 111.430 89.690 112.130 ;
        RECT 86.700 109.930 87.400 110.630 ;
        RECT 86.935 104.780 87.165 109.930 ;
        RECT 89.225 104.780 89.455 111.430 ;
        RECT 90.565 106.130 90.795 112.780 ;
        RECT 90.330 105.430 91.030 106.130 ;
        RECT 90.565 104.780 90.795 105.430 ;
        RECT 72.805 103.885 77.615 104.780 ;
        RECT 92.855 104.575 93.085 112.780 ;
        RECT 95.145 106.130 95.375 112.780 ;
        RECT 96.485 112.130 96.715 112.780 ;
        RECT 96.250 111.430 96.950 112.130 ;
        RECT 94.910 105.430 95.610 106.130 ;
        RECT 95.145 104.780 95.375 105.430 ;
        RECT 96.485 104.780 96.715 111.430 ;
        RECT 98.775 110.630 99.005 112.780 ;
        RECT 101.065 112.130 101.295 112.780 ;
        RECT 100.830 111.430 101.530 112.130 ;
        RECT 98.540 109.930 99.240 110.630 ;
        RECT 98.775 104.780 99.005 109.930 ;
        RECT 101.065 104.780 101.295 111.430 ;
        RECT 102.405 107.630 102.635 112.780 ;
        RECT 104.695 109.130 104.925 112.780 ;
        RECT 104.460 108.430 105.160 109.130 ;
        RECT 102.170 106.930 102.870 107.630 ;
        RECT 102.405 104.780 102.635 106.930 ;
        RECT 104.695 104.780 104.925 108.430 ;
        RECT 106.985 107.630 107.215 112.780 ;
        RECT 106.750 106.930 107.450 107.630 ;
        RECT 106.985 104.780 107.215 106.930 ;
        RECT 108.325 104.780 108.555 112.780 ;
        RECT 110.615 104.780 110.845 112.780 ;
        RECT 112.905 104.780 113.135 112.780 ;
        RECT 79.005 104.275 80.965 104.575 ;
        RECT 81.295 104.275 83.255 104.575 ;
        RECT 84.925 104.275 86.885 104.575 ;
        RECT 87.215 104.275 89.175 104.575 ;
        RECT 90.845 104.275 95.095 104.575 ;
        RECT 96.765 104.275 98.725 104.575 ;
        RECT 99.055 104.275 101.015 104.575 ;
        RECT 102.685 104.275 104.645 104.575 ;
        RECT 104.975 104.275 106.935 104.575 ;
        RECT 108.325 103.885 113.135 104.780 ;
        RECT 113.575 103.885 114.165 123.695 ;
        RECT 128.935 123.505 135.120 124.285 ;
        RECT 138.080 128.380 145.960 128.970 ;
        RECT 138.080 124.680 138.670 128.380 ;
        RECT 139.205 127.290 139.435 127.530 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.205 125.530 139.435 125.690 ;
        RECT 140.495 125.530 140.725 128.380 ;
        RECT 143.725 127.920 144.425 127.990 ;
        RECT 143.595 127.690 144.555 127.920 ;
        RECT 141.785 127.290 142.015 127.530 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 143.315 126.865 143.545 127.530 ;
        RECT 143.280 126.165 143.580 126.865 ;
        RECT 141.785 125.530 142.015 125.690 ;
        RECT 143.315 125.370 143.545 126.165 ;
        RECT 139.390 125.140 143.545 125.370 ;
        RECT 144.605 124.680 144.835 127.530 ;
        RECT 145.370 124.680 145.960 128.380 ;
        RECT 138.080 124.090 145.960 124.680 ;
        RECT 71.775 102.705 114.165 103.885 ;
        RECT 115.905 122.915 135.120 123.505 ;
        RECT 115.905 122.475 116.495 122.915 ;
        RECT 115.905 122.245 118.390 122.475 ;
        RECT 115.905 114.185 117.185 122.245 ;
        RECT 118.595 114.235 118.825 122.195 ;
        RECT 119.975 118.645 120.205 122.195 ;
        RECT 120.410 122.010 121.410 122.710 ;
        RECT 121.615 118.645 121.845 122.195 ;
        RECT 119.975 117.075 121.845 118.645 ;
        RECT 115.905 113.955 118.390 114.185 ;
        RECT 115.905 112.845 116.495 113.955 ;
        RECT 115.905 112.615 118.390 112.845 ;
        RECT 115.905 104.555 117.185 112.615 ;
        RECT 118.595 104.605 118.825 112.565 ;
        RECT 119.975 109.685 120.205 117.075 ;
        RECT 121.615 114.235 121.845 117.075 ;
        RECT 122.995 118.645 123.225 122.195 ;
        RECT 123.430 122.010 124.430 122.710 ;
        RECT 128.345 122.475 135.120 122.915 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 126.450 122.245 135.120 122.475 ;
        RECT 124.635 118.645 124.865 122.195 ;
        RECT 122.995 117.075 124.865 118.645 ;
        RECT 122.995 114.235 123.225 117.075 ;
        RECT 120.410 112.615 121.410 114.185 ;
        RECT 123.430 112.615 124.430 114.185 ;
        RECT 121.615 109.685 121.845 112.565 ;
        RECT 119.975 108.115 121.845 109.685 ;
        RECT 119.975 104.605 120.205 108.115 ;
        RECT 115.905 104.325 118.390 104.555 ;
        RECT 115.905 103.885 116.495 104.325 ;
        RECT 120.410 104.090 121.410 104.790 ;
        RECT 121.615 104.605 121.845 108.115 ;
        RECT 122.995 109.685 123.225 112.565 ;
        RECT 124.635 109.685 124.865 117.075 ;
        RECT 126.015 114.235 126.245 122.195 ;
        RECT 127.655 114.185 135.120 122.245 ;
        RECT 126.450 113.955 135.120 114.185 ;
        RECT 128.345 112.845 135.120 113.955 ;
        RECT 126.450 112.615 135.120 112.845 ;
        RECT 122.995 108.115 124.865 109.685 ;
        RECT 122.995 104.605 123.225 108.115 ;
        RECT 123.430 104.090 124.430 104.790 ;
        RECT 124.635 104.605 124.865 108.115 ;
        RECT 126.015 104.605 126.245 112.565 ;
        RECT 127.655 107.765 135.120 112.615 ;
        RECT 136.295 108.925 142.995 109.515 ;
        RECT 127.655 104.835 138.400 107.765 ;
        RECT 127.655 104.555 135.710 104.835 ;
        RECT 126.450 104.325 135.710 104.555 ;
        RECT 128.345 103.885 135.710 104.325 ;
        RECT 115.905 102.705 135.710 103.885 ;
        RECT 8.665 102.115 135.710 102.705 ;
        RECT 136.295 102.495 138.400 104.255 ;
        RECT 8.665 44.835 10.615 102.115 ;
        RECT 4.100 42.225 10.615 44.835 ;
        RECT 11.055 101.425 29.605 102.115 ;
        RECT 11.055 93.015 11.285 101.425 ;
        RECT 13.345 93.015 13.575 101.425 ;
        RECT 15.635 93.015 15.865 101.425 ;
        RECT 17.925 93.015 18.155 101.425 ;
        RECT 20.215 93.015 20.445 101.425 ;
        RECT 22.505 93.015 22.735 101.425 ;
        RECT 24.795 93.015 25.025 101.425 ;
        RECT 27.085 93.015 27.315 101.425 ;
        RECT 29.375 93.015 29.605 101.425 ;
        RECT 30.715 101.425 49.265 102.115 ;
        RECT 30.715 93.220 30.945 101.425 ;
        RECT 33.005 93.220 33.235 101.425 ;
        RECT 35.295 93.220 35.525 101.425 ;
        RECT 37.585 93.220 37.815 101.425 ;
        RECT 39.875 93.220 40.105 101.425 ;
        RECT 42.165 93.220 42.395 101.425 ;
        RECT 44.455 93.220 44.685 101.425 ;
        RECT 46.745 93.220 46.975 101.425 ;
        RECT 49.035 93.220 49.265 101.425 ;
        RECT 50.375 101.425 68.925 102.115 ;
        RECT 50.375 93.220 50.605 101.425 ;
        RECT 52.665 93.220 52.895 101.425 ;
        RECT 54.955 93.220 55.185 101.425 ;
        RECT 57.245 93.220 57.475 101.425 ;
        RECT 59.535 93.220 59.765 101.425 ;
        RECT 61.825 93.220 62.055 101.425 ;
        RECT 64.115 93.220 64.345 101.425 ;
        RECT 66.405 93.220 66.635 101.425 ;
        RECT 68.695 93.220 68.925 101.425 ;
        RECT 70.035 101.425 88.585 102.115 ;
        RECT 70.035 93.220 70.265 101.425 ;
        RECT 72.325 93.220 72.555 101.425 ;
        RECT 74.615 93.220 74.845 101.425 ;
        RECT 76.905 93.220 77.135 101.425 ;
        RECT 79.195 93.220 79.425 101.425 ;
        RECT 81.485 93.220 81.715 101.425 ;
        RECT 83.775 93.220 84.005 101.425 ;
        RECT 86.065 93.220 86.295 101.425 ;
        RECT 88.355 93.220 88.585 101.425 ;
        RECT 89.695 101.425 108.245 102.115 ;
        RECT 89.695 93.220 89.925 101.425 ;
        RECT 91.985 93.220 92.215 101.425 ;
        RECT 94.275 93.220 94.505 101.425 ;
        RECT 96.565 93.220 96.795 101.425 ;
        RECT 98.855 93.220 99.085 101.425 ;
        RECT 101.145 93.220 101.375 101.425 ;
        RECT 103.435 93.220 103.665 101.425 ;
        RECT 105.725 93.220 105.955 101.425 ;
        RECT 108.015 93.220 108.245 101.425 ;
        RECT 109.355 101.425 127.905 102.115 ;
        RECT 109.355 93.015 109.585 101.425 ;
        RECT 111.645 93.015 111.875 101.425 ;
        RECT 113.935 93.015 114.165 101.425 ;
        RECT 116.225 93.015 116.455 101.425 ;
        RECT 118.515 93.015 118.745 101.425 ;
        RECT 120.805 93.015 121.035 101.425 ;
        RECT 123.095 93.015 123.325 101.425 ;
        RECT 125.385 93.015 125.615 101.425 ;
        RECT 127.675 93.015 127.905 101.425 ;
        RECT 11.055 91.405 29.605 93.015 ;
        RECT 30.995 92.785 32.955 93.015 ;
        RECT 33.285 92.785 35.245 93.015 ;
        RECT 35.575 92.785 37.535 93.015 ;
        RECT 37.865 92.785 39.825 93.015 ;
        RECT 40.155 92.785 42.115 93.015 ;
        RECT 42.445 92.785 44.405 93.015 ;
        RECT 44.735 92.785 46.695 93.015 ;
        RECT 47.025 92.785 48.985 93.015 ;
        RECT 50.655 92.785 52.615 93.015 ;
        RECT 52.945 92.785 54.905 93.015 ;
        RECT 55.235 92.785 57.195 93.015 ;
        RECT 57.525 92.785 59.485 93.015 ;
        RECT 59.815 92.785 61.775 93.015 ;
        RECT 62.105 92.785 64.065 93.015 ;
        RECT 64.395 92.785 66.355 93.015 ;
        RECT 66.685 92.785 68.645 93.015 ;
        RECT 70.315 92.785 72.275 93.015 ;
        RECT 72.605 92.785 74.565 93.015 ;
        RECT 74.895 92.785 76.855 93.015 ;
        RECT 77.185 92.785 79.145 93.015 ;
        RECT 79.475 92.785 81.435 93.015 ;
        RECT 81.765 92.785 83.725 93.015 ;
        RECT 84.055 92.785 86.015 93.015 ;
        RECT 86.345 92.785 88.305 93.015 ;
        RECT 89.975 92.785 91.935 93.015 ;
        RECT 92.265 92.785 94.225 93.015 ;
        RECT 94.555 92.785 96.515 93.015 ;
        RECT 96.845 92.785 98.805 93.015 ;
        RECT 99.135 92.785 101.095 93.015 ;
        RECT 101.425 92.785 103.385 93.015 ;
        RECT 103.715 92.785 105.675 93.015 ;
        RECT 106.005 92.785 107.965 93.015 ;
        RECT 30.995 91.405 32.955 91.635 ;
        RECT 11.055 82.995 11.285 91.405 ;
        RECT 13.345 82.995 13.575 91.405 ;
        RECT 15.635 82.995 15.865 91.405 ;
        RECT 17.925 82.995 18.155 91.405 ;
        RECT 20.215 82.995 20.445 91.405 ;
        RECT 22.505 82.995 22.735 91.405 ;
        RECT 24.795 82.995 25.025 91.405 ;
        RECT 27.085 82.995 27.315 91.405 ;
        RECT 29.375 82.995 29.605 91.405 ;
        RECT 33.285 91.345 35.245 91.875 ;
        RECT 35.575 91.345 37.535 91.875 ;
        RECT 37.865 91.405 39.825 91.635 ;
        RECT 40.155 91.405 42.115 91.635 ;
        RECT 42.445 91.345 44.405 91.875 ;
        RECT 44.735 91.345 46.695 91.875 ;
        RECT 47.025 91.405 48.985 91.635 ;
        RECT 50.655 91.345 52.615 91.875 ;
        RECT 52.945 91.405 54.905 91.635 ;
        RECT 55.235 91.405 57.195 91.635 ;
        RECT 57.525 91.345 59.485 91.875 ;
        RECT 59.815 91.345 61.775 91.875 ;
        RECT 62.105 91.405 64.065 91.635 ;
        RECT 64.395 91.405 66.355 91.635 ;
        RECT 66.685 91.345 68.645 91.875 ;
        RECT 70.315 91.345 72.275 91.875 ;
        RECT 72.605 91.405 74.565 91.635 ;
        RECT 74.895 91.405 76.855 91.635 ;
        RECT 77.185 91.345 79.145 91.875 ;
        RECT 79.475 91.345 81.435 91.875 ;
        RECT 81.765 91.405 83.725 91.635 ;
        RECT 84.055 91.405 86.015 91.635 ;
        RECT 86.345 91.345 88.305 91.875 ;
        RECT 89.975 91.405 91.935 91.635 ;
        RECT 92.265 91.345 94.225 91.875 ;
        RECT 94.555 91.345 96.515 91.875 ;
        RECT 96.845 91.405 98.805 91.635 ;
        RECT 99.135 91.405 101.095 91.635 ;
        RECT 101.425 91.345 103.385 91.875 ;
        RECT 103.715 91.345 105.675 91.875 ;
        RECT 106.005 91.405 107.965 91.635 ;
        RECT 109.355 91.405 127.905 93.015 ;
        RECT 30.715 84.590 30.945 91.200 ;
        RECT 33.005 88.540 33.235 91.200 ;
        RECT 35.295 91.090 35.525 91.200 ;
        RECT 35.260 89.690 35.560 91.090 ;
        RECT 32.970 85.740 33.270 88.540 ;
        RECT 30.680 83.190 30.980 84.590 ;
        RECT 33.005 83.200 33.235 85.740 ;
        RECT 35.295 83.200 35.525 89.690 ;
        RECT 37.585 88.540 37.815 91.200 ;
        RECT 37.550 85.740 37.850 88.540 ;
        RECT 37.585 83.200 37.815 85.740 ;
        RECT 39.875 84.590 40.105 91.200 ;
        RECT 42.165 88.540 42.395 91.200 ;
        RECT 44.455 91.090 44.685 91.200 ;
        RECT 44.420 89.690 44.720 91.090 ;
        RECT 42.130 85.740 42.430 88.540 ;
        RECT 39.840 83.190 40.140 84.590 ;
        RECT 42.165 83.200 42.395 85.740 ;
        RECT 44.455 83.200 44.685 89.690 ;
        RECT 46.745 88.540 46.975 91.200 ;
        RECT 46.710 85.740 47.010 88.540 ;
        RECT 46.745 83.200 46.975 85.740 ;
        RECT 49.035 84.590 49.265 91.200 ;
        RECT 50.375 91.090 50.605 91.200 ;
        RECT 50.340 89.690 50.640 91.090 ;
        RECT 49.000 83.190 49.300 84.590 ;
        RECT 50.375 83.200 50.605 89.690 ;
        RECT 52.665 88.540 52.895 91.200 ;
        RECT 52.630 85.740 52.930 88.540 ;
        RECT 52.665 83.200 52.895 85.740 ;
        RECT 54.955 84.590 55.185 91.200 ;
        RECT 57.245 88.540 57.475 91.200 ;
        RECT 59.535 91.090 59.765 91.200 ;
        RECT 59.500 89.690 59.800 91.090 ;
        RECT 57.210 85.740 57.510 88.540 ;
        RECT 54.920 83.190 55.220 84.590 ;
        RECT 57.245 83.200 57.475 85.740 ;
        RECT 59.535 83.200 59.765 89.690 ;
        RECT 61.825 88.540 62.055 91.200 ;
        RECT 61.790 85.740 62.090 88.540 ;
        RECT 61.825 83.200 62.055 85.740 ;
        RECT 64.115 84.590 64.345 91.200 ;
        RECT 66.405 88.540 66.635 91.200 ;
        RECT 68.695 91.090 68.925 91.200 ;
        RECT 70.035 91.090 70.265 91.200 ;
        RECT 68.660 89.690 68.960 91.090 ;
        RECT 70.000 89.690 70.300 91.090 ;
        RECT 66.370 85.740 66.670 88.540 ;
        RECT 64.080 83.190 64.380 84.590 ;
        RECT 66.405 83.200 66.635 85.740 ;
        RECT 68.695 83.200 68.925 89.690 ;
        RECT 70.035 83.200 70.265 89.690 ;
        RECT 72.325 88.540 72.555 91.200 ;
        RECT 72.290 85.740 72.590 88.540 ;
        RECT 72.325 83.200 72.555 85.740 ;
        RECT 74.615 84.590 74.845 91.200 ;
        RECT 76.905 88.540 77.135 91.200 ;
        RECT 79.195 91.090 79.425 91.200 ;
        RECT 79.160 89.690 79.460 91.090 ;
        RECT 76.870 85.740 77.170 88.540 ;
        RECT 74.580 83.190 74.880 84.590 ;
        RECT 76.905 83.200 77.135 85.740 ;
        RECT 79.195 83.200 79.425 89.690 ;
        RECT 81.485 88.540 81.715 91.200 ;
        RECT 81.450 85.740 81.750 88.540 ;
        RECT 81.485 83.200 81.715 85.740 ;
        RECT 83.775 84.590 84.005 91.200 ;
        RECT 86.065 88.540 86.295 91.200 ;
        RECT 88.355 91.090 88.585 91.200 ;
        RECT 88.320 89.690 88.620 91.090 ;
        RECT 86.030 85.740 86.330 88.540 ;
        RECT 83.740 83.190 84.040 84.590 ;
        RECT 86.065 83.200 86.295 85.740 ;
        RECT 88.355 83.200 88.585 89.690 ;
        RECT 89.695 84.590 89.925 91.200 ;
        RECT 91.985 88.540 92.215 91.200 ;
        RECT 94.275 91.090 94.505 91.200 ;
        RECT 94.240 89.690 94.540 91.090 ;
        RECT 91.950 85.740 92.250 88.540 ;
        RECT 89.660 83.190 89.960 84.590 ;
        RECT 91.985 83.200 92.215 85.740 ;
        RECT 94.275 83.200 94.505 89.690 ;
        RECT 96.565 88.540 96.795 91.200 ;
        RECT 96.530 85.740 96.830 88.540 ;
        RECT 96.565 83.200 96.795 85.740 ;
        RECT 98.855 84.590 99.085 91.200 ;
        RECT 101.145 88.540 101.375 91.200 ;
        RECT 103.435 91.090 103.665 91.200 ;
        RECT 103.400 89.690 103.700 91.090 ;
        RECT 101.110 85.740 101.410 88.540 ;
        RECT 98.820 83.190 99.120 84.590 ;
        RECT 101.145 83.200 101.375 85.740 ;
        RECT 103.435 83.200 103.665 89.690 ;
        RECT 105.725 88.540 105.955 91.200 ;
        RECT 105.690 85.740 105.990 88.540 ;
        RECT 105.725 83.200 105.955 85.740 ;
        RECT 108.015 84.590 108.245 91.200 ;
        RECT 107.980 83.190 108.280 84.590 ;
        RECT 109.355 82.995 109.585 91.405 ;
        RECT 111.645 82.995 111.875 91.405 ;
        RECT 113.935 82.995 114.165 91.405 ;
        RECT 116.225 82.995 116.455 91.405 ;
        RECT 118.515 82.995 118.745 91.405 ;
        RECT 120.805 82.995 121.035 91.405 ;
        RECT 123.095 82.995 123.325 91.405 ;
        RECT 125.385 82.995 125.615 91.405 ;
        RECT 127.675 82.995 127.905 91.405 ;
        RECT 11.055 81.385 29.605 82.995 ;
        RECT 30.995 82.405 32.955 82.995 ;
        RECT 33.285 82.765 35.245 82.995 ;
        RECT 35.575 82.765 37.535 82.995 ;
        RECT 37.865 82.405 39.825 82.995 ;
        RECT 40.155 82.405 42.115 82.995 ;
        RECT 42.445 82.765 44.405 82.995 ;
        RECT 44.735 82.765 46.695 82.995 ;
        RECT 47.025 82.405 48.985 82.995 ;
        RECT 50.655 82.765 52.615 82.995 ;
        RECT 52.945 82.405 54.905 82.995 ;
        RECT 55.235 82.405 57.195 82.995 ;
        RECT 57.525 82.765 59.485 82.995 ;
        RECT 59.815 82.765 61.775 82.995 ;
        RECT 62.105 82.405 64.065 82.995 ;
        RECT 64.395 82.405 66.355 82.995 ;
        RECT 66.685 82.765 68.645 82.995 ;
        RECT 70.315 82.765 72.275 82.995 ;
        RECT 72.605 82.405 74.565 82.995 ;
        RECT 74.895 82.405 76.855 82.995 ;
        RECT 77.185 82.765 79.145 82.995 ;
        RECT 79.475 82.765 81.435 82.995 ;
        RECT 81.765 82.405 83.725 82.995 ;
        RECT 84.055 82.405 86.015 82.995 ;
        RECT 86.345 82.765 88.305 82.995 ;
        RECT 89.975 82.405 91.935 82.995 ;
        RECT 92.265 82.765 94.225 82.995 ;
        RECT 94.555 82.765 96.515 82.995 ;
        RECT 96.845 82.405 98.805 82.995 ;
        RECT 99.135 82.405 101.095 82.995 ;
        RECT 101.425 82.765 103.385 82.995 ;
        RECT 103.715 82.765 105.675 82.995 ;
        RECT 106.005 82.405 107.965 82.995 ;
        RECT 30.995 81.385 32.955 81.615 ;
        RECT 11.055 72.975 11.285 81.385 ;
        RECT 13.345 72.975 13.575 81.385 ;
        RECT 15.635 72.975 15.865 81.385 ;
        RECT 17.925 72.975 18.155 81.385 ;
        RECT 20.215 72.975 20.445 81.385 ;
        RECT 22.505 72.975 22.735 81.385 ;
        RECT 24.795 72.975 25.025 81.385 ;
        RECT 27.085 72.975 27.315 81.385 ;
        RECT 29.375 72.975 29.605 81.385 ;
        RECT 33.285 81.325 35.245 81.855 ;
        RECT 35.575 81.325 37.535 81.855 ;
        RECT 37.865 81.385 39.825 81.615 ;
        RECT 40.155 81.385 42.115 81.615 ;
        RECT 42.445 81.325 44.405 81.855 ;
        RECT 44.735 81.325 46.695 81.855 ;
        RECT 47.025 81.385 48.985 81.615 ;
        RECT 50.655 81.325 52.615 81.855 ;
        RECT 52.945 81.385 54.905 81.615 ;
        RECT 55.235 81.385 57.195 81.615 ;
        RECT 57.525 81.325 59.485 81.855 ;
        RECT 59.815 81.325 61.775 81.855 ;
        RECT 62.105 81.385 64.065 81.615 ;
        RECT 64.395 81.385 66.355 81.615 ;
        RECT 66.685 81.325 68.645 81.855 ;
        RECT 70.315 81.325 72.275 81.855 ;
        RECT 72.605 81.385 74.565 81.615 ;
        RECT 74.895 81.385 76.855 81.615 ;
        RECT 77.185 81.325 79.145 81.855 ;
        RECT 79.475 81.325 81.435 81.855 ;
        RECT 81.765 81.385 83.725 81.615 ;
        RECT 84.055 81.385 86.015 81.615 ;
        RECT 86.345 81.325 88.305 81.855 ;
        RECT 89.975 81.385 91.935 81.615 ;
        RECT 92.265 81.325 94.225 81.855 ;
        RECT 94.555 81.325 96.515 81.855 ;
        RECT 96.845 81.385 98.805 81.615 ;
        RECT 99.135 81.385 101.095 81.615 ;
        RECT 101.425 81.325 103.385 81.855 ;
        RECT 103.715 81.325 105.675 81.855 ;
        RECT 106.005 81.385 107.965 81.615 ;
        RECT 109.355 81.385 127.905 82.995 ;
        RECT 30.715 81.070 30.945 81.180 ;
        RECT 30.680 79.670 30.980 81.070 ;
        RECT 30.715 73.180 30.945 79.670 ;
        RECT 33.005 78.520 33.235 81.180 ;
        RECT 32.970 75.720 33.270 78.520 ;
        RECT 33.005 73.180 33.235 75.720 ;
        RECT 35.295 74.570 35.525 81.180 ;
        RECT 37.585 78.520 37.815 81.180 ;
        RECT 39.875 81.070 40.105 81.180 ;
        RECT 39.840 79.670 40.140 81.070 ;
        RECT 37.550 75.720 37.850 78.520 ;
        RECT 35.260 73.170 35.560 74.570 ;
        RECT 37.585 73.180 37.815 75.720 ;
        RECT 39.875 73.180 40.105 79.670 ;
        RECT 42.165 78.520 42.395 81.180 ;
        RECT 42.130 75.720 42.430 78.520 ;
        RECT 42.165 73.180 42.395 75.720 ;
        RECT 44.455 74.570 44.685 81.180 ;
        RECT 46.745 78.520 46.975 81.180 ;
        RECT 49.035 81.070 49.265 81.180 ;
        RECT 49.000 79.670 49.300 81.070 ;
        RECT 46.710 75.720 47.010 78.520 ;
        RECT 44.420 73.170 44.720 74.570 ;
        RECT 46.745 73.180 46.975 75.720 ;
        RECT 49.035 73.180 49.265 79.670 ;
        RECT 50.375 74.570 50.605 81.180 ;
        RECT 52.665 78.520 52.895 81.180 ;
        RECT 54.955 81.070 55.185 81.180 ;
        RECT 54.920 79.670 55.220 81.070 ;
        RECT 52.630 75.720 52.930 78.520 ;
        RECT 50.340 73.170 50.640 74.570 ;
        RECT 52.665 73.180 52.895 75.720 ;
        RECT 54.955 73.180 55.185 79.670 ;
        RECT 57.245 78.520 57.475 81.180 ;
        RECT 57.210 75.720 57.510 78.520 ;
        RECT 57.245 73.180 57.475 75.720 ;
        RECT 59.535 74.570 59.765 81.180 ;
        RECT 61.825 78.520 62.055 81.180 ;
        RECT 64.115 81.070 64.345 81.180 ;
        RECT 64.080 79.670 64.380 81.070 ;
        RECT 61.790 75.720 62.090 78.520 ;
        RECT 59.500 73.170 59.800 74.570 ;
        RECT 61.825 73.180 62.055 75.720 ;
        RECT 64.115 73.180 64.345 79.670 ;
        RECT 66.405 78.520 66.635 81.180 ;
        RECT 66.370 75.720 66.670 78.520 ;
        RECT 66.405 73.180 66.635 75.720 ;
        RECT 68.695 74.570 68.925 81.180 ;
        RECT 70.035 74.570 70.265 81.180 ;
        RECT 72.325 78.520 72.555 81.180 ;
        RECT 74.615 81.070 74.845 81.180 ;
        RECT 74.580 79.670 74.880 81.070 ;
        RECT 72.290 75.720 72.590 78.520 ;
        RECT 68.660 73.170 68.960 74.570 ;
        RECT 70.000 73.170 70.300 74.570 ;
        RECT 72.325 73.180 72.555 75.720 ;
        RECT 74.615 73.180 74.845 79.670 ;
        RECT 76.905 78.520 77.135 81.180 ;
        RECT 76.870 75.720 77.170 78.520 ;
        RECT 76.905 73.180 77.135 75.720 ;
        RECT 79.195 74.570 79.425 81.180 ;
        RECT 81.485 78.520 81.715 81.180 ;
        RECT 83.775 81.070 84.005 81.180 ;
        RECT 83.740 79.670 84.040 81.070 ;
        RECT 81.450 75.720 81.750 78.520 ;
        RECT 79.160 73.170 79.460 74.570 ;
        RECT 81.485 73.180 81.715 75.720 ;
        RECT 83.775 73.180 84.005 79.670 ;
        RECT 86.065 78.520 86.295 81.180 ;
        RECT 86.030 75.720 86.330 78.520 ;
        RECT 86.065 73.180 86.295 75.720 ;
        RECT 88.355 74.570 88.585 81.180 ;
        RECT 89.695 81.070 89.925 81.180 ;
        RECT 89.660 79.670 89.960 81.070 ;
        RECT 88.320 73.170 88.620 74.570 ;
        RECT 89.695 73.180 89.925 79.670 ;
        RECT 91.985 78.520 92.215 81.180 ;
        RECT 91.950 75.720 92.250 78.520 ;
        RECT 91.985 73.180 92.215 75.720 ;
        RECT 94.275 74.570 94.505 81.180 ;
        RECT 96.565 78.520 96.795 81.180 ;
        RECT 98.855 81.070 99.085 81.180 ;
        RECT 98.820 79.670 99.120 81.070 ;
        RECT 96.530 75.720 96.830 78.520 ;
        RECT 94.240 73.170 94.540 74.570 ;
        RECT 96.565 73.180 96.795 75.720 ;
        RECT 98.855 73.180 99.085 79.670 ;
        RECT 101.145 78.520 101.375 81.180 ;
        RECT 101.110 75.720 101.410 78.520 ;
        RECT 101.145 73.180 101.375 75.720 ;
        RECT 103.435 74.570 103.665 81.180 ;
        RECT 105.725 78.520 105.955 81.180 ;
        RECT 108.015 81.070 108.245 81.180 ;
        RECT 107.980 79.670 108.280 81.070 ;
        RECT 105.690 75.720 105.990 78.520 ;
        RECT 103.400 73.170 103.700 74.570 ;
        RECT 105.725 73.180 105.955 75.720 ;
        RECT 108.015 73.180 108.245 79.670 ;
        RECT 109.355 72.975 109.585 81.385 ;
        RECT 111.645 72.975 111.875 81.385 ;
        RECT 113.935 72.975 114.165 81.385 ;
        RECT 116.225 72.975 116.455 81.385 ;
        RECT 118.515 72.975 118.745 81.385 ;
        RECT 120.805 72.975 121.035 81.385 ;
        RECT 123.095 72.975 123.325 81.385 ;
        RECT 125.385 72.975 125.615 81.385 ;
        RECT 127.675 72.975 127.905 81.385 ;
        RECT 11.055 71.365 29.605 72.975 ;
        RECT 30.995 72.385 32.955 72.975 ;
        RECT 33.285 72.745 35.245 72.975 ;
        RECT 35.575 72.745 37.535 72.975 ;
        RECT 37.865 72.385 39.825 72.975 ;
        RECT 40.155 72.385 42.115 72.975 ;
        RECT 42.445 72.745 44.405 72.975 ;
        RECT 44.735 72.745 46.695 72.975 ;
        RECT 47.025 72.385 48.985 72.975 ;
        RECT 50.655 72.745 52.615 72.975 ;
        RECT 52.945 72.385 54.905 72.975 ;
        RECT 55.235 72.385 57.195 72.975 ;
        RECT 57.525 72.745 59.485 72.975 ;
        RECT 59.815 72.745 61.775 72.975 ;
        RECT 62.105 72.385 64.065 72.975 ;
        RECT 64.395 72.385 66.355 72.975 ;
        RECT 66.685 72.745 68.645 72.975 ;
        RECT 70.315 72.745 72.275 72.975 ;
        RECT 72.605 72.385 74.565 72.975 ;
        RECT 74.895 72.385 76.855 72.975 ;
        RECT 77.185 72.745 79.145 72.975 ;
        RECT 79.475 72.745 81.435 72.975 ;
        RECT 81.765 72.385 83.725 72.975 ;
        RECT 84.055 72.385 86.015 72.975 ;
        RECT 86.345 72.745 88.305 72.975 ;
        RECT 89.975 72.385 91.935 72.975 ;
        RECT 92.265 72.745 94.225 72.975 ;
        RECT 94.555 72.745 96.515 72.975 ;
        RECT 96.845 72.385 98.805 72.975 ;
        RECT 99.135 72.385 101.095 72.975 ;
        RECT 101.425 72.745 103.385 72.975 ;
        RECT 103.715 72.745 105.675 72.975 ;
        RECT 106.005 72.385 107.965 72.975 ;
        RECT 11.055 62.955 11.285 71.365 ;
        RECT 13.345 62.955 13.575 71.365 ;
        RECT 15.635 62.955 15.865 71.365 ;
        RECT 17.925 62.955 18.155 71.365 ;
        RECT 20.215 62.955 20.445 71.365 ;
        RECT 22.505 62.955 22.735 71.365 ;
        RECT 24.795 62.955 25.025 71.365 ;
        RECT 27.085 62.955 27.315 71.365 ;
        RECT 29.375 62.955 29.605 71.365 ;
        RECT 30.995 71.305 32.955 71.835 ;
        RECT 33.285 71.365 35.245 71.595 ;
        RECT 35.575 71.365 37.535 71.595 ;
        RECT 37.865 71.305 39.825 71.835 ;
        RECT 40.155 71.305 42.115 71.835 ;
        RECT 42.445 71.365 44.405 71.595 ;
        RECT 44.735 71.365 46.695 71.595 ;
        RECT 47.025 71.305 48.985 71.835 ;
        RECT 50.655 71.365 52.615 71.595 ;
        RECT 52.945 71.305 54.905 71.835 ;
        RECT 55.235 71.305 57.195 71.835 ;
        RECT 57.525 71.365 59.485 71.595 ;
        RECT 59.815 71.365 61.775 71.595 ;
        RECT 62.105 71.305 64.065 71.835 ;
        RECT 64.395 71.305 66.355 71.835 ;
        RECT 66.685 71.365 68.645 71.595 ;
        RECT 70.315 71.365 72.275 71.595 ;
        RECT 72.605 71.305 74.565 71.835 ;
        RECT 74.895 71.305 76.855 71.835 ;
        RECT 77.185 71.365 79.145 71.595 ;
        RECT 79.475 71.365 81.435 71.595 ;
        RECT 81.765 71.305 83.725 71.835 ;
        RECT 84.055 71.305 86.015 71.835 ;
        RECT 86.345 71.365 88.305 71.595 ;
        RECT 89.975 71.305 91.935 71.835 ;
        RECT 92.265 71.365 94.225 71.595 ;
        RECT 94.555 71.365 96.515 71.595 ;
        RECT 96.845 71.305 98.805 71.835 ;
        RECT 99.135 71.305 101.095 71.835 ;
        RECT 101.425 71.365 103.385 71.595 ;
        RECT 103.715 71.365 105.675 71.595 ;
        RECT 106.005 71.305 107.965 71.835 ;
        RECT 109.355 71.365 127.905 72.975 ;
        RECT 30.715 71.050 30.945 71.160 ;
        RECT 30.680 69.650 30.980 71.050 ;
        RECT 30.715 63.160 30.945 69.650 ;
        RECT 33.005 68.500 33.235 71.160 ;
        RECT 32.970 65.700 33.270 68.500 ;
        RECT 33.005 63.160 33.235 65.700 ;
        RECT 35.295 64.550 35.525 71.160 ;
        RECT 37.585 68.500 37.815 71.160 ;
        RECT 39.875 71.050 40.105 71.160 ;
        RECT 39.840 69.650 40.140 71.050 ;
        RECT 37.550 65.700 37.850 68.500 ;
        RECT 35.260 63.150 35.560 64.550 ;
        RECT 37.585 63.160 37.815 65.700 ;
        RECT 39.875 63.160 40.105 69.650 ;
        RECT 42.165 68.500 42.395 71.160 ;
        RECT 42.130 65.700 42.430 68.500 ;
        RECT 42.165 63.160 42.395 65.700 ;
        RECT 44.455 64.550 44.685 71.160 ;
        RECT 46.745 68.500 46.975 71.160 ;
        RECT 49.035 71.050 49.265 71.160 ;
        RECT 49.000 69.650 49.300 71.050 ;
        RECT 46.710 65.700 47.010 68.500 ;
        RECT 44.420 63.150 44.720 64.550 ;
        RECT 46.745 63.160 46.975 65.700 ;
        RECT 49.035 63.160 49.265 69.650 ;
        RECT 50.375 64.550 50.605 71.160 ;
        RECT 52.665 68.500 52.895 71.160 ;
        RECT 54.955 71.050 55.185 71.160 ;
        RECT 54.920 69.650 55.220 71.050 ;
        RECT 52.630 65.700 52.930 68.500 ;
        RECT 50.340 63.150 50.640 64.550 ;
        RECT 52.665 63.160 52.895 65.700 ;
        RECT 54.955 63.160 55.185 69.650 ;
        RECT 57.245 68.500 57.475 71.160 ;
        RECT 57.210 65.700 57.510 68.500 ;
        RECT 57.245 63.160 57.475 65.700 ;
        RECT 59.535 64.550 59.765 71.160 ;
        RECT 61.825 68.500 62.055 71.160 ;
        RECT 64.115 71.050 64.345 71.160 ;
        RECT 64.080 69.650 64.380 71.050 ;
        RECT 61.790 65.700 62.090 68.500 ;
        RECT 59.500 63.150 59.800 64.550 ;
        RECT 61.825 63.160 62.055 65.700 ;
        RECT 64.115 63.160 64.345 69.650 ;
        RECT 66.405 68.500 66.635 71.160 ;
        RECT 66.370 65.700 66.670 68.500 ;
        RECT 66.405 63.160 66.635 65.700 ;
        RECT 68.695 64.550 68.925 71.160 ;
        RECT 70.035 64.550 70.265 71.160 ;
        RECT 72.325 68.500 72.555 71.160 ;
        RECT 74.615 71.050 74.845 71.160 ;
        RECT 74.580 69.650 74.880 71.050 ;
        RECT 72.290 65.700 72.590 68.500 ;
        RECT 68.660 63.150 68.960 64.550 ;
        RECT 70.000 63.150 70.300 64.550 ;
        RECT 72.325 63.160 72.555 65.700 ;
        RECT 74.615 63.160 74.845 69.650 ;
        RECT 76.905 68.500 77.135 71.160 ;
        RECT 76.870 65.700 77.170 68.500 ;
        RECT 76.905 63.160 77.135 65.700 ;
        RECT 79.195 64.550 79.425 71.160 ;
        RECT 81.485 68.500 81.715 71.160 ;
        RECT 83.775 71.050 84.005 71.160 ;
        RECT 83.740 69.650 84.040 71.050 ;
        RECT 81.450 65.700 81.750 68.500 ;
        RECT 79.160 63.150 79.460 64.550 ;
        RECT 81.485 63.160 81.715 65.700 ;
        RECT 83.775 63.160 84.005 69.650 ;
        RECT 86.065 68.500 86.295 71.160 ;
        RECT 86.030 65.700 86.330 68.500 ;
        RECT 86.065 63.160 86.295 65.700 ;
        RECT 88.355 64.550 88.585 71.160 ;
        RECT 89.695 71.050 89.925 71.160 ;
        RECT 89.660 69.650 89.960 71.050 ;
        RECT 88.320 63.150 88.620 64.550 ;
        RECT 89.695 63.160 89.925 69.650 ;
        RECT 91.985 68.500 92.215 71.160 ;
        RECT 91.950 65.700 92.250 68.500 ;
        RECT 91.985 63.160 92.215 65.700 ;
        RECT 94.275 64.550 94.505 71.160 ;
        RECT 96.565 68.500 96.795 71.160 ;
        RECT 98.855 71.050 99.085 71.160 ;
        RECT 98.820 69.650 99.120 71.050 ;
        RECT 96.530 65.700 96.830 68.500 ;
        RECT 94.240 63.150 94.540 64.550 ;
        RECT 96.565 63.160 96.795 65.700 ;
        RECT 98.855 63.160 99.085 69.650 ;
        RECT 101.145 68.500 101.375 71.160 ;
        RECT 101.110 65.700 101.410 68.500 ;
        RECT 101.145 63.160 101.375 65.700 ;
        RECT 103.435 64.550 103.665 71.160 ;
        RECT 105.725 68.500 105.955 71.160 ;
        RECT 108.015 71.050 108.245 71.160 ;
        RECT 107.980 69.650 108.280 71.050 ;
        RECT 105.690 65.700 105.990 68.500 ;
        RECT 103.400 63.150 103.700 64.550 ;
        RECT 105.725 63.160 105.955 65.700 ;
        RECT 108.015 63.160 108.245 69.650 ;
        RECT 109.355 62.955 109.585 71.365 ;
        RECT 111.645 62.955 111.875 71.365 ;
        RECT 113.935 62.955 114.165 71.365 ;
        RECT 116.225 62.955 116.455 71.365 ;
        RECT 118.515 62.955 118.745 71.365 ;
        RECT 120.805 62.955 121.035 71.365 ;
        RECT 123.095 62.955 123.325 71.365 ;
        RECT 125.385 62.955 125.615 71.365 ;
        RECT 127.675 62.955 127.905 71.365 ;
        RECT 11.055 61.345 29.605 62.955 ;
        RECT 30.995 62.725 32.955 62.955 ;
        RECT 33.285 62.365 35.245 62.955 ;
        RECT 35.575 62.365 37.535 62.955 ;
        RECT 37.865 62.725 39.825 62.955 ;
        RECT 40.155 62.725 42.115 62.955 ;
        RECT 42.445 62.365 44.405 62.955 ;
        RECT 44.735 62.365 46.695 62.955 ;
        RECT 47.025 62.725 48.985 62.955 ;
        RECT 50.655 62.365 52.615 62.955 ;
        RECT 52.945 62.725 54.905 62.955 ;
        RECT 55.235 62.725 57.195 62.955 ;
        RECT 57.525 62.365 59.485 62.955 ;
        RECT 59.815 62.365 61.775 62.955 ;
        RECT 62.105 62.725 64.065 62.955 ;
        RECT 64.395 62.725 66.355 62.955 ;
        RECT 66.685 62.365 68.645 62.955 ;
        RECT 70.315 62.365 72.275 62.955 ;
        RECT 72.605 62.725 74.565 62.955 ;
        RECT 74.895 62.725 76.855 62.955 ;
        RECT 77.185 62.365 79.145 62.955 ;
        RECT 79.475 62.365 81.435 62.955 ;
        RECT 81.765 62.725 83.725 62.955 ;
        RECT 84.055 62.725 86.015 62.955 ;
        RECT 86.345 62.365 88.305 62.955 ;
        RECT 89.975 62.725 91.935 62.955 ;
        RECT 92.265 62.365 94.225 62.955 ;
        RECT 94.555 62.365 96.515 62.955 ;
        RECT 96.845 62.725 98.805 62.955 ;
        RECT 99.135 62.725 101.095 62.955 ;
        RECT 101.425 62.365 103.385 62.955 ;
        RECT 103.715 62.365 105.675 62.955 ;
        RECT 106.005 62.725 107.965 62.955 ;
        RECT 11.055 52.935 11.285 61.345 ;
        RECT 13.345 52.935 13.575 61.345 ;
        RECT 15.635 52.935 15.865 61.345 ;
        RECT 17.925 52.935 18.155 61.345 ;
        RECT 20.215 52.935 20.445 61.345 ;
        RECT 22.505 52.935 22.735 61.345 ;
        RECT 24.795 52.935 25.025 61.345 ;
        RECT 27.085 52.935 27.315 61.345 ;
        RECT 29.375 52.935 29.605 61.345 ;
        RECT 30.995 61.285 32.955 61.815 ;
        RECT 33.285 61.345 35.245 61.575 ;
        RECT 35.575 61.345 37.535 61.575 ;
        RECT 37.865 61.285 39.825 61.815 ;
        RECT 40.155 61.285 42.115 61.815 ;
        RECT 42.445 61.345 44.405 61.575 ;
        RECT 44.735 61.345 46.695 61.575 ;
        RECT 47.025 61.285 48.985 61.815 ;
        RECT 50.655 61.345 52.615 61.575 ;
        RECT 52.945 61.285 54.905 61.815 ;
        RECT 55.235 61.285 57.195 61.815 ;
        RECT 57.525 61.345 59.485 61.575 ;
        RECT 59.815 61.345 61.775 61.575 ;
        RECT 62.105 61.285 64.065 61.815 ;
        RECT 64.395 61.285 66.355 61.815 ;
        RECT 66.685 61.345 68.645 61.575 ;
        RECT 70.315 61.345 72.275 61.575 ;
        RECT 72.605 61.285 74.565 61.815 ;
        RECT 74.895 61.285 76.855 61.815 ;
        RECT 77.185 61.345 79.145 61.575 ;
        RECT 79.475 61.345 81.435 61.575 ;
        RECT 81.765 61.285 83.725 61.815 ;
        RECT 84.055 61.285 86.015 61.815 ;
        RECT 86.345 61.345 88.305 61.575 ;
        RECT 89.975 61.285 91.935 61.815 ;
        RECT 92.265 61.345 94.225 61.575 ;
        RECT 94.555 61.345 96.515 61.575 ;
        RECT 96.845 61.285 98.805 61.815 ;
        RECT 99.135 61.285 101.095 61.815 ;
        RECT 101.425 61.345 103.385 61.575 ;
        RECT 103.715 61.345 105.675 61.575 ;
        RECT 106.005 61.285 107.965 61.815 ;
        RECT 109.355 61.345 127.905 62.955 ;
        RECT 30.715 54.530 30.945 61.140 ;
        RECT 33.005 58.480 33.235 61.140 ;
        RECT 35.295 61.030 35.525 61.140 ;
        RECT 35.260 59.630 35.560 61.030 ;
        RECT 32.970 55.680 33.270 58.480 ;
        RECT 30.680 53.130 30.980 54.530 ;
        RECT 33.005 53.140 33.235 55.680 ;
        RECT 35.295 53.140 35.525 59.630 ;
        RECT 37.585 58.480 37.815 61.140 ;
        RECT 37.550 55.680 37.850 58.480 ;
        RECT 37.585 53.140 37.815 55.680 ;
        RECT 39.875 54.530 40.105 61.140 ;
        RECT 42.165 58.480 42.395 61.140 ;
        RECT 44.455 61.030 44.685 61.140 ;
        RECT 44.420 59.630 44.720 61.030 ;
        RECT 42.130 55.680 42.430 58.480 ;
        RECT 39.840 53.130 40.140 54.530 ;
        RECT 42.165 53.140 42.395 55.680 ;
        RECT 44.455 53.140 44.685 59.630 ;
        RECT 46.745 58.480 46.975 61.140 ;
        RECT 46.710 55.680 47.010 58.480 ;
        RECT 46.745 53.140 46.975 55.680 ;
        RECT 49.035 54.530 49.265 61.140 ;
        RECT 50.375 61.030 50.605 61.140 ;
        RECT 50.340 59.630 50.640 61.030 ;
        RECT 49.000 53.130 49.300 54.530 ;
        RECT 50.375 53.140 50.605 59.630 ;
        RECT 52.665 58.480 52.895 61.140 ;
        RECT 52.630 55.680 52.930 58.480 ;
        RECT 52.665 53.140 52.895 55.680 ;
        RECT 54.955 54.530 55.185 61.140 ;
        RECT 57.245 58.480 57.475 61.140 ;
        RECT 59.535 61.030 59.765 61.140 ;
        RECT 59.500 59.630 59.800 61.030 ;
        RECT 57.210 55.680 57.510 58.480 ;
        RECT 54.920 53.130 55.220 54.530 ;
        RECT 57.245 53.140 57.475 55.680 ;
        RECT 59.535 53.140 59.765 59.630 ;
        RECT 61.825 58.480 62.055 61.140 ;
        RECT 61.790 55.680 62.090 58.480 ;
        RECT 61.825 53.140 62.055 55.680 ;
        RECT 64.115 54.530 64.345 61.140 ;
        RECT 66.405 58.480 66.635 61.140 ;
        RECT 68.695 61.030 68.925 61.140 ;
        RECT 70.035 61.030 70.265 61.140 ;
        RECT 68.660 59.630 68.960 61.030 ;
        RECT 70.000 59.630 70.300 61.030 ;
        RECT 66.370 55.680 66.670 58.480 ;
        RECT 64.080 53.130 64.380 54.530 ;
        RECT 66.405 53.140 66.635 55.680 ;
        RECT 68.695 53.140 68.925 59.630 ;
        RECT 70.035 53.140 70.265 59.630 ;
        RECT 72.325 58.480 72.555 61.140 ;
        RECT 72.290 55.680 72.590 58.480 ;
        RECT 72.325 53.140 72.555 55.680 ;
        RECT 74.615 54.530 74.845 61.140 ;
        RECT 76.905 58.480 77.135 61.140 ;
        RECT 79.195 61.030 79.425 61.140 ;
        RECT 79.160 59.630 79.460 61.030 ;
        RECT 76.870 55.680 77.170 58.480 ;
        RECT 74.580 53.130 74.880 54.530 ;
        RECT 76.905 53.140 77.135 55.680 ;
        RECT 79.195 53.140 79.425 59.630 ;
        RECT 81.485 58.480 81.715 61.140 ;
        RECT 81.450 55.680 81.750 58.480 ;
        RECT 81.485 53.140 81.715 55.680 ;
        RECT 83.775 54.530 84.005 61.140 ;
        RECT 86.065 58.480 86.295 61.140 ;
        RECT 88.355 61.030 88.585 61.140 ;
        RECT 88.320 59.630 88.620 61.030 ;
        RECT 86.030 55.680 86.330 58.480 ;
        RECT 83.740 53.130 84.040 54.530 ;
        RECT 86.065 53.140 86.295 55.680 ;
        RECT 88.355 53.140 88.585 59.630 ;
        RECT 89.695 54.530 89.925 61.140 ;
        RECT 91.985 58.480 92.215 61.140 ;
        RECT 94.275 61.030 94.505 61.140 ;
        RECT 94.240 59.630 94.540 61.030 ;
        RECT 91.950 55.680 92.250 58.480 ;
        RECT 89.660 53.130 89.960 54.530 ;
        RECT 91.985 53.140 92.215 55.680 ;
        RECT 94.275 53.140 94.505 59.630 ;
        RECT 96.565 58.480 96.795 61.140 ;
        RECT 96.530 55.680 96.830 58.480 ;
        RECT 96.565 53.140 96.795 55.680 ;
        RECT 98.855 54.530 99.085 61.140 ;
        RECT 101.145 58.480 101.375 61.140 ;
        RECT 103.435 61.030 103.665 61.140 ;
        RECT 103.400 59.630 103.700 61.030 ;
        RECT 101.110 55.680 101.410 58.480 ;
        RECT 98.820 53.130 99.120 54.530 ;
        RECT 101.145 53.140 101.375 55.680 ;
        RECT 103.435 53.140 103.665 59.630 ;
        RECT 105.725 58.480 105.955 61.140 ;
        RECT 105.690 55.680 105.990 58.480 ;
        RECT 105.725 53.140 105.955 55.680 ;
        RECT 108.015 54.530 108.245 61.140 ;
        RECT 107.980 53.130 108.280 54.530 ;
        RECT 109.355 52.935 109.585 61.345 ;
        RECT 111.645 52.935 111.875 61.345 ;
        RECT 113.935 52.935 114.165 61.345 ;
        RECT 116.225 52.935 116.455 61.345 ;
        RECT 118.515 52.935 118.745 61.345 ;
        RECT 120.805 52.935 121.035 61.345 ;
        RECT 123.095 52.935 123.325 61.345 ;
        RECT 125.385 52.935 125.615 61.345 ;
        RECT 127.675 52.935 127.905 61.345 ;
        RECT 11.055 51.325 29.605 52.935 ;
        RECT 30.995 52.705 32.955 52.935 ;
        RECT 33.285 52.345 35.245 52.935 ;
        RECT 35.575 52.345 37.535 52.935 ;
        RECT 37.865 52.705 39.825 52.935 ;
        RECT 40.155 52.705 42.115 52.935 ;
        RECT 42.445 52.345 44.405 52.935 ;
        RECT 44.735 52.345 46.695 52.935 ;
        RECT 47.025 52.705 48.985 52.935 ;
        RECT 50.655 52.345 52.615 52.935 ;
        RECT 52.945 52.705 54.905 52.935 ;
        RECT 55.235 52.705 57.195 52.935 ;
        RECT 57.525 52.345 59.485 52.935 ;
        RECT 59.815 52.345 61.775 52.935 ;
        RECT 62.105 52.705 64.065 52.935 ;
        RECT 64.395 52.705 66.355 52.935 ;
        RECT 66.685 52.345 68.645 52.935 ;
        RECT 70.315 52.345 72.275 52.935 ;
        RECT 72.605 52.705 74.565 52.935 ;
        RECT 74.895 52.705 76.855 52.935 ;
        RECT 77.185 52.345 79.145 52.935 ;
        RECT 79.475 52.345 81.435 52.935 ;
        RECT 81.765 52.705 83.725 52.935 ;
        RECT 84.055 52.705 86.015 52.935 ;
        RECT 86.345 52.345 88.305 52.935 ;
        RECT 89.975 52.705 91.935 52.935 ;
        RECT 92.265 52.345 94.225 52.935 ;
        RECT 94.555 52.345 96.515 52.935 ;
        RECT 96.845 52.705 98.805 52.935 ;
        RECT 99.135 52.705 101.095 52.935 ;
        RECT 101.425 52.345 103.385 52.935 ;
        RECT 103.715 52.345 105.675 52.935 ;
        RECT 106.005 52.705 107.965 52.935 ;
        RECT 30.995 51.325 32.955 51.555 ;
        RECT 33.285 51.325 35.245 51.555 ;
        RECT 35.575 51.325 37.535 51.555 ;
        RECT 37.865 51.325 39.825 51.555 ;
        RECT 40.155 51.325 42.115 51.555 ;
        RECT 42.445 51.325 44.405 51.555 ;
        RECT 44.735 51.325 46.695 51.555 ;
        RECT 47.025 51.325 48.985 51.555 ;
        RECT 50.655 51.325 52.615 51.555 ;
        RECT 52.945 51.325 54.905 51.555 ;
        RECT 55.235 51.325 57.195 51.555 ;
        RECT 57.525 51.325 59.485 51.555 ;
        RECT 59.815 51.325 61.775 51.555 ;
        RECT 62.105 51.325 64.065 51.555 ;
        RECT 64.395 51.325 66.355 51.555 ;
        RECT 66.685 51.325 68.645 51.555 ;
        RECT 70.315 51.325 72.275 51.555 ;
        RECT 72.605 51.325 74.565 51.555 ;
        RECT 74.895 51.325 76.855 51.555 ;
        RECT 77.185 51.325 79.145 51.555 ;
        RECT 79.475 51.325 81.435 51.555 ;
        RECT 81.765 51.325 83.725 51.555 ;
        RECT 84.055 51.325 86.015 51.555 ;
        RECT 86.345 51.325 88.305 51.555 ;
        RECT 89.975 51.325 91.935 51.555 ;
        RECT 92.265 51.325 94.225 51.555 ;
        RECT 94.555 51.325 96.515 51.555 ;
        RECT 96.845 51.325 98.805 51.555 ;
        RECT 99.135 51.325 101.095 51.555 ;
        RECT 101.425 51.325 103.385 51.555 ;
        RECT 103.715 51.325 105.675 51.555 ;
        RECT 106.005 51.325 107.965 51.555 ;
        RECT 109.355 51.325 127.905 52.935 ;
        RECT 11.055 42.915 11.285 51.325 ;
        RECT 13.345 42.915 13.575 51.325 ;
        RECT 15.635 42.915 15.865 51.325 ;
        RECT 17.925 42.915 18.155 51.325 ;
        RECT 20.215 42.915 20.445 51.325 ;
        RECT 22.505 42.915 22.735 51.325 ;
        RECT 24.795 42.915 25.025 51.325 ;
        RECT 27.085 42.915 27.315 51.325 ;
        RECT 29.375 42.915 29.605 51.325 ;
        RECT 11.055 42.225 29.605 42.915 ;
        RECT 30.715 42.915 30.945 51.120 ;
        RECT 33.005 42.915 33.235 51.120 ;
        RECT 35.295 42.915 35.525 51.120 ;
        RECT 37.585 42.915 37.815 51.120 ;
        RECT 39.875 42.915 40.105 51.120 ;
        RECT 42.165 42.915 42.395 51.120 ;
        RECT 44.455 42.915 44.685 51.120 ;
        RECT 46.745 42.915 46.975 51.120 ;
        RECT 49.035 42.915 49.265 51.120 ;
        RECT 30.715 42.225 49.265 42.915 ;
        RECT 50.375 42.915 50.605 51.120 ;
        RECT 52.665 42.915 52.895 51.120 ;
        RECT 54.955 42.915 55.185 51.120 ;
        RECT 57.245 42.915 57.475 51.120 ;
        RECT 59.535 42.915 59.765 51.120 ;
        RECT 61.825 42.915 62.055 51.120 ;
        RECT 64.115 42.915 64.345 51.120 ;
        RECT 66.405 42.915 66.635 51.120 ;
        RECT 68.695 42.915 68.925 51.120 ;
        RECT 50.375 42.225 68.925 42.915 ;
        RECT 70.035 42.915 70.265 51.120 ;
        RECT 72.325 42.915 72.555 51.120 ;
        RECT 74.615 42.915 74.845 51.120 ;
        RECT 76.905 42.915 77.135 51.120 ;
        RECT 79.195 42.915 79.425 51.120 ;
        RECT 81.485 42.915 81.715 51.120 ;
        RECT 83.775 42.915 84.005 51.120 ;
        RECT 86.065 42.915 86.295 51.120 ;
        RECT 88.355 42.915 88.585 51.120 ;
        RECT 70.035 42.225 88.585 42.915 ;
        RECT 89.695 42.915 89.925 51.120 ;
        RECT 91.985 42.915 92.215 51.120 ;
        RECT 94.275 42.915 94.505 51.120 ;
        RECT 96.565 42.915 96.795 51.120 ;
        RECT 98.855 42.915 99.085 51.120 ;
        RECT 101.145 42.915 101.375 51.120 ;
        RECT 103.435 42.915 103.665 51.120 ;
        RECT 105.725 42.915 105.955 51.120 ;
        RECT 108.015 42.915 108.245 51.120 ;
        RECT 89.695 42.225 108.245 42.915 ;
        RECT 109.355 42.915 109.585 51.325 ;
        RECT 111.645 42.915 111.875 51.325 ;
        RECT 113.935 42.915 114.165 51.325 ;
        RECT 116.225 42.915 116.455 51.325 ;
        RECT 118.515 42.915 118.745 51.325 ;
        RECT 120.805 42.915 121.035 51.325 ;
        RECT 123.095 42.915 123.325 51.325 ;
        RECT 125.385 42.915 125.615 51.325 ;
        RECT 127.675 42.915 127.905 51.325 ;
        RECT 109.355 42.225 127.905 42.915 ;
        RECT 128.345 42.225 135.710 102.115 ;
        RECT 136.295 100.155 138.400 101.915 ;
        RECT 136.295 97.815 138.400 99.575 ;
        RECT 136.295 95.475 138.400 97.235 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 141.695 93.725 142.995 108.925 ;
        RECT 149.570 107.765 155.900 137.690 ;
        RECT 146.290 104.835 155.900 107.765 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 146.290 101.325 148.395 103.085 ;
        RECT 146.290 98.985 148.395 100.745 ;
        RECT 146.290 96.645 148.395 98.405 ;
        RECT 146.290 94.305 148.395 96.065 ;
        RECT 136.295 91.965 138.400 93.725 ;
        RECT 141.695 93.135 148.395 93.725 ;
        RECT 146.290 91.965 148.395 92.555 ;
        RECT 136.295 90.795 143.395 91.385 ;
        RECT 136.295 89.625 138.400 90.215 ;
        RECT 146.290 89.625 148.395 91.385 ;
        RECT 136.295 87.285 138.400 89.045 ;
        RECT 146.290 88.455 148.395 89.045 ;
        RECT 146.290 87.285 148.395 87.875 ;
        RECT 136.295 86.115 138.400 86.705 ;
        RECT 136.295 84.945 138.400 85.535 ;
        RECT 146.290 84.945 148.395 86.705 ;
        RECT 136.295 82.605 138.400 84.365 ;
        RECT 146.290 83.775 148.395 84.365 ;
        RECT 146.290 82.605 148.395 83.195 ;
        RECT 136.295 81.435 141.260 82.025 ;
        RECT 143.790 81.435 148.395 82.025 ;
        RECT 136.295 80.265 138.400 80.855 ;
        RECT 136.295 79.095 138.400 79.685 ;
        RECT 136.295 76.755 138.400 78.515 ;
        RECT 136.295 75.585 138.400 76.175 ;
        RECT 136.295 74.415 138.400 75.005 ;
        RECT 136.295 72.075 138.400 73.835 ;
        RECT 136.295 70.905 138.400 71.495 ;
        RECT 136.295 69.735 138.400 70.325 ;
        RECT 136.295 67.395 138.400 69.155 ;
        RECT 136.295 66.225 138.400 66.815 ;
        RECT 136.295 65.055 138.400 65.645 ;
        RECT 136.295 62.715 138.400 64.475 ;
        RECT 143.790 62.135 145.190 81.435 ;
        RECT 146.290 79.095 148.395 80.855 ;
        RECT 146.290 77.925 148.395 78.515 ;
        RECT 146.290 76.755 148.395 77.345 ;
        RECT 146.290 74.415 148.395 76.175 ;
        RECT 146.290 73.245 148.395 73.835 ;
        RECT 146.290 72.075 148.395 72.665 ;
        RECT 146.290 69.735 148.395 71.495 ;
        RECT 146.290 68.565 148.395 69.155 ;
        RECT 146.290 67.395 148.395 67.985 ;
        RECT 146.290 65.055 148.395 66.815 ;
        RECT 146.290 63.885 148.395 64.475 ;
        RECT 146.290 62.715 148.395 63.305 ;
        RECT 136.295 61.545 140.910 62.135 ;
        RECT 143.790 61.545 148.395 62.135 ;
        RECT 136.295 60.375 138.400 60.965 ;
        RECT 136.295 59.205 138.400 59.795 ;
        RECT 136.295 56.865 138.400 58.625 ;
        RECT 136.295 55.695 138.400 56.285 ;
        RECT 136.295 54.525 138.400 55.115 ;
        RECT 136.295 52.185 138.400 53.945 ;
        RECT 136.295 51.015 138.400 51.605 ;
        RECT 136.295 49.845 138.400 50.435 ;
        RECT 136.295 47.505 138.400 49.265 ;
        RECT 136.295 46.335 138.400 46.925 ;
        RECT 136.295 45.165 138.400 45.755 ;
        RECT 136.295 42.825 138.400 44.585 ;
        RECT 139.510 42.245 140.910 61.545 ;
        RECT 146.290 59.205 148.395 60.965 ;
        RECT 146.290 58.035 148.395 58.625 ;
        RECT 146.290 56.865 148.395 57.455 ;
        RECT 146.290 54.525 148.395 56.285 ;
        RECT 146.290 53.355 148.395 53.945 ;
        RECT 146.290 52.185 148.395 52.775 ;
        RECT 146.290 49.845 148.395 51.605 ;
        RECT 146.290 48.675 148.395 49.265 ;
        RECT 146.290 47.505 148.395 48.095 ;
        RECT 146.290 45.165 148.395 46.925 ;
        RECT 146.290 43.995 148.395 44.585 ;
        RECT 146.290 42.825 148.395 43.415 ;
        RECT 4.100 41.635 135.710 42.225 ;
        RECT 136.295 41.655 140.910 42.245 ;
        RECT 143.435 41.655 148.395 42.245 ;
        RECT 4.100 4.900 4.900 41.635 ;
        RECT 7.065 39.040 130.565 39.630 ;
        RECT 7.065 36.430 10.615 39.040 ;
        RECT 8.665 9.480 10.615 36.430 ;
        RECT 11.115 38.350 20.505 38.580 ;
        RECT 22.015 38.350 30.845 38.650 ;
        RECT 32.635 38.350 41.465 38.650 ;
        RECT 43.255 38.350 52.085 38.650 ;
        RECT 53.875 38.350 62.705 38.650 ;
        RECT 64.215 38.350 73.605 38.580 ;
        RECT 11.115 34.890 11.345 38.350 ;
        RECT 13.405 34.890 13.635 38.190 ;
        RECT 15.695 34.890 15.925 38.350 ;
        RECT 17.985 34.890 18.215 38.190 ;
        RECT 20.275 34.890 20.505 38.350 ;
        RECT 11.020 33.490 11.345 34.890 ;
        RECT 13.370 33.490 13.670 34.890 ;
        RECT 15.660 33.490 15.960 34.890 ;
        RECT 17.950 33.490 18.250 34.890 ;
        RECT 20.240 33.490 20.540 34.890 ;
        RECT 11.115 30.030 11.345 33.490 ;
        RECT 13.405 30.190 13.635 33.490 ;
        RECT 15.695 30.030 15.925 33.490 ;
        RECT 17.985 30.190 18.215 33.490 ;
        RECT 20.275 30.030 20.505 33.490 ;
        RECT 21.735 32.890 21.965 38.190 ;
        RECT 24.025 34.890 24.255 38.190 ;
        RECT 26.315 36.890 26.545 38.190 ;
        RECT 26.280 35.490 26.580 36.890 ;
        RECT 23.990 33.490 24.290 34.890 ;
        RECT 21.700 31.490 22.000 32.890 ;
        RECT 21.735 30.190 21.965 31.490 ;
        RECT 24.025 30.190 24.255 33.490 ;
        RECT 26.315 30.190 26.545 35.490 ;
        RECT 28.605 34.890 28.835 38.190 ;
        RECT 28.570 33.490 28.870 34.890 ;
        RECT 28.605 30.190 28.835 33.490 ;
        RECT 30.895 32.890 31.125 38.190 ;
        RECT 32.355 36.890 32.585 38.190 ;
        RECT 32.320 35.490 32.620 36.890 ;
        RECT 30.860 31.490 31.160 32.890 ;
        RECT 30.895 30.190 31.125 31.490 ;
        RECT 32.355 30.190 32.585 35.490 ;
        RECT 34.645 34.890 34.875 38.190 ;
        RECT 34.610 33.490 34.910 34.890 ;
        RECT 34.645 30.190 34.875 33.490 ;
        RECT 36.935 32.890 37.165 38.190 ;
        RECT 39.225 34.890 39.455 38.190 ;
        RECT 41.515 36.890 41.745 38.190 ;
        RECT 41.480 35.490 41.780 36.890 ;
        RECT 39.190 33.490 39.490 34.890 ;
        RECT 36.900 31.490 37.200 32.890 ;
        RECT 36.935 30.190 37.165 31.490 ;
        RECT 39.225 30.190 39.455 33.490 ;
        RECT 41.515 30.190 41.745 35.490 ;
        RECT 42.975 32.890 43.205 38.190 ;
        RECT 45.265 34.890 45.495 38.190 ;
        RECT 47.555 36.890 47.785 38.190 ;
        RECT 47.520 35.490 47.820 36.890 ;
        RECT 45.230 33.490 45.530 34.890 ;
        RECT 42.940 31.490 43.240 32.890 ;
        RECT 42.975 30.190 43.205 31.490 ;
        RECT 45.265 30.190 45.495 33.490 ;
        RECT 47.555 30.190 47.785 35.490 ;
        RECT 49.845 34.890 50.075 38.190 ;
        RECT 49.810 33.490 50.110 34.890 ;
        RECT 49.845 30.190 50.075 33.490 ;
        RECT 52.135 32.890 52.365 38.190 ;
        RECT 53.595 36.890 53.825 38.190 ;
        RECT 53.560 35.490 53.860 36.890 ;
        RECT 52.100 31.490 52.400 32.890 ;
        RECT 52.135 30.190 52.365 31.490 ;
        RECT 53.595 30.190 53.825 35.490 ;
        RECT 55.885 34.890 56.115 38.190 ;
        RECT 55.850 33.490 56.150 34.890 ;
        RECT 55.885 30.190 56.115 33.490 ;
        RECT 58.175 32.890 58.405 38.190 ;
        RECT 60.465 34.890 60.695 38.190 ;
        RECT 62.755 36.890 62.985 38.190 ;
        RECT 62.720 35.490 63.020 36.890 ;
        RECT 60.430 33.490 60.730 34.890 ;
        RECT 58.140 31.490 58.440 32.890 ;
        RECT 58.175 30.190 58.405 31.490 ;
        RECT 60.465 30.190 60.695 33.490 ;
        RECT 62.755 30.190 62.985 35.490 ;
        RECT 64.215 34.890 64.445 38.350 ;
        RECT 66.505 34.890 66.735 38.190 ;
        RECT 68.795 34.890 69.025 38.350 ;
        RECT 71.085 34.890 71.315 38.190 ;
        RECT 73.375 34.890 73.605 38.350 ;
        RECT 64.180 33.490 64.480 34.890 ;
        RECT 66.470 33.490 66.770 34.890 ;
        RECT 68.760 33.490 69.060 34.890 ;
        RECT 71.050 33.490 71.350 34.890 ;
        RECT 73.340 33.490 73.640 34.890 ;
        RECT 64.215 30.030 64.445 33.490 ;
        RECT 66.505 30.190 66.735 33.490 ;
        RECT 68.795 30.030 69.025 33.490 ;
        RECT 71.085 30.190 71.315 33.490 ;
        RECT 73.375 30.030 73.605 33.490 ;
        RECT 11.115 29.800 20.505 30.030 ;
        RECT 22.015 29.730 30.845 30.030 ;
        RECT 32.635 29.730 41.465 30.030 ;
        RECT 43.255 29.730 52.085 30.030 ;
        RECT 53.875 29.730 62.705 30.030 ;
        RECT 64.215 29.800 73.605 30.030 ;
        RECT 11.115 28.420 20.505 28.650 ;
        RECT 22.015 28.420 30.845 28.720 ;
        RECT 32.635 28.650 41.465 28.720 ;
        RECT 43.255 28.650 52.085 28.720 ;
        RECT 32.355 28.420 41.745 28.650 ;
        RECT 11.115 24.960 11.345 28.420 ;
        RECT 13.405 24.960 13.635 28.260 ;
        RECT 15.695 24.960 15.925 28.420 ;
        RECT 17.985 24.960 18.215 28.260 ;
        RECT 20.275 24.960 20.505 28.420 ;
        RECT 21.735 26.960 21.965 28.260 ;
        RECT 21.700 25.560 22.000 26.960 ;
        RECT 11.020 23.560 11.345 24.960 ;
        RECT 13.370 23.560 13.670 24.960 ;
        RECT 15.660 23.560 15.960 24.960 ;
        RECT 17.950 23.560 18.250 24.960 ;
        RECT 20.240 23.560 20.540 24.960 ;
        RECT 11.115 20.100 11.345 23.560 ;
        RECT 13.405 20.260 13.635 23.560 ;
        RECT 15.695 20.100 15.925 23.560 ;
        RECT 17.985 20.260 18.215 23.560 ;
        RECT 20.275 20.100 20.505 23.560 ;
        RECT 21.735 20.260 21.965 25.560 ;
        RECT 24.025 24.960 24.255 28.260 ;
        RECT 23.990 23.560 24.290 24.960 ;
        RECT 24.025 20.260 24.255 23.560 ;
        RECT 26.315 22.960 26.545 28.260 ;
        RECT 28.605 24.960 28.835 28.260 ;
        RECT 30.895 26.960 31.125 28.260 ;
        RECT 30.860 25.560 31.160 26.960 ;
        RECT 28.570 23.560 28.870 24.960 ;
        RECT 26.280 21.560 26.580 22.960 ;
        RECT 26.315 20.260 26.545 21.560 ;
        RECT 28.605 20.260 28.835 23.560 ;
        RECT 30.895 20.260 31.125 25.560 ;
        RECT 32.355 20.100 32.585 28.420 ;
        RECT 34.645 24.960 34.875 28.260 ;
        RECT 34.610 23.560 34.910 24.960 ;
        RECT 34.645 20.260 34.875 23.560 ;
        RECT 36.935 20.100 37.165 28.420 ;
        RECT 39.225 24.960 39.455 28.260 ;
        RECT 39.190 23.560 39.490 24.960 ;
        RECT 39.225 20.260 39.455 23.560 ;
        RECT 41.515 20.100 41.745 28.420 ;
        RECT 11.115 19.870 20.505 20.100 ;
        RECT 22.015 19.800 30.845 20.100 ;
        RECT 32.355 19.870 41.745 20.100 ;
        RECT 42.975 28.420 52.365 28.650 ;
        RECT 53.875 28.420 62.705 28.720 ;
        RECT 64.215 28.420 73.605 28.650 ;
        RECT 42.975 20.100 43.205 28.420 ;
        RECT 45.265 24.960 45.495 28.260 ;
        RECT 45.230 23.560 45.530 24.960 ;
        RECT 45.265 20.260 45.495 23.560 ;
        RECT 47.555 20.100 47.785 28.420 ;
        RECT 49.845 24.960 50.075 28.260 ;
        RECT 49.810 23.560 50.110 24.960 ;
        RECT 49.845 20.260 50.075 23.560 ;
        RECT 52.135 20.100 52.365 28.420 ;
        RECT 53.595 22.960 53.825 28.260 ;
        RECT 55.885 24.960 56.115 28.260 ;
        RECT 58.175 26.960 58.405 28.260 ;
        RECT 58.140 25.560 58.440 26.960 ;
        RECT 55.850 23.560 56.150 24.960 ;
        RECT 53.560 21.560 53.860 22.960 ;
        RECT 53.595 20.260 53.825 21.560 ;
        RECT 55.885 20.260 56.115 23.560 ;
        RECT 58.175 20.260 58.405 25.560 ;
        RECT 60.465 24.960 60.695 28.260 ;
        RECT 60.430 23.560 60.730 24.960 ;
        RECT 60.465 20.260 60.695 23.560 ;
        RECT 62.755 22.960 62.985 28.260 ;
        RECT 64.215 24.960 64.445 28.420 ;
        RECT 66.505 24.960 66.735 28.260 ;
        RECT 68.795 24.960 69.025 28.420 ;
        RECT 71.085 24.960 71.315 28.260 ;
        RECT 73.375 24.960 73.605 28.420 ;
        RECT 64.180 23.560 64.480 24.960 ;
        RECT 66.470 23.560 66.770 24.960 ;
        RECT 68.760 23.560 69.060 24.960 ;
        RECT 71.050 23.560 71.350 24.960 ;
        RECT 73.340 23.560 73.640 24.960 ;
        RECT 62.720 21.560 63.020 22.960 ;
        RECT 62.755 20.260 62.985 21.560 ;
        RECT 64.215 20.100 64.445 23.560 ;
        RECT 66.505 20.260 66.735 23.560 ;
        RECT 68.795 20.100 69.025 23.560 ;
        RECT 71.085 20.260 71.315 23.560 ;
        RECT 73.375 20.100 73.605 23.560 ;
        RECT 42.975 19.870 52.365 20.100 ;
        RECT 32.635 19.800 41.465 19.870 ;
        RECT 43.255 19.800 52.085 19.870 ;
        RECT 53.875 19.800 62.705 20.100 ;
        RECT 64.215 19.870 73.605 20.100 ;
        RECT 11.115 18.490 20.505 18.720 ;
        RECT 22.015 18.490 30.845 18.790 ;
        RECT 32.635 18.490 41.465 18.790 ;
        RECT 43.255 18.490 52.085 18.790 ;
        RECT 53.875 18.490 62.705 18.790 ;
        RECT 64.215 18.490 73.605 18.720 ;
        RECT 11.115 15.030 11.345 18.490 ;
        RECT 13.405 15.030 13.635 18.330 ;
        RECT 15.695 15.030 15.925 18.490 ;
        RECT 17.985 15.030 18.215 18.330 ;
        RECT 20.275 15.030 20.505 18.490 ;
        RECT 11.020 13.630 11.345 15.030 ;
        RECT 13.370 13.630 13.670 15.030 ;
        RECT 15.660 13.630 15.960 15.030 ;
        RECT 17.950 13.630 18.250 15.030 ;
        RECT 20.240 13.630 20.540 15.030 ;
        RECT 11.115 10.170 11.345 13.630 ;
        RECT 13.405 10.330 13.635 13.630 ;
        RECT 15.695 10.170 15.925 13.630 ;
        RECT 17.985 10.330 18.215 13.630 ;
        RECT 20.275 10.170 20.505 13.630 ;
        RECT 21.735 13.030 21.965 18.330 ;
        RECT 24.025 15.030 24.255 18.330 ;
        RECT 26.315 17.030 26.545 18.330 ;
        RECT 26.280 15.630 26.580 17.030 ;
        RECT 23.990 13.630 24.290 15.030 ;
        RECT 21.700 11.630 22.000 13.030 ;
        RECT 21.735 10.330 21.965 11.630 ;
        RECT 24.025 10.330 24.255 13.630 ;
        RECT 26.315 10.330 26.545 15.630 ;
        RECT 28.605 15.030 28.835 18.330 ;
        RECT 28.570 13.630 28.870 15.030 ;
        RECT 28.605 10.330 28.835 13.630 ;
        RECT 30.895 13.030 31.125 18.330 ;
        RECT 32.355 17.030 32.585 18.330 ;
        RECT 32.320 15.630 32.620 17.030 ;
        RECT 30.860 11.630 31.160 13.030 ;
        RECT 30.895 10.330 31.125 11.630 ;
        RECT 32.355 10.330 32.585 15.630 ;
        RECT 34.645 15.030 34.875 18.330 ;
        RECT 34.610 13.630 34.910 15.030 ;
        RECT 34.645 10.330 34.875 13.630 ;
        RECT 36.935 13.030 37.165 18.330 ;
        RECT 39.225 15.030 39.455 18.330 ;
        RECT 41.515 17.030 41.745 18.330 ;
        RECT 41.480 15.630 41.780 17.030 ;
        RECT 39.190 13.630 39.490 15.030 ;
        RECT 36.900 11.630 37.200 13.030 ;
        RECT 36.935 10.330 37.165 11.630 ;
        RECT 39.225 10.330 39.455 13.630 ;
        RECT 41.515 10.330 41.745 15.630 ;
        RECT 42.975 13.030 43.205 18.330 ;
        RECT 45.265 15.030 45.495 18.330 ;
        RECT 47.555 17.030 47.785 18.330 ;
        RECT 47.520 15.630 47.820 17.030 ;
        RECT 45.230 13.630 45.530 15.030 ;
        RECT 42.940 11.630 43.240 13.030 ;
        RECT 42.975 10.330 43.205 11.630 ;
        RECT 45.265 10.330 45.495 13.630 ;
        RECT 47.555 10.330 47.785 15.630 ;
        RECT 49.845 15.030 50.075 18.330 ;
        RECT 49.810 13.630 50.110 15.030 ;
        RECT 49.845 10.330 50.075 13.630 ;
        RECT 52.135 13.030 52.365 18.330 ;
        RECT 53.595 17.030 53.825 18.330 ;
        RECT 53.560 15.630 53.860 17.030 ;
        RECT 52.100 11.630 52.400 13.030 ;
        RECT 52.135 10.330 52.365 11.630 ;
        RECT 53.595 10.330 53.825 15.630 ;
        RECT 55.885 15.030 56.115 18.330 ;
        RECT 55.850 13.630 56.150 15.030 ;
        RECT 55.885 10.330 56.115 13.630 ;
        RECT 58.175 13.030 58.405 18.330 ;
        RECT 60.465 15.030 60.695 18.330 ;
        RECT 62.755 17.030 62.985 18.330 ;
        RECT 62.720 15.630 63.020 17.030 ;
        RECT 60.430 13.630 60.730 15.030 ;
        RECT 58.140 11.630 58.440 13.030 ;
        RECT 58.175 10.330 58.405 11.630 ;
        RECT 60.465 10.330 60.695 13.630 ;
        RECT 62.755 10.330 62.985 15.630 ;
        RECT 64.215 15.030 64.445 18.490 ;
        RECT 66.505 15.030 66.735 18.330 ;
        RECT 68.795 15.030 69.025 18.490 ;
        RECT 71.085 15.030 71.315 18.330 ;
        RECT 73.375 15.030 73.605 18.490 ;
        RECT 64.180 13.630 64.480 15.030 ;
        RECT 66.470 13.630 66.770 15.030 ;
        RECT 68.760 13.630 69.060 15.030 ;
        RECT 71.050 13.630 71.350 15.030 ;
        RECT 73.340 13.630 73.640 15.030 ;
        RECT 64.215 10.170 64.445 13.630 ;
        RECT 66.505 10.330 66.735 13.630 ;
        RECT 68.795 10.170 69.025 13.630 ;
        RECT 71.085 10.330 71.315 13.630 ;
        RECT 73.375 10.170 73.605 13.630 ;
        RECT 11.115 9.940 20.505 10.170 ;
        RECT 22.015 9.870 30.845 10.170 ;
        RECT 32.635 9.870 41.465 10.170 ;
        RECT 43.255 9.870 52.085 10.170 ;
        RECT 53.875 9.870 62.705 10.170 ;
        RECT 64.215 9.940 73.605 10.170 ;
        RECT 74.105 9.480 80.255 39.040 ;
        RECT 81.035 38.350 82.995 38.580 ;
        RECT 83.325 38.350 85.285 38.580 ;
        RECT 87.075 38.350 89.035 38.700 ;
        RECT 89.365 38.350 91.325 38.700 ;
        RECT 93.115 38.350 97.365 38.700 ;
        RECT 99.155 38.350 101.115 38.700 ;
        RECT 101.445 38.350 103.405 38.700 ;
        RECT 105.195 38.350 107.155 38.700 ;
        RECT 107.485 38.350 109.445 38.700 ;
        RECT 111.235 38.350 115.485 38.700 ;
        RECT 117.275 38.350 119.235 38.700 ;
        RECT 119.565 38.350 121.525 38.700 ;
        RECT 123.315 38.350 125.275 38.580 ;
        RECT 125.605 38.350 127.565 38.580 ;
        RECT 80.755 30.190 80.985 38.190 ;
        RECT 83.045 30.190 83.275 38.190 ;
        RECT 85.335 30.190 85.565 38.190 ;
        RECT 86.795 35.995 87.025 38.190 ;
        RECT 86.560 35.295 87.260 35.995 ;
        RECT 86.795 30.190 87.025 35.295 ;
        RECT 89.085 34.495 89.315 38.190 ;
        RECT 91.375 35.995 91.605 38.190 ;
        RECT 92.835 37.495 93.065 38.190 ;
        RECT 92.600 36.795 93.300 37.495 ;
        RECT 91.140 35.295 91.840 35.995 ;
        RECT 88.850 33.795 89.550 34.495 ;
        RECT 89.085 30.190 89.315 33.795 ;
        RECT 91.375 30.190 91.605 35.295 ;
        RECT 92.835 30.190 93.065 36.795 ;
        RECT 95.125 30.190 95.355 38.350 ;
        RECT 97.415 37.495 97.645 38.190 ;
        RECT 97.180 36.795 97.880 37.495 ;
        RECT 97.415 30.190 97.645 36.795 ;
        RECT 98.875 31.495 99.105 38.190 ;
        RECT 101.165 32.995 101.395 38.190 ;
        RECT 100.930 32.295 101.630 32.995 ;
        RECT 98.640 30.795 99.340 31.495 ;
        RECT 98.875 30.190 99.105 30.795 ;
        RECT 101.165 30.190 101.395 32.295 ;
        RECT 103.455 31.495 103.685 38.190 ;
        RECT 104.915 31.495 105.145 38.190 ;
        RECT 107.205 32.995 107.435 38.190 ;
        RECT 106.970 32.295 107.670 32.995 ;
        RECT 103.220 30.795 103.920 31.495 ;
        RECT 104.680 30.795 105.380 31.495 ;
        RECT 103.455 30.190 103.685 30.795 ;
        RECT 104.915 30.190 105.145 30.795 ;
        RECT 107.205 30.190 107.435 32.295 ;
        RECT 109.495 31.495 109.725 38.190 ;
        RECT 110.955 37.495 111.185 38.190 ;
        RECT 110.720 36.795 111.420 37.495 ;
        RECT 109.260 30.795 109.960 31.495 ;
        RECT 109.495 30.190 109.725 30.795 ;
        RECT 110.955 30.190 111.185 36.795 ;
        RECT 113.245 30.190 113.475 38.350 ;
        RECT 115.535 37.495 115.765 38.190 ;
        RECT 115.300 36.795 116.000 37.495 ;
        RECT 115.535 30.190 115.765 36.795 ;
        RECT 116.995 35.995 117.225 38.190 ;
        RECT 116.760 35.295 117.460 35.995 ;
        RECT 116.995 30.190 117.225 35.295 ;
        RECT 119.285 34.495 119.515 38.190 ;
        RECT 121.575 35.995 121.805 38.190 ;
        RECT 121.340 35.295 122.040 35.995 ;
        RECT 119.050 33.795 119.750 34.495 ;
        RECT 119.285 30.190 119.515 33.795 ;
        RECT 121.575 30.190 121.805 35.295 ;
        RECT 123.035 30.190 123.265 38.190 ;
        RECT 125.325 30.190 125.555 38.190 ;
        RECT 127.615 30.190 127.845 38.190 ;
        RECT 81.035 29.800 82.995 30.030 ;
        RECT 83.325 29.800 85.285 30.030 ;
        RECT 87.075 29.680 89.035 30.030 ;
        RECT 89.365 29.680 91.325 30.030 ;
        RECT 93.115 29.680 95.075 30.030 ;
        RECT 95.405 29.680 97.365 30.030 ;
        RECT 99.155 29.680 101.115 30.030 ;
        RECT 101.445 29.680 103.405 30.030 ;
        RECT 105.195 29.680 107.155 30.030 ;
        RECT 107.485 29.680 109.445 30.030 ;
        RECT 111.235 29.680 113.195 30.030 ;
        RECT 113.525 29.680 115.485 30.030 ;
        RECT 117.275 29.680 119.235 30.030 ;
        RECT 119.565 29.680 121.525 30.030 ;
        RECT 123.315 29.800 125.275 30.030 ;
        RECT 125.605 29.800 127.565 30.030 ;
        RECT 81.035 28.420 82.995 28.650 ;
        RECT 83.325 28.420 85.285 28.650 ;
        RECT 87.075 28.420 89.035 28.770 ;
        RECT 89.365 28.420 91.325 28.770 ;
        RECT 93.115 28.420 95.075 28.770 ;
        RECT 95.405 28.420 97.365 28.770 ;
        RECT 99.155 28.420 101.115 28.770 ;
        RECT 101.445 28.420 103.405 28.770 ;
        RECT 105.195 28.420 107.155 28.770 ;
        RECT 107.485 28.420 109.445 28.770 ;
        RECT 111.235 28.420 113.195 28.770 ;
        RECT 113.525 28.420 115.485 28.770 ;
        RECT 117.275 28.420 119.235 28.770 ;
        RECT 119.565 28.420 121.525 28.770 ;
        RECT 123.315 28.420 125.275 28.650 ;
        RECT 125.605 28.420 127.565 28.650 ;
        RECT 80.755 20.260 80.985 28.260 ;
        RECT 83.045 20.260 83.275 28.260 ;
        RECT 85.335 20.260 85.565 28.260 ;
        RECT 86.795 23.065 87.025 28.260 ;
        RECT 89.085 24.565 89.315 28.260 ;
        RECT 88.850 23.865 89.550 24.565 ;
        RECT 86.560 22.365 87.260 23.065 ;
        RECT 86.795 20.260 87.025 22.365 ;
        RECT 89.085 20.260 89.315 23.865 ;
        RECT 91.375 23.065 91.605 28.260 ;
        RECT 91.140 22.365 91.840 23.065 ;
        RECT 91.375 20.260 91.605 22.365 ;
        RECT 92.835 21.565 93.065 28.260 ;
        RECT 92.600 20.865 93.300 21.565 ;
        RECT 92.835 20.260 93.065 20.865 ;
        RECT 95.125 20.100 95.355 28.260 ;
        RECT 97.415 21.565 97.645 28.260 ;
        RECT 98.875 27.565 99.105 28.260 ;
        RECT 98.640 26.865 99.340 27.565 ;
        RECT 97.180 20.865 97.880 21.565 ;
        RECT 97.415 20.260 97.645 20.865 ;
        RECT 98.875 20.260 99.105 26.865 ;
        RECT 101.165 26.065 101.395 28.260 ;
        RECT 103.455 27.565 103.685 28.260 ;
        RECT 104.915 27.565 105.145 28.260 ;
        RECT 103.220 26.865 103.920 27.565 ;
        RECT 104.680 26.865 105.380 27.565 ;
        RECT 100.930 25.365 101.630 26.065 ;
        RECT 101.165 20.260 101.395 25.365 ;
        RECT 103.455 20.260 103.685 26.865 ;
        RECT 104.915 20.260 105.145 26.865 ;
        RECT 107.205 26.065 107.435 28.260 ;
        RECT 109.495 27.565 109.725 28.260 ;
        RECT 109.260 26.865 109.960 27.565 ;
        RECT 106.970 25.365 107.670 26.065 ;
        RECT 107.205 20.260 107.435 25.365 ;
        RECT 109.495 20.260 109.725 26.865 ;
        RECT 110.955 21.565 111.185 28.260 ;
        RECT 110.720 20.865 111.420 21.565 ;
        RECT 110.955 20.260 111.185 20.865 ;
        RECT 113.245 20.100 113.475 28.260 ;
        RECT 115.535 21.565 115.765 28.260 ;
        RECT 116.995 23.065 117.225 28.260 ;
        RECT 119.285 24.565 119.515 28.260 ;
        RECT 119.050 23.865 119.750 24.565 ;
        RECT 116.760 22.365 117.460 23.065 ;
        RECT 115.300 20.865 116.000 21.565 ;
        RECT 115.535 20.260 115.765 20.865 ;
        RECT 116.995 20.260 117.225 22.365 ;
        RECT 119.285 20.260 119.515 23.865 ;
        RECT 121.575 23.065 121.805 28.260 ;
        RECT 121.340 22.365 122.040 23.065 ;
        RECT 121.575 20.260 121.805 22.365 ;
        RECT 123.035 20.260 123.265 28.260 ;
        RECT 125.325 20.260 125.555 28.260 ;
        RECT 127.615 20.260 127.845 28.260 ;
        RECT 81.035 19.870 82.995 20.100 ;
        RECT 83.325 19.870 85.285 20.100 ;
        RECT 87.075 19.750 89.035 20.100 ;
        RECT 89.365 19.750 91.325 20.100 ;
        RECT 93.115 19.750 97.365 20.100 ;
        RECT 99.155 19.750 101.115 20.100 ;
        RECT 101.445 19.750 103.405 20.100 ;
        RECT 105.195 19.750 107.155 20.100 ;
        RECT 107.485 19.750 109.445 20.100 ;
        RECT 111.235 19.750 115.485 20.100 ;
        RECT 117.275 19.750 119.235 20.100 ;
        RECT 119.565 19.750 121.525 20.100 ;
        RECT 123.315 19.870 125.275 20.100 ;
        RECT 125.605 19.870 127.565 20.100 ;
        RECT 81.035 18.490 82.995 18.720 ;
        RECT 83.325 18.490 85.285 18.720 ;
        RECT 87.075 18.490 89.035 18.720 ;
        RECT 89.365 18.490 91.325 18.720 ;
        RECT 93.115 18.490 95.075 18.720 ;
        RECT 95.405 18.490 97.365 18.720 ;
        RECT 99.155 18.490 101.115 18.720 ;
        RECT 101.445 18.490 103.405 18.720 ;
        RECT 105.195 18.490 107.155 18.720 ;
        RECT 107.485 18.490 109.445 18.720 ;
        RECT 111.235 18.490 113.195 18.720 ;
        RECT 113.525 18.490 115.485 18.720 ;
        RECT 117.275 18.490 119.235 18.720 ;
        RECT 119.565 18.490 121.525 18.720 ;
        RECT 123.315 18.490 125.275 18.720 ;
        RECT 125.605 18.490 127.565 18.720 ;
        RECT 80.755 10.330 80.985 18.330 ;
        RECT 83.045 10.330 83.275 18.330 ;
        RECT 85.335 10.330 85.565 18.330 ;
        RECT 86.795 10.330 87.025 18.330 ;
        RECT 89.085 10.330 89.315 18.330 ;
        RECT 91.375 10.330 91.605 18.330 ;
        RECT 92.835 10.330 93.065 18.330 ;
        RECT 95.125 10.330 95.355 18.330 ;
        RECT 97.415 10.330 97.645 18.330 ;
        RECT 98.875 10.330 99.105 18.330 ;
        RECT 101.165 10.330 101.395 18.330 ;
        RECT 103.455 10.330 103.685 18.330 ;
        RECT 104.915 10.330 105.145 18.330 ;
        RECT 107.205 10.330 107.435 18.330 ;
        RECT 109.495 10.330 109.725 18.330 ;
        RECT 110.955 10.330 111.185 18.330 ;
        RECT 113.245 10.330 113.475 18.330 ;
        RECT 115.535 10.330 115.765 18.330 ;
        RECT 116.995 10.330 117.225 18.330 ;
        RECT 119.285 10.330 119.515 18.330 ;
        RECT 121.575 10.330 121.805 18.330 ;
        RECT 123.035 10.330 123.265 18.330 ;
        RECT 125.325 10.330 125.555 18.330 ;
        RECT 127.615 10.330 127.845 18.330 ;
        RECT 81.035 9.940 82.995 10.170 ;
        RECT 83.325 9.940 85.285 10.170 ;
        RECT 87.075 9.940 89.035 10.170 ;
        RECT 89.365 9.940 91.325 10.170 ;
        RECT 93.115 9.940 95.075 10.170 ;
        RECT 95.405 9.940 97.365 10.170 ;
        RECT 99.155 9.940 101.115 10.170 ;
        RECT 101.445 9.940 103.405 10.170 ;
        RECT 105.195 9.940 107.155 10.170 ;
        RECT 107.485 9.940 109.445 10.170 ;
        RECT 111.235 9.940 113.195 10.170 ;
        RECT 113.525 9.940 115.485 10.170 ;
        RECT 117.275 9.940 119.235 10.170 ;
        RECT 119.565 9.940 121.525 10.170 ;
        RECT 123.315 9.940 125.275 10.170 ;
        RECT 125.605 9.940 127.565 10.170 ;
        RECT 128.345 9.480 130.565 39.040 ;
        RECT 8.665 8.890 130.565 9.480 ;
        RECT 7.065 5.690 130.565 8.890 ;
        RECT 135.120 18.845 135.710 41.635 ;
        RECT 136.295 40.485 138.400 41.075 ;
        RECT 136.295 39.315 138.400 39.905 ;
        RECT 146.290 39.315 148.395 41.075 ;
        RECT 136.295 36.975 138.400 38.735 ;
        RECT 146.290 38.145 148.395 38.735 ;
        RECT 146.290 36.975 148.395 37.565 ;
        RECT 136.295 35.805 138.400 36.395 ;
        RECT 136.295 34.635 138.400 35.225 ;
        RECT 146.290 34.635 148.395 36.395 ;
        RECT 136.295 32.295 138.400 34.055 ;
        RECT 146.290 33.465 148.395 34.055 ;
        RECT 143.640 32.295 148.395 32.885 ;
        RECT 136.295 31.125 138.400 31.715 ;
        RECT 136.295 29.955 141.055 30.545 ;
        RECT 146.290 29.955 148.395 31.715 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 136.295 26.445 138.400 28.205 ;
        RECT 146.290 27.615 148.395 29.375 ;
        RECT 136.295 24.105 138.400 25.865 ;
        RECT 146.290 25.275 148.395 27.035 ;
        RECT 136.295 21.765 138.400 23.525 ;
        RECT 146.290 22.935 148.395 24.695 ;
        RECT 136.295 19.425 138.400 21.185 ;
        RECT 146.290 20.595 148.395 22.355 ;
        RECT 141.295 19.425 148.395 20.015 ;
        RECT 148.980 18.845 155.900 104.835 ;
        RECT 135.120 14.050 138.400 18.845 ;
        RECT 146.290 14.050 155.900 18.845 ;
        RECT 135.120 4.900 155.900 14.050 ;
        RECT 4.100 4.100 155.900 4.900 ;
      LAYER met2 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.495 208.765 51.905 210.765 ;
        RECT 9.495 205.765 45.165 207.765 ;
        RECT 51.315 207.460 51.905 208.765 ;
        RECT 9.495 202.765 48.270 204.765 ;
        RECT 9.495 198.745 48.270 200.745 ;
        RECT 9.495 195.745 45.165 197.745 ;
        RECT 9.495 192.745 46.670 194.745 ;
        RECT 9.495 187.420 15.245 188.980 ;
        RECT 16.515 188.295 45.165 190.295 ;
        RECT 52.860 188.465 54.245 190.570 ;
        RECT 16.515 184.775 56.920 186.775 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.495 182.570 15.245 184.130 ;
        RECT 16.515 181.255 46.670 183.255 ;
        RECT 5.910 176.050 7.510 179.250 ;
        RECT 57.020 178.865 57.820 178.990 ;
        RECT 9.500 177.365 58.420 178.865 ;
        RECT 53.870 176.720 54.670 176.890 ;
        RECT 9.500 175.220 54.670 176.720 ;
        RECT 9.500 172.820 54.670 174.320 ;
        RECT 53.870 172.640 54.670 172.820 ;
        RECT 52.220 171.920 53.020 172.040 ;
        RECT 9.500 170.420 53.020 171.920 ;
        RECT 63.470 170.855 65.220 217.105 ;
        RECT 66.220 170.855 67.970 217.105 ;
        RECT 68.970 170.855 70.720 217.105 ;
        RECT 71.720 170.855 73.470 217.105 ;
        RECT 74.470 170.855 76.220 217.105 ;
        RECT 77.220 170.855 78.970 217.105 ;
        RECT 79.970 170.115 81.970 217.845 ;
        RECT 106.340 217.515 107.940 220.715 ;
        RECT 109.240 219.705 111.675 220.105 ;
        RECT 113.270 219.705 115.705 220.105 ;
        RECT 117.300 219.705 119.735 220.105 ;
        RECT 121.330 219.705 123.765 220.105 ;
        RECT 125.360 219.705 127.795 220.105 ;
        RECT 129.390 219.705 131.825 220.105 ;
        RECT 133.420 219.705 135.855 220.105 ;
        RECT 137.450 219.705 139.885 220.105 ;
        RECT 141.480 219.705 143.915 220.105 ;
        RECT 145.510 219.705 147.945 220.105 ;
        RECT 149.540 219.705 151.975 220.105 ;
        RECT 109.240 217.705 109.640 219.705 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 111.820 217.295 112.220 219.305 ;
        RECT 113.270 217.705 113.670 219.705 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 115.850 217.295 116.250 219.305 ;
        RECT 117.300 217.705 117.700 219.705 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 119.880 217.295 120.280 219.305 ;
        RECT 121.330 217.705 121.730 219.705 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 123.910 217.295 124.310 219.305 ;
        RECT 125.360 217.705 125.760 219.705 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 127.940 217.295 128.340 219.305 ;
        RECT 129.390 217.705 129.790 219.705 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 131.970 217.295 132.370 219.305 ;
        RECT 133.420 217.705 133.820 219.705 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 136.000 217.295 136.400 219.305 ;
        RECT 137.450 217.705 137.850 219.705 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 140.030 217.295 140.430 219.305 ;
        RECT 141.480 217.705 141.880 219.705 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 144.060 217.295 144.460 219.305 ;
        RECT 145.510 217.705 145.910 219.705 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 148.090 217.295 148.490 219.305 ;
        RECT 149.540 217.705 149.940 219.705 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 152.120 217.295 152.520 219.305 ;
        RECT 82.970 170.855 84.720 217.105 ;
        RECT 85.720 170.855 87.470 217.105 ;
        RECT 88.470 170.855 90.220 217.105 ;
        RECT 91.220 170.855 92.970 217.105 ;
        RECT 93.970 170.855 95.720 217.105 ;
        RECT 96.720 170.855 98.470 217.105 ;
        RECT 109.785 216.895 112.220 217.295 ;
        RECT 113.815 216.895 116.250 217.295 ;
        RECT 117.845 216.895 120.280 217.295 ;
        RECT 121.875 216.895 124.310 217.295 ;
        RECT 125.905 216.895 128.340 217.295 ;
        RECT 129.935 216.895 132.370 217.295 ;
        RECT 133.965 216.895 136.400 217.295 ;
        RECT 137.995 216.895 140.430 217.295 ;
        RECT 142.025 216.895 144.460 217.295 ;
        RECT 146.055 216.895 148.490 217.295 ;
        RECT 150.085 216.895 152.520 217.295 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 111.820 205.955 112.220 206.755 ;
        RECT 115.850 205.955 116.250 206.755 ;
        RECT 119.880 205.955 120.280 206.755 ;
        RECT 123.910 205.955 124.310 206.755 ;
        RECT 127.940 205.955 128.340 206.755 ;
        RECT 131.970 205.955 132.370 206.755 ;
        RECT 136.000 205.955 136.400 206.755 ;
        RECT 140.030 205.955 140.430 206.755 ;
        RECT 144.060 205.955 144.460 206.755 ;
        RECT 148.090 205.955 148.490 206.755 ;
        RECT 152.120 205.955 152.520 206.755 ;
        RECT 109.240 204.745 111.675 205.545 ;
        RECT 113.270 204.745 115.705 205.545 ;
        RECT 117.300 204.745 119.735 205.545 ;
        RECT 121.330 204.745 123.765 205.545 ;
        RECT 125.360 204.745 127.795 205.545 ;
        RECT 129.390 204.745 131.825 205.545 ;
        RECT 133.420 204.745 135.855 205.545 ;
        RECT 137.450 204.745 139.885 205.545 ;
        RECT 141.480 204.745 143.915 205.545 ;
        RECT 145.510 204.745 147.945 205.545 ;
        RECT 149.540 204.745 151.975 205.545 ;
        RECT 108.540 202.425 108.940 202.625 ;
        RECT 109.785 202.425 110.385 204.345 ;
        RECT 108.540 202.025 110.385 202.425 ;
        RECT 108.540 201.825 108.940 202.025 ;
        RECT 109.785 199.970 110.385 202.025 ;
        RECT 111.075 199.970 111.675 204.745 ;
        RECT 112.570 202.425 112.970 202.625 ;
        RECT 113.815 202.425 114.415 204.345 ;
        RECT 112.570 202.025 114.415 202.425 ;
        RECT 112.570 201.825 112.970 202.025 ;
        RECT 113.815 199.970 114.415 202.025 ;
        RECT 115.105 199.970 115.705 204.745 ;
        RECT 116.600 202.425 117.000 202.625 ;
        RECT 117.845 202.425 118.445 204.345 ;
        RECT 116.600 202.025 118.445 202.425 ;
        RECT 116.600 201.825 117.000 202.025 ;
        RECT 117.845 199.970 118.445 202.025 ;
        RECT 119.135 199.970 119.735 204.745 ;
        RECT 120.630 202.425 121.030 202.625 ;
        RECT 121.875 202.425 122.475 204.345 ;
        RECT 120.630 202.025 122.475 202.425 ;
        RECT 120.630 201.825 121.030 202.025 ;
        RECT 121.875 199.970 122.475 202.025 ;
        RECT 123.165 199.970 123.765 204.745 ;
        RECT 124.660 202.425 125.060 202.625 ;
        RECT 125.905 202.425 126.505 204.345 ;
        RECT 124.660 202.025 126.505 202.425 ;
        RECT 124.660 201.825 125.060 202.025 ;
        RECT 125.905 199.970 126.505 202.025 ;
        RECT 127.195 199.970 127.795 204.745 ;
        RECT 128.690 202.425 129.090 202.625 ;
        RECT 129.935 202.425 130.535 204.345 ;
        RECT 128.690 202.025 130.535 202.425 ;
        RECT 128.690 201.825 129.090 202.025 ;
        RECT 129.935 199.970 130.535 202.025 ;
        RECT 131.225 199.970 131.825 204.745 ;
        RECT 132.720 202.425 133.120 202.625 ;
        RECT 133.965 202.425 134.565 204.345 ;
        RECT 132.720 202.025 134.565 202.425 ;
        RECT 132.720 201.825 133.120 202.025 ;
        RECT 133.965 199.970 134.565 202.025 ;
        RECT 135.255 199.970 135.855 204.745 ;
        RECT 136.750 202.425 137.150 202.625 ;
        RECT 137.995 202.425 138.595 204.345 ;
        RECT 136.750 202.025 138.595 202.425 ;
        RECT 136.750 201.825 137.150 202.025 ;
        RECT 137.995 199.970 138.595 202.025 ;
        RECT 139.285 199.970 139.885 204.745 ;
        RECT 140.780 202.425 141.180 202.625 ;
        RECT 142.025 202.425 142.625 204.345 ;
        RECT 140.780 202.025 142.625 202.425 ;
        RECT 140.780 201.825 141.180 202.025 ;
        RECT 142.025 199.970 142.625 202.025 ;
        RECT 143.315 199.970 143.915 204.745 ;
        RECT 144.810 202.425 145.210 202.625 ;
        RECT 146.055 202.425 146.655 204.345 ;
        RECT 144.810 202.025 146.655 202.425 ;
        RECT 144.810 201.825 145.210 202.025 ;
        RECT 146.055 199.970 146.655 202.025 ;
        RECT 147.345 199.970 147.945 204.745 ;
        RECT 148.840 202.425 149.240 202.625 ;
        RECT 150.085 202.425 150.685 204.345 ;
        RECT 148.840 202.025 150.685 202.425 ;
        RECT 148.840 201.825 149.240 202.025 ;
        RECT 150.085 199.970 150.685 202.025 ;
        RECT 151.375 199.970 151.975 204.745 ;
        RECT 109.240 194.440 109.640 199.685 ;
        RECT 109.240 194.040 110.255 194.440 ;
        RECT 109.240 191.285 109.640 192.885 ;
        RECT 110.530 187.540 110.930 198.905 ;
        RECT 111.820 194.440 112.220 199.685 ;
        RECT 111.205 194.040 112.220 194.440 ;
        RECT 113.270 194.440 113.670 199.685 ;
        RECT 113.270 194.040 114.285 194.440 ;
        RECT 111.820 191.285 112.220 192.885 ;
        RECT 113.270 191.285 113.670 192.885 ;
        RECT 114.560 187.540 114.960 198.905 ;
        RECT 115.850 194.440 116.250 199.685 ;
        RECT 115.235 194.040 116.250 194.440 ;
        RECT 117.300 194.440 117.700 199.685 ;
        RECT 117.300 194.040 118.315 194.440 ;
        RECT 115.850 191.285 116.250 192.885 ;
        RECT 117.300 191.285 117.700 192.885 ;
        RECT 118.590 187.540 118.990 198.905 ;
        RECT 119.880 194.440 120.280 199.685 ;
        RECT 119.265 194.040 120.280 194.440 ;
        RECT 121.330 194.440 121.730 199.685 ;
        RECT 121.330 194.040 122.345 194.440 ;
        RECT 119.880 191.285 120.280 192.885 ;
        RECT 121.330 191.285 121.730 192.885 ;
        RECT 122.620 187.540 123.020 198.905 ;
        RECT 123.910 194.440 124.310 199.685 ;
        RECT 123.295 194.040 124.310 194.440 ;
        RECT 125.360 194.440 125.760 199.685 ;
        RECT 125.360 194.040 126.375 194.440 ;
        RECT 123.910 191.285 124.310 192.885 ;
        RECT 125.360 191.285 125.760 192.885 ;
        RECT 126.650 187.540 127.050 198.905 ;
        RECT 127.940 194.440 128.340 199.685 ;
        RECT 127.325 194.040 128.340 194.440 ;
        RECT 129.390 194.440 129.790 199.685 ;
        RECT 129.390 194.040 130.405 194.440 ;
        RECT 127.940 191.285 128.340 192.885 ;
        RECT 129.390 191.285 129.790 192.885 ;
        RECT 130.680 187.540 131.080 198.905 ;
        RECT 131.970 194.440 132.370 199.685 ;
        RECT 131.355 194.040 132.370 194.440 ;
        RECT 133.420 194.440 133.820 199.685 ;
        RECT 133.420 194.040 134.435 194.440 ;
        RECT 131.970 191.285 132.370 192.885 ;
        RECT 133.420 191.285 133.820 192.885 ;
        RECT 134.710 187.540 135.110 198.905 ;
        RECT 136.000 194.440 136.400 199.685 ;
        RECT 135.385 194.040 136.400 194.440 ;
        RECT 137.450 194.440 137.850 199.685 ;
        RECT 137.450 194.040 138.465 194.440 ;
        RECT 136.000 191.285 136.400 192.885 ;
        RECT 137.450 191.285 137.850 192.885 ;
        RECT 138.740 187.540 139.140 198.905 ;
        RECT 140.030 194.440 140.430 199.685 ;
        RECT 139.415 194.040 140.430 194.440 ;
        RECT 141.480 194.440 141.880 199.685 ;
        RECT 141.480 194.040 142.495 194.440 ;
        RECT 140.030 191.285 140.430 192.885 ;
        RECT 141.480 191.285 141.880 192.885 ;
        RECT 142.770 187.540 143.170 198.905 ;
        RECT 144.060 194.440 144.460 199.685 ;
        RECT 143.445 194.040 144.460 194.440 ;
        RECT 145.510 194.440 145.910 199.685 ;
        RECT 145.510 194.040 146.525 194.440 ;
        RECT 144.060 191.285 144.460 192.885 ;
        RECT 145.510 191.285 145.910 192.885 ;
        RECT 146.800 187.540 147.200 198.905 ;
        RECT 148.090 194.440 148.490 199.685 ;
        RECT 147.475 194.040 148.490 194.440 ;
        RECT 149.540 194.440 149.940 199.685 ;
        RECT 149.540 194.040 150.555 194.440 ;
        RECT 148.090 191.285 148.490 192.885 ;
        RECT 149.540 191.285 149.940 192.885 ;
        RECT 150.830 187.540 151.230 198.905 ;
        RECT 152.120 194.440 152.520 199.685 ;
        RECT 151.505 194.040 152.520 194.440 ;
        RECT 152.120 191.285 152.520 192.885 ;
        RECT 109.240 184.370 109.640 184.770 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 109.240 183.970 154.345 184.370 ;
        RECT 153.945 183.570 154.345 183.970 ;
        RECT 115.265 175.815 117.965 176.215 ;
        RECT 119.885 175.815 122.585 176.215 ;
        RECT 124.505 175.815 127.205 176.215 ;
        RECT 129.125 175.815 131.825 176.215 ;
        RECT 133.745 175.815 136.445 176.215 ;
        RECT 138.365 175.815 141.065 176.215 ;
        RECT 142.985 175.815 145.685 176.215 ;
        RECT 147.605 175.815 150.305 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 114.835 172.120 118.395 174.820 ;
        RECT 119.155 172.120 123.015 174.820 ;
        RECT 123.775 172.120 127.635 174.820 ;
        RECT 128.395 172.120 132.255 174.820 ;
        RECT 133.015 172.120 136.875 174.820 ;
        RECT 137.635 172.120 141.495 174.820 ;
        RECT 142.255 172.120 146.115 174.820 ;
        RECT 146.875 172.120 150.735 174.820 ;
        RECT 57.020 169.775 57.820 169.890 ;
        RECT 9.500 168.275 58.420 169.775 ;
        RECT 9.500 165.715 56.920 166.715 ;
        RECT 103.350 164.990 103.750 170.890 ;
        RECT 105.930 168.490 106.330 170.890 ;
        RECT 9.500 163.915 55.070 164.915 ;
        RECT 102.625 164.590 103.750 164.990 ;
        RECT 104.640 164.790 105.040 167.190 ;
        RECT 107.380 164.990 107.780 170.890 ;
        RECT 109.960 168.490 110.360 170.890 ;
        RECT 115.625 169.795 117.605 170.845 ;
        RECT 119.155 169.795 119.755 172.120 ;
        RECT 115.625 169.195 119.755 169.795 ;
        RECT 120.245 169.795 122.225 170.845 ;
        RECT 123.775 169.795 124.375 172.120 ;
        RECT 120.245 169.195 124.375 169.795 ;
        RECT 124.865 169.795 126.845 170.845 ;
        RECT 128.395 169.795 128.995 172.120 ;
        RECT 124.865 169.195 128.995 169.795 ;
        RECT 129.485 169.795 131.465 170.845 ;
        RECT 133.015 169.795 133.615 172.120 ;
        RECT 129.485 169.195 133.615 169.795 ;
        RECT 134.105 169.795 136.085 170.845 ;
        RECT 137.635 169.795 138.235 172.120 ;
        RECT 134.105 169.195 138.235 169.795 ;
        RECT 138.725 169.795 140.705 170.845 ;
        RECT 142.255 169.795 142.855 172.120 ;
        RECT 138.725 169.195 142.855 169.795 ;
        RECT 143.345 169.795 145.325 170.845 ;
        RECT 146.875 169.795 147.475 172.120 ;
        RECT 143.345 169.195 147.475 169.795 ;
        RECT 115.625 168.145 117.605 169.195 ;
        RECT 120.245 168.145 122.225 169.195 ;
        RECT 124.865 168.145 126.845 169.195 ;
        RECT 129.485 168.145 131.465 169.195 ;
        RECT 134.105 168.145 136.085 169.195 ;
        RECT 138.725 168.145 140.705 169.195 ;
        RECT 143.345 168.145 145.325 169.195 ;
        RECT 147.965 168.145 150.345 170.845 ;
        RECT 106.655 164.590 107.780 164.990 ;
        RECT 108.670 164.790 109.070 167.190 ;
        RECT 9.500 162.115 51.610 163.115 ;
        RECT 9.500 159.815 53.170 161.315 ;
        RECT 2.705 157.015 51.610 159.015 ;
        RECT 2.705 1.285 3.505 157.015 ;
        RECT 9.500 154.715 53.170 156.215 ;
        RECT 9.500 152.915 51.610 153.915 ;
        RECT 9.500 151.115 55.070 152.115 ;
        RECT 74.940 151.875 86.100 155.595 ;
        RECT 9.500 149.315 56.520 150.315 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 148.155 78.660 151.875 ;
        RECT 80.100 149.595 80.930 150.425 ;
        RECT 82.380 148.155 86.100 151.875 ;
        RECT 102.625 149.850 103.025 164.590 ;
        RECT 103.350 162.940 104.365 163.340 ;
        RECT 105.315 162.940 106.330 163.340 ;
        RECT 103.350 159.695 103.750 162.940 ;
        RECT 105.930 160.395 106.330 162.940 ;
        RECT 104.190 159.795 106.330 160.395 ;
        RECT 104.190 159.410 104.495 159.795 ;
        RECT 105.930 159.695 106.330 159.795 ;
        RECT 103.895 154.535 104.495 159.410 ;
        RECT 105.185 155.035 105.785 159.410 ;
        RECT 103.895 153.935 106.330 154.535 ;
        RECT 103.350 150.640 103.750 153.565 ;
        RECT 105.930 152.190 106.330 153.935 ;
        RECT 103.895 151.790 106.330 152.190 ;
        RECT 103.895 151.015 104.495 151.790 ;
        RECT 105.185 150.640 105.785 151.415 ;
        RECT 103.350 150.240 105.785 150.640 ;
        RECT 106.655 149.850 107.055 164.590 ;
        RECT 107.380 162.940 108.395 163.340 ;
        RECT 109.345 162.940 110.360 163.340 ;
        RECT 107.380 159.695 107.780 162.940 ;
        RECT 109.960 160.395 110.360 162.940 ;
        RECT 108.220 159.795 110.360 160.395 ;
        RECT 108.220 159.410 108.525 159.795 ;
        RECT 109.960 159.695 110.360 159.795 ;
        RECT 107.925 154.535 108.525 159.410 ;
        RECT 109.215 155.035 109.815 159.410 ;
        RECT 107.925 153.935 110.360 154.535 ;
        RECT 107.380 150.640 107.780 153.565 ;
        RECT 109.960 152.190 110.360 153.935 ;
        RECT 107.925 151.790 110.360 152.190 ;
        RECT 107.925 151.015 108.525 151.790 ;
        RECT 109.215 150.640 109.815 151.415 ;
        RECT 107.380 150.240 109.815 150.640 ;
        RECT 102.625 149.450 103.750 149.850 ;
        RECT 74.940 144.435 86.100 148.155 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 11.195 139.800 23.015 140.200 ;
        RECT 11.195 137.185 11.795 139.800 ;
        RECT 14.860 138.370 21.050 138.770 ;
        RECT 14.860 137.585 15.260 138.370 ;
        RECT 20.650 137.970 21.050 138.370 ;
        RECT 14.130 137.185 16.020 137.585 ;
        RECT 16.805 137.185 18.955 137.585 ;
        RECT 16.805 136.875 17.205 137.185 ;
        RECT 11.940 136.275 15.275 136.875 ;
        RECT 16.165 136.275 17.205 136.875 ;
        RECT 5.910 132.225 7.510 135.425 ;
        RECT 13.485 133.130 14.085 135.875 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 16.805 129.110 17.205 136.275 ;
        RECT 19.100 136.125 20.750 136.725 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 19.100 128.925 19.500 136.125 ;
        RECT 22.615 134.120 23.015 139.800 ;
        RECT 24.255 135.155 25.755 143.745 ;
        RECT 27.765 135.155 29.265 143.745 ;
        RECT 36.055 135.155 37.555 143.745 ;
        RECT 44.345 135.155 45.845 143.745 ;
        RECT 52.635 135.155 54.135 143.745 ;
        RECT 56.145 135.155 57.645 143.745 ;
        RECT 103.350 143.435 103.750 149.450 ;
        RECT 104.640 147.135 105.040 149.535 ;
        RECT 106.655 149.450 107.780 149.850 ;
        RECT 105.930 143.435 106.330 145.835 ;
        RECT 107.380 143.435 107.780 149.450 ;
        RECT 108.670 147.135 109.070 149.535 ;
        RECT 109.960 143.435 110.360 145.835 ;
        RECT 116.310 143.410 116.910 168.145 ;
        RECT 120.930 147.550 121.530 168.145 ;
        RECT 125.550 159.440 126.150 168.145 ;
        RECT 125.550 158.840 128.940 159.440 ;
        RECT 120.930 146.950 126.935 147.550 ;
        RECT 122.645 144.030 124.245 144.830 ;
        RECT 128.340 144.540 128.940 158.840 ;
        RECT 130.170 148.610 130.770 168.145 ;
        RECT 134.795 164.330 135.395 168.145 ;
        RECT 133.685 163.140 134.485 163.740 ;
        RECT 133.785 155.610 134.385 163.140 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 139.410 157.075 140.010 168.145 ;
        RECT 144.035 163.040 144.635 168.145 ;
        RECT 146.855 164.430 147.655 165.030 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 141.615 158.550 142.415 159.150 ;
        RECT 138.070 156.475 140.010 157.075 ;
        RECT 133.285 155.010 134.885 155.610 ;
        RECT 133.275 151.400 134.875 152.200 ;
        RECT 133.275 150.230 134.875 151.030 ;
        RECT 138.070 149.760 138.670 156.475 ;
        RECT 141.715 152.110 142.315 158.550 ;
        RECT 141.215 151.905 142.815 152.110 ;
        RECT 140.950 151.505 143.050 151.905 ;
        RECT 133.285 149.160 138.670 149.760 ;
        RECT 130.170 148.010 134.430 148.610 ;
        RECT 130.615 146.830 132.215 147.630 ;
        RECT 133.285 147.410 134.885 148.010 ;
        RECT 138.525 147.310 140.125 148.110 ;
        RECT 128.340 143.940 134.885 144.540 ;
        RECT 138.525 143.820 140.125 144.620 ;
        RECT 116.310 142.810 132.215 143.410 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 141.990 142.815 142.790 ;
        RECT 146.955 142.730 147.555 164.430 ;
        RECT 148.655 158.450 149.255 168.145 ;
        RECT 146.455 142.640 148.055 142.730 ;
        RECT 146.195 142.240 148.295 142.640 ;
        RECT 146.455 142.130 148.055 142.240 ;
        RECT 104.640 139.365 152.360 140.165 ;
        RECT 97.200 137.420 147.750 138.220 ;
        RECT 107.380 135.525 132.465 136.325 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 56.145 133.555 77.110 135.155 ;
        RECT 80.120 133.320 137.265 134.120 ;
        RECT 137.945 133.410 144.375 133.810 ;
        RECT 21.615 131.745 135.665 132.545 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 142.980 131.990 143.630 132.590 ;
        RECT 27.065 129.995 134.065 130.795 ;
        RECT 19.100 128.125 101.315 128.925 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 142.980 126.815 143.230 131.990 ;
        RECT 144.025 131.050 144.375 133.410 ;
        RECT 143.725 129.545 144.425 131.050 ;
        RECT 153.945 129.545 154.345 129.945 ;
        RECT 143.725 129.145 154.345 129.545 ;
        RECT 143.725 127.640 144.425 129.145 ;
        RECT 142.980 126.215 143.630 126.815 ;
        RECT 10.025 122.800 70.175 123.810 ;
        RECT 71.775 122.750 114.165 123.850 ;
        RECT 10.025 120.300 70.175 122.300 ;
        RECT 71.775 121.250 114.165 122.350 ;
        RECT 115.905 121.575 128.935 123.145 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 10.025 117.800 70.175 119.800 ;
        RECT 71.775 119.750 114.165 120.850 ;
        RECT 71.775 118.250 114.165 119.350 ;
        RECT 10.025 115.300 70.175 117.300 ;
        RECT 71.775 116.750 114.165 117.850 ;
        RECT 115.905 117.075 128.935 118.645 ;
        RECT 141.900 116.370 150.745 117.170 ;
        RECT 71.775 115.250 114.165 116.350 ;
        RECT 10.025 112.780 70.175 114.800 ;
        RECT 71.775 112.730 114.165 114.850 ;
        RECT 136.465 114.770 144.870 115.570 ;
        RECT 115.905 112.615 128.935 114.185 ;
        RECT 10.025 110.280 70.175 112.280 ;
        RECT 71.775 111.230 114.165 112.330 ;
        RECT 133.265 111.795 141.675 112.595 ;
        RECT 10.025 107.780 70.175 109.780 ;
        RECT 71.775 109.730 114.165 110.830 ;
        RECT 140.875 110.315 141.675 111.795 ;
        RECT 144.070 110.315 144.870 114.770 ;
        RECT 71.775 108.230 114.165 109.330 ;
        RECT 115.905 108.115 128.935 109.685 ;
        RECT 139.560 109.515 142.995 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 10.025 105.280 70.175 107.280 ;
        RECT 71.775 106.730 114.165 107.830 ;
        RECT 71.775 105.230 114.165 106.330 ;
        RECT 10.025 103.770 70.175 104.780 ;
        RECT 71.775 103.730 114.165 104.830 ;
        RECT 115.905 103.655 128.935 105.225 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 10.025 91.525 128.935 92.775 ;
        RECT 10.025 89.640 128.935 91.140 ;
        RECT 10.025 85.640 128.935 88.640 ;
        RECT 136.295 86.115 138.400 90.215 ;
        RECT 10.025 83.140 128.935 84.640 ;
        RECT 10.025 81.505 128.935 82.755 ;
        RECT 10.025 79.620 128.935 81.120 ;
        RECT 136.295 80.265 138.400 85.535 ;
        RECT 139.560 82.025 140.860 109.515 ;
        RECT 141.695 91.385 142.995 109.515 ;
        RECT 141.290 90.795 143.395 91.385 ;
        RECT 139.155 81.435 141.260 82.025 ;
        RECT 10.025 75.620 128.935 78.620 ;
        RECT 136.295 75.585 138.400 79.685 ;
        RECT 10.025 73.120 128.935 74.620 ;
        RECT 10.025 71.485 128.935 72.735 ;
        RECT 10.025 69.600 128.935 71.100 ;
        RECT 136.295 70.905 138.400 75.005 ;
        RECT 10.025 65.600 128.935 68.600 ;
        RECT 136.295 66.225 138.400 70.325 ;
        RECT 10.025 63.100 128.935 64.600 ;
        RECT 10.025 61.465 128.935 62.715 ;
        RECT 10.025 59.580 128.935 61.080 ;
        RECT 136.295 60.375 138.400 65.645 ;
        RECT 10.025 55.580 128.935 58.580 ;
        RECT 136.295 55.695 138.400 59.795 ;
        RECT 10.025 53.080 128.935 54.580 ;
        RECT 10.025 51.445 128.935 52.695 ;
        RECT 136.295 51.015 138.400 55.115 ;
        RECT 12.915 45.565 14.515 47.165 ;
        RECT 90.715 45.565 92.315 47.165 ;
        RECT 136.295 46.335 138.400 50.435 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 136.295 40.485 138.400 45.755 ;
        RECT 143.835 42.245 145.135 110.315 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 146.290 88.455 148.395 92.555 ;
        RECT 146.290 83.775 148.395 87.875 ;
        RECT 146.290 77.925 148.395 83.195 ;
        RECT 146.290 73.245 148.395 77.345 ;
        RECT 146.290 68.565 148.395 72.665 ;
        RECT 146.290 63.885 148.395 67.985 ;
        RECT 146.290 58.035 148.395 63.305 ;
        RECT 146.290 53.355 148.395 57.455 ;
        RECT 146.290 48.675 148.395 52.775 ;
        RECT 146.290 43.995 148.395 48.095 ;
        RECT 143.435 41.655 145.540 42.245 ;
        RECT 143.835 41.605 145.135 41.655 ;
        RECT 7.065 36.430 8.665 39.630 ;
        RECT 10.170 37.965 74.550 38.965 ;
        RECT 79.810 38.185 127.975 39.285 ;
        RECT 10.170 35.440 74.550 36.940 ;
        RECT 79.810 36.685 127.975 37.785 ;
        RECT 79.810 35.185 127.975 36.285 ;
        RECT 136.295 35.805 138.400 39.905 ;
        RECT 146.290 38.145 148.395 43.415 ;
        RECT 10.170 33.440 74.550 34.940 ;
        RECT 79.810 33.685 127.975 34.785 ;
        RECT 10.170 31.440 74.550 32.940 ;
        RECT 79.810 32.185 127.975 33.285 ;
        RECT 79.810 30.685 127.975 31.785 ;
        RECT 136.295 31.125 138.400 35.225 ;
        RECT 146.290 33.465 148.395 37.565 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 10.170 28.035 74.550 30.415 ;
        RECT 79.810 28.165 127.975 30.285 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 10.170 25.510 74.550 27.010 ;
        RECT 79.810 26.665 127.975 27.765 ;
        RECT 79.810 25.165 127.975 26.265 ;
        RECT 10.170 23.510 74.550 25.010 ;
        RECT 79.810 23.665 127.975 24.765 ;
        RECT 10.170 21.510 74.550 23.010 ;
        RECT 79.810 22.165 127.975 23.265 ;
        RECT 79.810 20.665 127.975 21.765 ;
        RECT 10.170 18.105 74.550 20.485 ;
        RECT 79.810 19.165 127.975 20.265 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 10.170 15.580 74.550 17.080 ;
        RECT 10.170 13.580 74.550 15.080 ;
        RECT 10.170 11.580 74.550 13.080 ;
        RECT 10.170 9.555 74.550 10.555 ;
        RECT 80.745 9.665 82.345 10.465 ;
        RECT 7.065 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.965 5.690 130.565 8.890 ;
      LAYER met3 ;
        RECT 108.865 224.515 109.665 224.615 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.915 106.460 224.450 ;
        RECT 108.865 224.215 129.040 224.515 ;
        RECT 95.070 221.515 95.370 223.650 ;
        RECT 97.830 222.115 98.130 223.650 ;
        RECT 100.590 222.715 100.890 223.650 ;
        RECT 103.350 223.315 103.650 223.650 ;
        RECT 106.060 223.615 125.010 223.915 ;
        RECT 103.350 223.015 120.980 223.315 ;
        RECT 100.590 222.415 116.950 222.715 ;
        RECT 97.830 221.815 112.920 222.115 ;
        RECT 95.070 221.215 108.890 221.515 ;
        RECT 1.000 218.590 12.150 220.190 ;
        RECT 106.340 217.515 107.940 220.715 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.920 188.640 10.720 211.890 ;
        RECT 15.720 198.970 38.920 209.370 ;
        RECT 9.520 187.840 11.120 188.640 ;
        RECT 15.720 186.970 38.920 197.370 ;
        RECT 44.120 188.440 44.920 211.890 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.520 182.990 11.120 183.790 ;
        RECT 3.600 176.050 7.510 179.250 ;
        RECT 9.920 163.040 10.720 182.990 ;
        RECT 15.720 174.970 38.920 185.370 ;
        RECT 45.870 181.190 46.670 210.555 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 47.470 182.790 48.270 204.590 ;
        RECT 108.590 202.625 108.890 221.215 ;
        RECT 109.240 207.925 109.640 219.305 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 111.820 207.925 112.220 219.305 ;
        RECT 109.240 207.525 110.490 207.925 ;
        RECT 108.540 201.825 108.940 202.625 ;
        RECT 63.550 200.610 98.400 200.615 ;
        RECT 63.550 199.815 106.330 200.610 ;
        RECT 98.400 199.810 106.330 199.815 ;
        RECT 68.970 196.830 100.300 197.630 ;
        RECT 74.545 193.735 98.000 194.535 ;
        RECT 66.295 190.655 95.650 191.455 ;
        RECT 52.860 188.465 53.660 190.065 ;
        RECT 55.320 184.940 56.920 186.540 ;
        RECT 47.470 181.990 54.670 182.790 ;
        RECT 45.870 180.390 53.020 181.190 ;
        RECT 9.520 162.240 11.120 163.040 ;
        RECT 15.720 162.970 38.920 173.370 ;
        RECT 52.220 170.440 53.020 180.390 ;
        RECT 53.870 175.290 54.670 181.990 ;
        RECT 53.870 164.840 54.670 174.240 ;
        RECT 55.720 166.640 56.520 184.940 ;
        RECT 57.020 177.390 57.820 178.990 ;
        RECT 61.980 174.370 90.220 175.170 ;
        RECT 57.020 168.290 57.820 169.890 ;
        RECT 55.320 165.840 56.920 166.640 ;
        RECT 53.470 164.040 55.070 164.840 ;
        RECT 9.920 153.790 10.720 162.240 ;
        RECT 9.520 152.990 11.120 153.790 ;
        RECT 9.920 152.915 10.720 152.990 ;
        RECT 15.720 150.970 38.920 161.370 ;
        RECT 51.570 160.190 53.170 160.990 ;
        RECT 51.970 155.790 52.770 160.190 ;
        RECT 51.570 154.990 53.170 155.790 ;
        RECT 41.830 149.410 46.630 150.210 ;
        RECT 51.970 148.290 52.770 154.990 ;
        RECT 53.870 151.990 54.670 164.040 ;
        RECT 53.470 151.190 55.070 151.990 ;
        RECT 55.720 150.240 56.520 165.840 ;
        RECT 54.920 149.440 56.520 150.240 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 61.980 143.690 62.780 174.370 ;
        RECT 3.600 132.225 7.510 135.425 ;
        RECT 9.095 134.635 18.955 143.035 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 28.140 142.890 62.780 143.690 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 20.650 131.410 21.050 138.770 ;
        RECT 61.980 135.095 62.780 142.890 ;
        RECT 70.165 172.130 84.650 172.930 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 12.915 45.565 14.515 119.215 ;
        RECT 16.165 56.765 17.765 121.615 ;
        RECT 21.615 95.165 22.415 132.545 ;
        RECT 27.065 95.165 27.865 130.795 ;
        RECT 70.165 128.125 70.965 172.130 ;
        RECT 74.940 154.795 86.100 155.595 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 145.235 75.740 154.795 ;
        RECT 94.850 150.520 95.650 190.655 ;
        RECT 80.010 149.520 95.650 150.520 ;
        RECT 74.940 144.435 86.100 145.235 ;
        RECT 63.315 103.770 64.915 123.715 ;
        RECT 65.865 110.280 67.465 127.485 ;
        RECT 75.510 123.715 77.110 135.155 ;
        RECT 80.125 133.320 80.925 144.435 ;
        RECT 94.850 131.745 95.650 149.520 ;
        RECT 97.200 137.420 98.000 193.735 ;
        RECT 99.500 129.995 100.300 196.830 ;
        RECT 102.950 168.255 103.750 186.540 ;
        RECT 105.530 170.890 106.330 199.810 ;
        RECT 109.240 198.885 109.640 205.545 ;
        RECT 110.090 197.895 110.490 207.525 ;
        RECT 109.240 197.495 110.490 197.895 ;
        RECT 110.970 207.525 112.220 207.925 ;
        RECT 110.970 197.895 111.370 207.525 ;
        RECT 111.820 198.885 112.220 206.755 ;
        RECT 112.620 202.625 112.920 221.815 ;
        RECT 113.270 207.925 113.670 219.305 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 115.850 207.925 116.250 219.305 ;
        RECT 113.270 207.525 114.520 207.925 ;
        RECT 112.570 201.825 112.970 202.625 ;
        RECT 113.270 198.885 113.670 205.545 ;
        RECT 114.120 197.895 114.520 207.525 ;
        RECT 110.970 197.495 112.220 197.895 ;
        RECT 109.240 183.970 109.640 197.495 ;
        RECT 111.820 191.285 112.220 197.495 ;
        RECT 113.270 197.495 114.520 197.895 ;
        RECT 115.000 207.525 116.250 207.925 ;
        RECT 115.000 197.895 115.400 207.525 ;
        RECT 115.850 198.885 116.250 206.755 ;
        RECT 116.650 202.625 116.950 222.415 ;
        RECT 117.300 207.925 117.700 219.305 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 119.880 207.925 120.280 219.305 ;
        RECT 117.300 207.525 118.550 207.925 ;
        RECT 116.600 201.825 117.000 202.625 ;
        RECT 117.300 198.885 117.700 205.545 ;
        RECT 118.150 197.895 118.550 207.525 ;
        RECT 115.000 197.495 116.250 197.895 ;
        RECT 110.530 187.540 110.930 189.140 ;
        RECT 113.270 183.990 113.670 197.495 ;
        RECT 115.850 191.285 116.250 197.495 ;
        RECT 117.300 197.495 118.550 197.895 ;
        RECT 119.030 207.525 120.280 207.925 ;
        RECT 119.030 197.895 119.430 207.525 ;
        RECT 119.880 198.885 120.280 206.755 ;
        RECT 120.680 202.625 120.980 223.015 ;
        RECT 121.330 207.925 121.730 219.305 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 123.910 207.925 124.310 219.305 ;
        RECT 121.330 207.525 122.580 207.925 ;
        RECT 120.630 201.825 121.030 202.625 ;
        RECT 121.330 198.885 121.730 205.545 ;
        RECT 122.180 197.895 122.580 207.525 ;
        RECT 119.030 197.495 120.280 197.895 ;
        RECT 114.560 187.540 114.960 189.140 ;
        RECT 111.685 183.590 113.670 183.990 ;
        RECT 105.530 168.255 106.730 170.890 ;
        RECT 107.380 168.490 107.780 170.890 ;
        RECT 103.350 152.765 103.750 160.495 ;
        RECT 103.350 143.435 103.750 145.835 ;
        RECT 104.640 140.165 105.040 167.190 ;
        RECT 105.385 157.365 105.785 158.165 ;
        RECT 106.330 145.835 106.730 168.255 ;
        RECT 107.380 152.765 107.780 160.495 ;
        RECT 108.670 147.135 109.070 178.990 ;
        RECT 109.960 168.490 110.760 170.890 ;
        RECT 109.415 156.165 109.815 156.965 ;
        RECT 110.360 145.835 110.760 168.490 ;
        RECT 111.685 157.765 112.085 183.590 ;
        RECT 117.300 182.580 117.700 197.495 ;
        RECT 119.880 191.285 120.280 197.495 ;
        RECT 121.330 197.495 122.580 197.895 ;
        RECT 123.060 207.525 124.310 207.925 ;
        RECT 123.060 197.895 123.460 207.525 ;
        RECT 123.910 198.885 124.310 206.755 ;
        RECT 124.710 202.625 125.010 223.615 ;
        RECT 125.360 207.925 125.760 219.305 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 127.940 207.925 128.340 219.305 ;
        RECT 125.360 207.525 126.610 207.925 ;
        RECT 124.660 201.825 125.060 202.625 ;
        RECT 125.360 198.885 125.760 205.545 ;
        RECT 126.210 197.895 126.610 207.525 ;
        RECT 123.060 197.495 124.310 197.895 ;
        RECT 118.590 187.540 118.990 189.140 ;
        RECT 113.085 182.180 117.700 182.580 ;
        RECT 113.085 156.165 113.485 182.180 ;
        RECT 121.330 181.545 121.730 197.495 ;
        RECT 123.910 191.285 124.310 197.495 ;
        RECT 125.360 197.495 126.610 197.895 ;
        RECT 127.090 207.525 128.340 207.925 ;
        RECT 127.090 197.895 127.490 207.525 ;
        RECT 127.940 198.885 128.340 206.755 ;
        RECT 128.740 202.625 129.040 224.215 ;
        RECT 132.720 220.715 133.120 221.515 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 129.390 207.925 129.790 219.305 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 131.970 207.925 132.370 219.305 ;
        RECT 129.390 207.525 130.640 207.925 ;
        RECT 128.690 201.825 129.090 202.625 ;
        RECT 129.390 198.885 129.790 205.545 ;
        RECT 130.240 197.895 130.640 207.525 ;
        RECT 127.090 197.495 128.340 197.895 ;
        RECT 122.620 187.540 123.020 189.140 ;
        RECT 116.415 181.145 121.730 181.545 ;
        RECT 116.415 176.215 116.815 181.145 ;
        RECT 125.360 180.565 125.760 197.495 ;
        RECT 127.940 191.285 128.340 197.495 ;
        RECT 129.390 197.495 130.640 197.895 ;
        RECT 131.120 207.525 132.370 207.925 ;
        RECT 131.120 197.895 131.520 207.525 ;
        RECT 131.970 198.885 132.370 206.755 ;
        RECT 132.770 202.625 133.070 220.715 ;
        RECT 133.420 207.925 133.820 219.305 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 136.000 207.925 136.400 219.305 ;
        RECT 133.420 207.525 134.670 207.925 ;
        RECT 132.720 201.825 133.120 202.625 ;
        RECT 133.420 198.885 133.820 205.545 ;
        RECT 134.270 197.895 134.670 207.525 ;
        RECT 131.120 197.495 132.370 197.895 ;
        RECT 126.650 187.540 127.050 189.140 ;
        RECT 121.035 180.165 125.760 180.565 ;
        RECT 121.035 176.215 121.435 180.165 ;
        RECT 129.390 179.490 129.790 197.495 ;
        RECT 131.970 191.285 132.370 197.495 ;
        RECT 133.420 197.495 134.670 197.895 ;
        RECT 135.150 207.525 136.400 207.925 ;
        RECT 135.150 197.895 135.550 207.525 ;
        RECT 136.000 198.885 136.400 206.755 ;
        RECT 136.800 202.625 137.100 220.715 ;
        RECT 137.450 207.925 137.850 219.305 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 140.030 207.925 140.430 219.305 ;
        RECT 137.450 207.525 138.700 207.925 ;
        RECT 136.750 201.825 137.150 202.625 ;
        RECT 137.450 198.885 137.850 205.545 ;
        RECT 138.300 197.895 138.700 207.525 ;
        RECT 135.150 197.495 136.400 197.895 ;
        RECT 130.680 187.540 131.080 189.140 ;
        RECT 125.660 179.090 129.790 179.490 ;
        RECT 125.660 176.215 126.060 179.090 ;
        RECT 133.420 178.920 133.820 197.495 ;
        RECT 136.000 191.285 136.400 197.495 ;
        RECT 137.450 197.495 138.700 197.895 ;
        RECT 139.180 207.525 140.430 207.925 ;
        RECT 139.180 197.895 139.580 207.525 ;
        RECT 140.030 198.885 140.430 206.755 ;
        RECT 140.830 202.625 141.130 220.715 ;
        RECT 141.480 207.925 141.880 219.305 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 144.060 207.925 144.460 219.305 ;
        RECT 141.480 207.525 142.730 207.925 ;
        RECT 140.780 201.825 141.180 202.625 ;
        RECT 141.480 198.885 141.880 205.545 ;
        RECT 142.330 197.895 142.730 207.525 ;
        RECT 139.180 197.495 140.430 197.895 ;
        RECT 134.710 187.540 135.110 189.140 ;
        RECT 137.450 178.920 137.850 197.495 ;
        RECT 140.030 191.285 140.430 197.495 ;
        RECT 141.480 197.495 142.730 197.895 ;
        RECT 143.210 207.525 144.460 207.925 ;
        RECT 143.210 197.895 143.610 207.525 ;
        RECT 144.060 198.885 144.460 206.755 ;
        RECT 144.860 202.625 145.160 220.715 ;
        RECT 145.510 207.925 145.910 219.305 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 148.090 207.925 148.490 219.305 ;
        RECT 145.510 207.525 146.760 207.925 ;
        RECT 144.810 201.825 145.210 202.625 ;
        RECT 145.510 198.885 145.910 205.545 ;
        RECT 146.360 197.895 146.760 207.525 ;
        RECT 143.210 197.495 144.460 197.895 ;
        RECT 138.740 187.540 139.140 189.140 ;
        RECT 141.480 178.920 141.880 197.495 ;
        RECT 144.060 191.285 144.460 197.495 ;
        RECT 145.510 197.495 146.760 197.895 ;
        RECT 147.240 207.525 148.490 207.925 ;
        RECT 147.240 197.895 147.640 207.525 ;
        RECT 148.090 198.885 148.490 206.755 ;
        RECT 148.890 202.625 149.190 220.715 ;
        RECT 149.540 207.925 149.940 219.305 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 152.120 207.925 152.520 219.305 ;
        RECT 149.540 207.525 150.790 207.925 ;
        RECT 148.840 201.825 149.240 202.625 ;
        RECT 149.540 198.885 149.940 205.545 ;
        RECT 150.390 197.895 150.790 207.525 ;
        RECT 147.240 197.495 148.490 197.895 ;
        RECT 142.770 187.540 143.170 189.140 ;
        RECT 145.510 178.920 145.910 197.495 ;
        RECT 148.090 191.285 148.490 197.495 ;
        RECT 149.540 197.495 150.790 197.895 ;
        RECT 151.270 207.525 152.520 207.925 ;
        RECT 151.270 197.895 151.670 207.525 ;
        RECT 152.120 198.885 152.520 206.755 ;
        RECT 151.270 197.495 152.520 197.895 ;
        RECT 146.800 187.540 147.200 189.140 ;
        RECT 149.540 178.920 149.940 197.495 ;
        RECT 152.120 191.285 152.520 197.495 ;
        RECT 150.830 187.540 151.230 189.140 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 130.275 178.520 133.820 178.920 ;
        RECT 134.895 178.520 137.850 178.920 ;
        RECT 139.510 178.520 141.880 178.920 ;
        RECT 144.135 178.520 145.910 178.920 ;
        RECT 148.755 178.520 149.940 178.920 ;
        RECT 130.275 176.215 130.675 178.520 ;
        RECT 134.895 176.215 135.295 178.520 ;
        RECT 139.510 176.215 139.910 178.520 ;
        RECT 144.135 176.215 144.535 178.520 ;
        RECT 148.755 176.215 149.155 178.520 ;
        RECT 116.215 175.815 117.015 176.215 ;
        RECT 120.835 175.815 121.635 176.215 ;
        RECT 125.455 175.815 126.255 176.215 ;
        RECT 130.075 175.815 130.875 176.215 ;
        RECT 134.695 175.815 135.495 176.215 ;
        RECT 139.315 175.815 140.115 176.215 ;
        RECT 143.935 175.815 144.735 176.215 ;
        RECT 148.555 175.815 149.355 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 115.815 173.070 117.415 173.870 ;
        RECT 120.435 173.070 122.035 173.870 ;
        RECT 125.055 173.070 126.655 173.870 ;
        RECT 129.675 173.070 131.275 173.870 ;
        RECT 134.295 173.070 135.895 173.870 ;
        RECT 138.915 173.070 140.515 173.870 ;
        RECT 143.535 173.070 145.135 173.870 ;
        RECT 148.155 173.070 149.755 173.870 ;
        RECT 105.930 143.435 106.730 145.835 ;
        RECT 104.640 139.365 105.440 140.165 ;
        RECT 107.380 136.325 107.780 145.835 ;
        RECT 109.960 143.435 110.760 145.835 ;
        RECT 116.310 144.730 116.910 173.070 ;
        RECT 120.930 147.530 121.530 173.070 ;
        RECT 125.550 148.690 126.150 173.070 ;
        RECT 130.175 149.890 130.775 173.070 ;
        RECT 134.795 160.260 135.395 173.070 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 133.275 152.100 134.875 152.200 ;
        RECT 136.875 152.100 137.475 161.650 ;
        RECT 133.275 151.500 137.475 152.100 ;
        RECT 133.275 151.400 134.875 151.500 ;
        RECT 133.275 150.930 134.875 151.030 ;
        RECT 139.410 150.930 140.010 173.070 ;
        RECT 144.035 162.450 144.635 173.070 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 148.655 161.210 149.255 173.070 ;
        RECT 133.275 150.330 140.010 150.930 ;
        RECT 141.715 160.610 149.255 161.210 ;
        RECT 133.275 150.230 134.875 150.330 ;
        RECT 130.175 149.290 136.695 149.890 ;
        RECT 125.550 148.090 133.635 148.690 ;
        RECT 130.615 147.530 132.215 147.630 ;
        RECT 120.930 146.930 132.215 147.530 ;
        RECT 130.615 146.830 132.215 146.930 ;
        RECT 122.645 144.730 124.245 144.830 ;
        RECT 116.310 144.130 124.245 144.730 ;
        RECT 122.645 144.030 124.245 144.130 ;
        RECT 133.035 144.520 133.635 148.090 ;
        RECT 136.095 148.010 136.695 149.290 ;
        RECT 138.525 148.010 140.125 148.110 ;
        RECT 136.095 147.410 140.125 148.010 ;
        RECT 138.525 147.310 140.125 147.410 ;
        RECT 138.525 144.520 140.125 144.620 ;
        RECT 133.035 143.920 140.125 144.520 ;
        RECT 141.715 144.040 142.315 160.610 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 138.525 143.820 140.125 143.920 ;
        RECT 109.960 138.220 110.360 143.435 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 142.690 142.815 142.790 ;
        RECT 145.625 142.690 146.225 159.460 ;
        RECT 141.215 142.090 146.225 142.690 ;
        RECT 141.215 141.990 142.815 142.090 ;
        RECT 109.560 137.420 110.760 138.220 ;
        RECT 107.380 135.525 108.180 136.325 ;
        RECT 72.765 103.865 74.365 122.215 ;
        RECT 75.510 114.215 77.115 123.715 ;
        RECT 75.515 100.215 77.115 114.215 ;
        RECT 21.215 51.675 22.815 95.165 ;
        RECT 26.665 61.465 28.265 95.165 ;
        RECT 97.165 93.265 98.765 119.215 ;
        RECT 100.515 117.715 101.315 128.925 ;
        RECT 100.115 96.415 101.715 117.715 ;
        RECT 103.315 111.365 104.915 123.165 ;
        RECT 116.915 121.965 118.515 122.765 ;
        RECT 105.965 103.965 107.565 120.665 ;
        RECT 109.865 108.365 111.465 119.215 ;
        RECT 117.115 108.365 118.715 118.265 ;
        RECT 121.565 113.015 123.165 127.485 ;
        RECT 116.965 104.015 118.565 104.815 ;
        RECT 42.740 71.190 53.140 83.050 ;
        RECT 55.740 71.190 66.140 83.050 ;
        RECT 68.740 71.190 79.140 83.050 ;
        RECT 81.740 71.190 92.140 83.050 ;
        RECT 94.740 71.190 105.140 83.050 ;
        RECT 42.740 57.830 53.140 69.690 ;
        RECT 55.740 57.830 66.140 69.690 ;
        RECT 68.740 57.830 79.140 69.690 ;
        RECT 81.740 57.830 92.140 69.690 ;
        RECT 94.740 57.830 105.140 69.690 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 3.600 36.430 8.665 39.630 ;
        RECT 3.600 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 34.940 ;
        RECT 65.765 15.915 67.365 44.215 ;
        RECT 68.865 11.965 70.465 41.615 ;
        RECT 72.095 9.665 73.695 38.865 ;
        RECT 80.745 9.665 82.345 37.635 ;
        RECT 84.015 22.315 85.615 41.615 ;
        RECT 87.165 26.815 88.765 44.215 ;
        RECT 90.715 19.315 92.315 47.165 ;
        RECT 116.115 42.615 117.715 90.815 ;
        RECT 119.215 40.015 120.815 84.315 ;
        RECT 123.215 23.815 124.815 94.865 ;
        RECT 126.165 25.365 127.765 98.015 ;
        RECT 128.965 5.690 130.565 8.890 ;
        RECT 2.705 1.285 98.380 2.085 ;
        RECT 131.665 1.800 132.465 136.325 ;
        RECT 133.265 111.795 134.065 130.795 ;
        RECT 134.865 110.315 135.665 132.545 ;
        RECT 136.465 114.770 137.265 134.120 ;
        RECT 137.945 133.410 138.745 133.810 ;
        RECT 137.945 131.410 138.345 133.410 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.970 125.690 142.100 127.290 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 133.525 109.515 138.400 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 136.495 29.375 138.195 94.305 ;
        RECT 139.355 30.545 141.055 114.150 ;
        RECT 141.900 110.315 142.700 117.170 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 141.495 20.015 143.195 110.315 ;
        RECT 143.640 32.885 145.340 114.150 ;
        RECT 146.950 110.315 147.750 138.220 ;
        RECT 149.945 116.370 150.745 170.845 ;
        RECT 146.490 104.255 148.190 110.315 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 151.560 1.800 152.360 140.165 ;
        RECT 153.945 129.145 154.345 184.370 ;
      LAYER met4 ;
        RECT 15.030 224.460 15.330 224.760 ;
        RECT 17.790 224.460 18.090 224.760 ;
        RECT 20.550 224.460 20.850 224.760 ;
        RECT 23.310 224.460 23.610 224.760 ;
        RECT 26.070 224.460 26.370 224.760 ;
        RECT 28.830 224.460 29.130 224.760 ;
        RECT 31.590 224.460 31.890 224.760 ;
        RECT 34.350 224.460 34.650 224.760 ;
        RECT 37.110 224.460 37.410 224.760 ;
        RECT 39.870 224.460 40.170 224.760 ;
        RECT 42.630 224.460 42.930 224.760 ;
        RECT 45.390 224.460 45.690 224.760 ;
        RECT 48.150 224.460 48.450 224.760 ;
        RECT 50.910 224.460 51.210 224.760 ;
        RECT 53.670 224.460 53.970 224.760 ;
        RECT 56.430 224.460 56.730 224.760 ;
        RECT 59.190 224.460 59.490 224.760 ;
        RECT 61.950 224.460 62.250 224.760 ;
        RECT 64.710 224.460 65.010 224.760 ;
        RECT 67.470 224.460 67.770 224.760 ;
        RECT 70.230 224.460 70.530 224.760 ;
        RECT 72.990 224.460 73.290 224.760 ;
        RECT 75.750 224.460 76.050 224.760 ;
        RECT 78.510 224.460 78.810 224.760 ;
        RECT 3.600 224.060 78.810 224.460 ;
        RECT 95.070 224.450 95.370 224.760 ;
        RECT 97.830 224.450 98.130 224.760 ;
        RECT 100.590 224.450 100.890 224.760 ;
        RECT 103.350 224.450 103.650 224.760 ;
        RECT 106.110 224.450 106.410 224.760 ;
        RECT 108.870 224.615 109.170 224.760 ;
        RECT 3.600 220.760 5.200 224.060 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.650 106.460 224.450 ;
        RECT 108.865 224.215 109.665 224.615 ;
        RECT 6.200 221.180 109.540 222.780 ;
        RECT 111.630 221.515 111.930 224.760 ;
        RECT 114.390 222.115 114.690 224.760 ;
        RECT 117.150 222.715 117.450 224.760 ;
        RECT 119.910 223.315 120.210 224.760 ;
        RECT 122.670 223.915 122.970 224.760 ;
        RECT 122.670 223.615 149.190 223.915 ;
        RECT 119.910 223.015 145.160 223.315 ;
        RECT 117.150 222.415 141.130 222.715 ;
        RECT 114.390 221.815 137.100 222.115 ;
        RECT 136.800 221.515 137.100 221.815 ;
        RECT 140.830 221.515 141.130 222.415 ;
        RECT 144.860 221.515 145.160 223.015 ;
        RECT 148.890 221.515 149.190 223.615 ;
        RECT 111.630 221.215 133.120 221.515 ;
        RECT 6.200 220.760 7.800 221.180 ;
        RECT 10.550 218.590 105.040 220.190 ;
        RECT 7.800 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 103.440 211.240 105.040 218.590 ;
        RECT 106.340 219.305 109.540 221.180 ;
        RECT 132.720 220.715 133.120 221.215 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 106.340 217.705 151.230 219.305 ;
        RECT 106.340 217.515 109.540 217.705 ;
        RECT 106.415 211.240 108.015 213.740 ;
        RECT 27.080 209.940 53.660 210.740 ;
        RECT 27.080 209.640 27.570 209.940 ;
        RECT 16.115 199.365 25.725 208.975 ;
        RECT 16.115 196.975 16.715 199.365 ;
        RECT 16.115 187.365 25.725 196.975 ;
        RECT 16.115 184.975 16.715 187.365 ;
        RECT 16.115 175.365 25.725 184.975 ;
        RECT 16.115 172.975 16.715 175.365 ;
        RECT 16.115 163.365 25.725 172.975 ;
        RECT 16.115 160.975 16.715 163.365 ;
        RECT 16.115 151.365 25.725 160.975 ;
        RECT 16.115 150.210 16.715 151.365 ;
        RECT 27.080 150.970 27.565 209.640 ;
        RECT 28.915 199.365 38.525 208.975 ;
        RECT 37.925 196.975 38.525 199.365 ;
        RECT 28.915 187.365 38.525 196.975 ;
        RECT 52.860 188.465 53.660 209.940 ;
        RECT 103.440 209.640 151.230 211.240 ;
        RECT 110.530 187.540 156.765 189.140 ;
        RECT 37.925 184.975 38.525 187.365 ;
        RECT 28.915 175.365 38.525 184.975 ;
        RECT 37.925 172.975 38.525 175.365 ;
        RECT 28.915 163.365 38.525 172.975 ;
        RECT 51.950 184.940 103.750 186.540 ;
        RECT 51.950 169.890 53.550 184.940 ;
        RECT 57.020 177.390 109.070 178.990 ;
        RECT 153.565 178.210 156.765 187.540 ;
        RECT 151.155 175.010 156.765 178.210 ;
        RECT 51.950 168.290 58.420 169.890 ;
        RECT 37.925 160.975 38.525 163.365 ;
        RECT 28.915 151.365 38.525 160.975 ;
        RECT 111.685 158.165 112.085 158.565 ;
        RECT 105.385 157.765 112.085 158.165 ;
        RECT 105.385 157.365 105.785 157.765 ;
        RECT 109.415 156.565 109.815 156.965 ;
        RECT 113.085 156.565 113.485 156.965 ;
        RECT 109.415 156.165 113.485 156.565 ;
        RECT 37.925 150.210 38.525 151.365 ;
        RECT 16.115 149.410 46.630 150.210 ;
        RECT 51.575 145.090 73.495 148.290 ;
        RECT 9.490 135.030 17.100 142.640 ;
        RECT 18.455 142.175 20.750 142.975 ;
        RECT 13.385 130.025 14.185 135.030 ;
        RECT 18.455 134.695 18.935 142.175 ;
        RECT 20.350 141.375 20.750 142.175 ;
        RECT 61.980 135.495 62.780 135.895 ;
        RECT 61.980 135.095 140.370 135.495 ;
        RECT 22.615 133.320 80.925 134.120 ;
        RECT 20.650 131.810 21.050 132.210 ;
        RECT 137.945 131.810 138.345 132.210 ;
        RECT 20.650 131.410 138.345 131.810 ;
        RECT 139.120 130.025 139.520 132.990 ;
        RECT 13.385 129.625 139.520 130.025 ;
        RECT 16.805 128.710 139.520 129.110 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 128.710 ;
        RECT 139.970 125.690 140.370 135.095 ;
        RECT 140.940 131.390 142.100 132.990 ;
        RECT 140.940 125.060 141.340 131.390 ;
        RECT 131.145 124.660 141.340 125.060 ;
        RECT 103.315 121.565 118.965 123.165 ;
        RECT 109.865 107.965 118.715 109.565 ;
        RECT 63.315 103.465 74.365 105.065 ;
        RECT 105.965 103.615 118.565 105.215 ;
        RECT 131.145 98.015 131.545 124.660 ;
        RECT 153.565 124.090 156.765 175.010 ;
        RECT 142.760 122.490 156.765 124.090 ;
        RECT 153.565 114.150 156.765 122.490 ;
        RECT 139.355 113.350 156.765 114.150 ;
        RECT 100.115 96.415 132.145 98.015 ;
        RECT 97.165 93.265 124.815 94.865 ;
        RECT 43.135 78.605 52.745 82.655 ;
        RECT 56.135 78.605 65.745 82.655 ;
        RECT 69.135 78.605 78.745 82.655 ;
        RECT 82.135 78.605 91.745 82.655 ;
        RECT 95.135 78.605 104.745 82.655 ;
        RECT 130.545 78.605 132.145 96.415 ;
        RECT 38.470 77.005 132.145 78.605 ;
        RECT 38.470 63.590 39.745 77.005 ;
        RECT 43.135 73.045 52.745 77.005 ;
        RECT 56.135 73.045 65.745 77.005 ;
        RECT 69.135 73.045 78.745 77.005 ;
        RECT 82.135 73.045 91.745 77.005 ;
        RECT 95.135 73.045 104.745 77.005 ;
        RECT 42.800 71.180 108.800 71.690 ;
        RECT 133.525 71.180 135.125 110.315 ;
        RECT 42.800 69.580 135.125 71.180 ;
        RECT 42.800 69.190 108.800 69.580 ;
        RECT 43.135 63.590 52.745 67.835 ;
        RECT 56.135 63.590 65.745 67.835 ;
        RECT 69.135 63.590 78.745 67.835 ;
        RECT 82.135 63.590 91.745 67.835 ;
        RECT 95.135 63.590 104.745 67.835 ;
        RECT 38.470 61.990 104.745 63.590 ;
        RECT 43.135 58.225 52.745 61.990 ;
        RECT 56.135 58.225 65.745 61.990 ;
        RECT 69.135 58.225 78.745 61.990 ;
        RECT 82.135 58.225 91.745 61.990 ;
        RECT 95.135 58.225 104.745 61.990 ;
        RECT 12.915 45.565 92.315 47.165 ;
        RECT 65.765 42.615 117.715 44.215 ;
        RECT 68.865 40.015 120.815 41.615 ;
        RECT 72.095 9.265 82.535 10.865 ;
        RECT 153.565 8.890 156.765 113.350 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.160 5.690 156.765 8.890 ;
        RECT 97.530 1.000 98.430 2.125 ;
        RECT 116.850 1.750 132.465 2.650 ;
        RECT 136.170 1.750 152.360 2.650 ;
        RECT 116.850 1.000 117.750 1.750 ;
        RECT 136.170 1.000 137.070 1.750 ;
  END
END tt_um_cw_vref
END LIBRARY

