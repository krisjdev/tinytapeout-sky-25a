module tt_um_delaychain (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire \thechain[0].chain1.dout ;
 wire \thechain[0].chain1.inv_chain[0] ;
 wire \thechain[0].chain1.inv_chain[1] ;
 wire \thechain[0].chain1.inv_chain[2] ;
 wire \thechain[0].chain2.dout ;
 wire \thechain[0].chain2.inv_chain[0] ;
 wire \thechain[0].chain2.inv_chain[1] ;
 wire \thechain[0].chain2.inv_chain[2] ;
 wire \thechain[0].chain2.inv_chain[3] ;
 wire \thechain[0].chain2.inv_chain[4] ;
 wire \thechain[0].chain3.dout ;
 wire \thechain[0].chain3.inv_chain[0] ;
 wire \thechain[0].chain3.inv_chain[1] ;
 wire \thechain[0].chain3.inv_chain[2] ;
 wire \thechain[0].chain3.inv_chain[3] ;
 wire \thechain[0].chain3.inv_chain[4] ;
 wire \thechain[0].chain3.inv_chain[5] ;
 wire \thechain[0].chain3.inv_chain[6] ;
 wire \thechain[0].chain3.inv_chain[7] ;
 wire \thechain[0].chain3.inv_chain[8] ;
 wire \thechain[0].chain4.dout ;
 wire \thechain[0].chain4.inv_chain[0] ;
 wire \thechain[0].chain4.inv_chain[10] ;
 wire \thechain[0].chain4.inv_chain[11] ;
 wire \thechain[0].chain4.inv_chain[12] ;
 wire \thechain[0].chain4.inv_chain[13] ;
 wire \thechain[0].chain4.inv_chain[14] ;
 wire \thechain[0].chain4.inv_chain[15] ;
 wire \thechain[0].chain4.inv_chain[16] ;
 wire \thechain[0].chain4.inv_chain[1] ;
 wire \thechain[0].chain4.inv_chain[2] ;
 wire \thechain[0].chain4.inv_chain[3] ;
 wire \thechain[0].chain4.inv_chain[4] ;
 wire \thechain[0].chain4.inv_chain[5] ;
 wire \thechain[0].chain4.inv_chain[6] ;
 wire \thechain[0].chain4.inv_chain[7] ;
 wire \thechain[0].chain4.inv_chain[8] ;
 wire \thechain[0].chain4.inv_chain[9] ;
 wire \thechain[0].chain5.dout ;
 wire \thechain[0].chain5.inv_chain[0] ;
 wire \thechain[0].chain5.inv_chain[10] ;
 wire \thechain[0].chain5.inv_chain[11] ;
 wire \thechain[0].chain5.inv_chain[12] ;
 wire \thechain[0].chain5.inv_chain[13] ;
 wire \thechain[0].chain5.inv_chain[14] ;
 wire \thechain[0].chain5.inv_chain[15] ;
 wire \thechain[0].chain5.inv_chain[16] ;
 wire \thechain[0].chain5.inv_chain[17] ;
 wire \thechain[0].chain5.inv_chain[18] ;
 wire \thechain[0].chain5.inv_chain[19] ;
 wire \thechain[0].chain5.inv_chain[1] ;
 wire \thechain[0].chain5.inv_chain[20] ;
 wire \thechain[0].chain5.inv_chain[21] ;
 wire \thechain[0].chain5.inv_chain[22] ;
 wire \thechain[0].chain5.inv_chain[23] ;
 wire \thechain[0].chain5.inv_chain[24] ;
 wire \thechain[0].chain5.inv_chain[25] ;
 wire \thechain[0].chain5.inv_chain[26] ;
 wire \thechain[0].chain5.inv_chain[27] ;
 wire \thechain[0].chain5.inv_chain[28] ;
 wire \thechain[0].chain5.inv_chain[29] ;
 wire \thechain[0].chain5.inv_chain[2] ;
 wire \thechain[0].chain5.inv_chain[30] ;
 wire \thechain[0].chain5.inv_chain[31] ;
 wire \thechain[0].chain5.inv_chain[32] ;
 wire \thechain[0].chain5.inv_chain[3] ;
 wire \thechain[0].chain5.inv_chain[4] ;
 wire \thechain[0].chain5.inv_chain[5] ;
 wire \thechain[0].chain5.inv_chain[6] ;
 wire \thechain[0].chain5.inv_chain[7] ;
 wire \thechain[0].chain5.inv_chain[8] ;
 wire \thechain[0].chain5.inv_chain[9] ;
 wire \thechain[0].chain6.dout ;
 wire \thechain[0].chain6.inv_chain[0] ;
 wire \thechain[0].chain6.inv_chain[10] ;
 wire \thechain[0].chain6.inv_chain[11] ;
 wire \thechain[0].chain6.inv_chain[12] ;
 wire \thechain[0].chain6.inv_chain[13] ;
 wire \thechain[0].chain6.inv_chain[14] ;
 wire \thechain[0].chain6.inv_chain[15] ;
 wire \thechain[0].chain6.inv_chain[16] ;
 wire \thechain[0].chain6.inv_chain[17] ;
 wire \thechain[0].chain6.inv_chain[18] ;
 wire \thechain[0].chain6.inv_chain[19] ;
 wire \thechain[0].chain6.inv_chain[1] ;
 wire \thechain[0].chain6.inv_chain[20] ;
 wire \thechain[0].chain6.inv_chain[21] ;
 wire \thechain[0].chain6.inv_chain[22] ;
 wire \thechain[0].chain6.inv_chain[23] ;
 wire \thechain[0].chain6.inv_chain[24] ;
 wire \thechain[0].chain6.inv_chain[25] ;
 wire \thechain[0].chain6.inv_chain[26] ;
 wire \thechain[0].chain6.inv_chain[27] ;
 wire \thechain[0].chain6.inv_chain[28] ;
 wire \thechain[0].chain6.inv_chain[29] ;
 wire \thechain[0].chain6.inv_chain[2] ;
 wire \thechain[0].chain6.inv_chain[30] ;
 wire \thechain[0].chain6.inv_chain[31] ;
 wire \thechain[0].chain6.inv_chain[32] ;
 wire \thechain[0].chain6.inv_chain[33] ;
 wire \thechain[0].chain6.inv_chain[34] ;
 wire \thechain[0].chain6.inv_chain[35] ;
 wire \thechain[0].chain6.inv_chain[36] ;
 wire \thechain[0].chain6.inv_chain[37] ;
 wire \thechain[0].chain6.inv_chain[38] ;
 wire \thechain[0].chain6.inv_chain[39] ;
 wire \thechain[0].chain6.inv_chain[3] ;
 wire \thechain[0].chain6.inv_chain[40] ;
 wire \thechain[0].chain6.inv_chain[41] ;
 wire \thechain[0].chain6.inv_chain[42] ;
 wire \thechain[0].chain6.inv_chain[43] ;
 wire \thechain[0].chain6.inv_chain[44] ;
 wire \thechain[0].chain6.inv_chain[45] ;
 wire \thechain[0].chain6.inv_chain[46] ;
 wire \thechain[0].chain6.inv_chain[47] ;
 wire \thechain[0].chain6.inv_chain[48] ;
 wire \thechain[0].chain6.inv_chain[49] ;
 wire \thechain[0].chain6.inv_chain[4] ;
 wire \thechain[0].chain6.inv_chain[50] ;
 wire \thechain[0].chain6.inv_chain[51] ;
 wire \thechain[0].chain6.inv_chain[52] ;
 wire \thechain[0].chain6.inv_chain[53] ;
 wire \thechain[0].chain6.inv_chain[54] ;
 wire \thechain[0].chain6.inv_chain[55] ;
 wire \thechain[0].chain6.inv_chain[56] ;
 wire \thechain[0].chain6.inv_chain[57] ;
 wire \thechain[0].chain6.inv_chain[58] ;
 wire \thechain[0].chain6.inv_chain[59] ;
 wire \thechain[0].chain6.inv_chain[5] ;
 wire \thechain[0].chain6.inv_chain[60] ;
 wire \thechain[0].chain6.inv_chain[61] ;
 wire \thechain[0].chain6.inv_chain[62] ;
 wire \thechain[0].chain6.inv_chain[63] ;
 wire \thechain[0].chain6.inv_chain[64] ;
 wire \thechain[0].chain6.inv_chain[6] ;
 wire \thechain[0].chain6.inv_chain[7] ;
 wire \thechain[0].chain6.inv_chain[8] ;
 wire \thechain[0].chain6.inv_chain[9] ;
 wire \thechain[0].chain7.dout ;
 wire \thechain[0].chain7.inv_chain[0] ;
 wire \thechain[0].chain7.inv_chain[100] ;
 wire \thechain[0].chain7.inv_chain[101] ;
 wire \thechain[0].chain7.inv_chain[102] ;
 wire \thechain[0].chain7.inv_chain[103] ;
 wire \thechain[0].chain7.inv_chain[104] ;
 wire \thechain[0].chain7.inv_chain[105] ;
 wire \thechain[0].chain7.inv_chain[106] ;
 wire \thechain[0].chain7.inv_chain[107] ;
 wire \thechain[0].chain7.inv_chain[108] ;
 wire \thechain[0].chain7.inv_chain[109] ;
 wire \thechain[0].chain7.inv_chain[10] ;
 wire \thechain[0].chain7.inv_chain[110] ;
 wire \thechain[0].chain7.inv_chain[111] ;
 wire \thechain[0].chain7.inv_chain[112] ;
 wire \thechain[0].chain7.inv_chain[113] ;
 wire \thechain[0].chain7.inv_chain[114] ;
 wire \thechain[0].chain7.inv_chain[115] ;
 wire \thechain[0].chain7.inv_chain[116] ;
 wire \thechain[0].chain7.inv_chain[117] ;
 wire \thechain[0].chain7.inv_chain[118] ;
 wire \thechain[0].chain7.inv_chain[119] ;
 wire \thechain[0].chain7.inv_chain[11] ;
 wire \thechain[0].chain7.inv_chain[120] ;
 wire \thechain[0].chain7.inv_chain[121] ;
 wire \thechain[0].chain7.inv_chain[122] ;
 wire \thechain[0].chain7.inv_chain[123] ;
 wire \thechain[0].chain7.inv_chain[124] ;
 wire \thechain[0].chain7.inv_chain[125] ;
 wire \thechain[0].chain7.inv_chain[126] ;
 wire \thechain[0].chain7.inv_chain[127] ;
 wire \thechain[0].chain7.inv_chain[128] ;
 wire \thechain[0].chain7.inv_chain[12] ;
 wire \thechain[0].chain7.inv_chain[13] ;
 wire \thechain[0].chain7.inv_chain[14] ;
 wire \thechain[0].chain7.inv_chain[15] ;
 wire \thechain[0].chain7.inv_chain[16] ;
 wire \thechain[0].chain7.inv_chain[17] ;
 wire \thechain[0].chain7.inv_chain[18] ;
 wire \thechain[0].chain7.inv_chain[19] ;
 wire \thechain[0].chain7.inv_chain[1] ;
 wire \thechain[0].chain7.inv_chain[20] ;
 wire \thechain[0].chain7.inv_chain[21] ;
 wire \thechain[0].chain7.inv_chain[22] ;
 wire \thechain[0].chain7.inv_chain[23] ;
 wire \thechain[0].chain7.inv_chain[24] ;
 wire \thechain[0].chain7.inv_chain[25] ;
 wire \thechain[0].chain7.inv_chain[26] ;
 wire \thechain[0].chain7.inv_chain[27] ;
 wire \thechain[0].chain7.inv_chain[28] ;
 wire \thechain[0].chain7.inv_chain[29] ;
 wire \thechain[0].chain7.inv_chain[2] ;
 wire \thechain[0].chain7.inv_chain[30] ;
 wire \thechain[0].chain7.inv_chain[31] ;
 wire \thechain[0].chain7.inv_chain[32] ;
 wire \thechain[0].chain7.inv_chain[33] ;
 wire \thechain[0].chain7.inv_chain[34] ;
 wire \thechain[0].chain7.inv_chain[35] ;
 wire \thechain[0].chain7.inv_chain[36] ;
 wire \thechain[0].chain7.inv_chain[37] ;
 wire \thechain[0].chain7.inv_chain[38] ;
 wire \thechain[0].chain7.inv_chain[39] ;
 wire \thechain[0].chain7.inv_chain[3] ;
 wire \thechain[0].chain7.inv_chain[40] ;
 wire \thechain[0].chain7.inv_chain[41] ;
 wire \thechain[0].chain7.inv_chain[42] ;
 wire \thechain[0].chain7.inv_chain[43] ;
 wire \thechain[0].chain7.inv_chain[44] ;
 wire \thechain[0].chain7.inv_chain[45] ;
 wire \thechain[0].chain7.inv_chain[46] ;
 wire \thechain[0].chain7.inv_chain[47] ;
 wire \thechain[0].chain7.inv_chain[48] ;
 wire \thechain[0].chain7.inv_chain[49] ;
 wire \thechain[0].chain7.inv_chain[4] ;
 wire \thechain[0].chain7.inv_chain[50] ;
 wire \thechain[0].chain7.inv_chain[51] ;
 wire \thechain[0].chain7.inv_chain[52] ;
 wire \thechain[0].chain7.inv_chain[53] ;
 wire \thechain[0].chain7.inv_chain[54] ;
 wire \thechain[0].chain7.inv_chain[55] ;
 wire \thechain[0].chain7.inv_chain[56] ;
 wire \thechain[0].chain7.inv_chain[57] ;
 wire \thechain[0].chain7.inv_chain[58] ;
 wire \thechain[0].chain7.inv_chain[59] ;
 wire \thechain[0].chain7.inv_chain[5] ;
 wire \thechain[0].chain7.inv_chain[60] ;
 wire \thechain[0].chain7.inv_chain[61] ;
 wire \thechain[0].chain7.inv_chain[62] ;
 wire \thechain[0].chain7.inv_chain[63] ;
 wire \thechain[0].chain7.inv_chain[64] ;
 wire \thechain[0].chain7.inv_chain[65] ;
 wire \thechain[0].chain7.inv_chain[66] ;
 wire \thechain[0].chain7.inv_chain[67] ;
 wire \thechain[0].chain7.inv_chain[68] ;
 wire \thechain[0].chain7.inv_chain[69] ;
 wire \thechain[0].chain7.inv_chain[6] ;
 wire \thechain[0].chain7.inv_chain[70] ;
 wire \thechain[0].chain7.inv_chain[71] ;
 wire \thechain[0].chain7.inv_chain[72] ;
 wire \thechain[0].chain7.inv_chain[73] ;
 wire \thechain[0].chain7.inv_chain[74] ;
 wire \thechain[0].chain7.inv_chain[75] ;
 wire \thechain[0].chain7.inv_chain[76] ;
 wire \thechain[0].chain7.inv_chain[77] ;
 wire \thechain[0].chain7.inv_chain[78] ;
 wire \thechain[0].chain7.inv_chain[79] ;
 wire \thechain[0].chain7.inv_chain[7] ;
 wire \thechain[0].chain7.inv_chain[80] ;
 wire \thechain[0].chain7.inv_chain[81] ;
 wire \thechain[0].chain7.inv_chain[82] ;
 wire \thechain[0].chain7.inv_chain[83] ;
 wire \thechain[0].chain7.inv_chain[84] ;
 wire \thechain[0].chain7.inv_chain[85] ;
 wire \thechain[0].chain7.inv_chain[86] ;
 wire \thechain[0].chain7.inv_chain[87] ;
 wire \thechain[0].chain7.inv_chain[88] ;
 wire \thechain[0].chain7.inv_chain[89] ;
 wire \thechain[0].chain7.inv_chain[8] ;
 wire \thechain[0].chain7.inv_chain[90] ;
 wire \thechain[0].chain7.inv_chain[91] ;
 wire \thechain[0].chain7.inv_chain[92] ;
 wire \thechain[0].chain7.inv_chain[93] ;
 wire \thechain[0].chain7.inv_chain[94] ;
 wire \thechain[0].chain7.inv_chain[95] ;
 wire \thechain[0].chain7.inv_chain[96] ;
 wire \thechain[0].chain7.inv_chain[97] ;
 wire \thechain[0].chain7.inv_chain[98] ;
 wire \thechain[0].chain7.inv_chain[99] ;
 wire \thechain[0].chain7.inv_chain[9] ;
 wire \thechain[0].chain8.dout ;
 wire \thechain[0].chain8.inv_chain[0] ;
 wire \thechain[0].chain8.inv_chain[100] ;
 wire \thechain[0].chain8.inv_chain[101] ;
 wire \thechain[0].chain8.inv_chain[102] ;
 wire \thechain[0].chain8.inv_chain[103] ;
 wire \thechain[0].chain8.inv_chain[104] ;
 wire \thechain[0].chain8.inv_chain[105] ;
 wire \thechain[0].chain8.inv_chain[106] ;
 wire \thechain[0].chain8.inv_chain[107] ;
 wire \thechain[0].chain8.inv_chain[108] ;
 wire \thechain[0].chain8.inv_chain[109] ;
 wire \thechain[0].chain8.inv_chain[10] ;
 wire \thechain[0].chain8.inv_chain[110] ;
 wire \thechain[0].chain8.inv_chain[111] ;
 wire \thechain[0].chain8.inv_chain[112] ;
 wire \thechain[0].chain8.inv_chain[113] ;
 wire \thechain[0].chain8.inv_chain[114] ;
 wire \thechain[0].chain8.inv_chain[115] ;
 wire \thechain[0].chain8.inv_chain[116] ;
 wire \thechain[0].chain8.inv_chain[117] ;
 wire \thechain[0].chain8.inv_chain[118] ;
 wire \thechain[0].chain8.inv_chain[119] ;
 wire \thechain[0].chain8.inv_chain[11] ;
 wire \thechain[0].chain8.inv_chain[120] ;
 wire \thechain[0].chain8.inv_chain[121] ;
 wire \thechain[0].chain8.inv_chain[122] ;
 wire \thechain[0].chain8.inv_chain[123] ;
 wire \thechain[0].chain8.inv_chain[124] ;
 wire \thechain[0].chain8.inv_chain[125] ;
 wire \thechain[0].chain8.inv_chain[126] ;
 wire \thechain[0].chain8.inv_chain[127] ;
 wire \thechain[0].chain8.inv_chain[128] ;
 wire \thechain[0].chain8.inv_chain[129] ;
 wire \thechain[0].chain8.inv_chain[12] ;
 wire \thechain[0].chain8.inv_chain[130] ;
 wire \thechain[0].chain8.inv_chain[131] ;
 wire \thechain[0].chain8.inv_chain[132] ;
 wire \thechain[0].chain8.inv_chain[133] ;
 wire \thechain[0].chain8.inv_chain[134] ;
 wire \thechain[0].chain8.inv_chain[135] ;
 wire \thechain[0].chain8.inv_chain[136] ;
 wire \thechain[0].chain8.inv_chain[137] ;
 wire \thechain[0].chain8.inv_chain[138] ;
 wire \thechain[0].chain8.inv_chain[139] ;
 wire \thechain[0].chain8.inv_chain[13] ;
 wire \thechain[0].chain8.inv_chain[140] ;
 wire \thechain[0].chain8.inv_chain[141] ;
 wire \thechain[0].chain8.inv_chain[142] ;
 wire \thechain[0].chain8.inv_chain[143] ;
 wire \thechain[0].chain8.inv_chain[144] ;
 wire \thechain[0].chain8.inv_chain[145] ;
 wire \thechain[0].chain8.inv_chain[146] ;
 wire \thechain[0].chain8.inv_chain[147] ;
 wire \thechain[0].chain8.inv_chain[148] ;
 wire \thechain[0].chain8.inv_chain[149] ;
 wire \thechain[0].chain8.inv_chain[14] ;
 wire \thechain[0].chain8.inv_chain[150] ;
 wire \thechain[0].chain8.inv_chain[151] ;
 wire \thechain[0].chain8.inv_chain[152] ;
 wire \thechain[0].chain8.inv_chain[153] ;
 wire \thechain[0].chain8.inv_chain[154] ;
 wire \thechain[0].chain8.inv_chain[155] ;
 wire \thechain[0].chain8.inv_chain[156] ;
 wire \thechain[0].chain8.inv_chain[157] ;
 wire \thechain[0].chain8.inv_chain[158] ;
 wire \thechain[0].chain8.inv_chain[159] ;
 wire \thechain[0].chain8.inv_chain[15] ;
 wire \thechain[0].chain8.inv_chain[160] ;
 wire \thechain[0].chain8.inv_chain[161] ;
 wire \thechain[0].chain8.inv_chain[162] ;
 wire \thechain[0].chain8.inv_chain[163] ;
 wire \thechain[0].chain8.inv_chain[164] ;
 wire \thechain[0].chain8.inv_chain[165] ;
 wire \thechain[0].chain8.inv_chain[166] ;
 wire \thechain[0].chain8.inv_chain[167] ;
 wire \thechain[0].chain8.inv_chain[168] ;
 wire \thechain[0].chain8.inv_chain[169] ;
 wire \thechain[0].chain8.inv_chain[16] ;
 wire \thechain[0].chain8.inv_chain[170] ;
 wire \thechain[0].chain8.inv_chain[171] ;
 wire \thechain[0].chain8.inv_chain[172] ;
 wire \thechain[0].chain8.inv_chain[173] ;
 wire \thechain[0].chain8.inv_chain[174] ;
 wire \thechain[0].chain8.inv_chain[175] ;
 wire \thechain[0].chain8.inv_chain[176] ;
 wire \thechain[0].chain8.inv_chain[177] ;
 wire \thechain[0].chain8.inv_chain[178] ;
 wire \thechain[0].chain8.inv_chain[179] ;
 wire \thechain[0].chain8.inv_chain[17] ;
 wire \thechain[0].chain8.inv_chain[180] ;
 wire \thechain[0].chain8.inv_chain[181] ;
 wire \thechain[0].chain8.inv_chain[182] ;
 wire \thechain[0].chain8.inv_chain[183] ;
 wire \thechain[0].chain8.inv_chain[184] ;
 wire \thechain[0].chain8.inv_chain[185] ;
 wire \thechain[0].chain8.inv_chain[186] ;
 wire \thechain[0].chain8.inv_chain[187] ;
 wire \thechain[0].chain8.inv_chain[188] ;
 wire \thechain[0].chain8.inv_chain[189] ;
 wire \thechain[0].chain8.inv_chain[18] ;
 wire \thechain[0].chain8.inv_chain[190] ;
 wire \thechain[0].chain8.inv_chain[191] ;
 wire \thechain[0].chain8.inv_chain[192] ;
 wire \thechain[0].chain8.inv_chain[19] ;
 wire \thechain[0].chain8.inv_chain[1] ;
 wire \thechain[0].chain8.inv_chain[20] ;
 wire \thechain[0].chain8.inv_chain[21] ;
 wire \thechain[0].chain8.inv_chain[22] ;
 wire \thechain[0].chain8.inv_chain[23] ;
 wire \thechain[0].chain8.inv_chain[24] ;
 wire \thechain[0].chain8.inv_chain[25] ;
 wire \thechain[0].chain8.inv_chain[26] ;
 wire \thechain[0].chain8.inv_chain[27] ;
 wire \thechain[0].chain8.inv_chain[28] ;
 wire \thechain[0].chain8.inv_chain[29] ;
 wire \thechain[0].chain8.inv_chain[2] ;
 wire \thechain[0].chain8.inv_chain[30] ;
 wire \thechain[0].chain8.inv_chain[31] ;
 wire \thechain[0].chain8.inv_chain[32] ;
 wire \thechain[0].chain8.inv_chain[33] ;
 wire \thechain[0].chain8.inv_chain[34] ;
 wire \thechain[0].chain8.inv_chain[35] ;
 wire \thechain[0].chain8.inv_chain[36] ;
 wire \thechain[0].chain8.inv_chain[37] ;
 wire \thechain[0].chain8.inv_chain[38] ;
 wire \thechain[0].chain8.inv_chain[39] ;
 wire \thechain[0].chain8.inv_chain[3] ;
 wire \thechain[0].chain8.inv_chain[40] ;
 wire \thechain[0].chain8.inv_chain[41] ;
 wire \thechain[0].chain8.inv_chain[42] ;
 wire \thechain[0].chain8.inv_chain[43] ;
 wire \thechain[0].chain8.inv_chain[44] ;
 wire \thechain[0].chain8.inv_chain[45] ;
 wire \thechain[0].chain8.inv_chain[46] ;
 wire \thechain[0].chain8.inv_chain[47] ;
 wire \thechain[0].chain8.inv_chain[48] ;
 wire \thechain[0].chain8.inv_chain[49] ;
 wire \thechain[0].chain8.inv_chain[4] ;
 wire \thechain[0].chain8.inv_chain[50] ;
 wire \thechain[0].chain8.inv_chain[51] ;
 wire \thechain[0].chain8.inv_chain[52] ;
 wire \thechain[0].chain8.inv_chain[53] ;
 wire \thechain[0].chain8.inv_chain[54] ;
 wire \thechain[0].chain8.inv_chain[55] ;
 wire \thechain[0].chain8.inv_chain[56] ;
 wire \thechain[0].chain8.inv_chain[57] ;
 wire \thechain[0].chain8.inv_chain[58] ;
 wire \thechain[0].chain8.inv_chain[59] ;
 wire \thechain[0].chain8.inv_chain[5] ;
 wire \thechain[0].chain8.inv_chain[60] ;
 wire \thechain[0].chain8.inv_chain[61] ;
 wire \thechain[0].chain8.inv_chain[62] ;
 wire \thechain[0].chain8.inv_chain[63] ;
 wire \thechain[0].chain8.inv_chain[64] ;
 wire \thechain[0].chain8.inv_chain[65] ;
 wire \thechain[0].chain8.inv_chain[66] ;
 wire \thechain[0].chain8.inv_chain[67] ;
 wire \thechain[0].chain8.inv_chain[68] ;
 wire \thechain[0].chain8.inv_chain[69] ;
 wire \thechain[0].chain8.inv_chain[6] ;
 wire \thechain[0].chain8.inv_chain[70] ;
 wire \thechain[0].chain8.inv_chain[71] ;
 wire \thechain[0].chain8.inv_chain[72] ;
 wire \thechain[0].chain8.inv_chain[73] ;
 wire \thechain[0].chain8.inv_chain[74] ;
 wire \thechain[0].chain8.inv_chain[75] ;
 wire \thechain[0].chain8.inv_chain[76] ;
 wire \thechain[0].chain8.inv_chain[77] ;
 wire \thechain[0].chain8.inv_chain[78] ;
 wire \thechain[0].chain8.inv_chain[79] ;
 wire \thechain[0].chain8.inv_chain[7] ;
 wire \thechain[0].chain8.inv_chain[80] ;
 wire \thechain[0].chain8.inv_chain[81] ;
 wire \thechain[0].chain8.inv_chain[82] ;
 wire \thechain[0].chain8.inv_chain[83] ;
 wire \thechain[0].chain8.inv_chain[84] ;
 wire \thechain[0].chain8.inv_chain[85] ;
 wire \thechain[0].chain8.inv_chain[86] ;
 wire \thechain[0].chain8.inv_chain[87] ;
 wire \thechain[0].chain8.inv_chain[88] ;
 wire \thechain[0].chain8.inv_chain[89] ;
 wire \thechain[0].chain8.inv_chain[8] ;
 wire \thechain[0].chain8.inv_chain[90] ;
 wire \thechain[0].chain8.inv_chain[91] ;
 wire \thechain[0].chain8.inv_chain[92] ;
 wire \thechain[0].chain8.inv_chain[93] ;
 wire \thechain[0].chain8.inv_chain[94] ;
 wire \thechain[0].chain8.inv_chain[95] ;
 wire \thechain[0].chain8.inv_chain[96] ;
 wire \thechain[0].chain8.inv_chain[97] ;
 wire \thechain[0].chain8.inv_chain[98] ;
 wire \thechain[0].chain8.inv_chain[99] ;
 wire \thechain[0].chain8.inv_chain[9] ;
 wire \thechain[0].chain9.dout ;
 wire \thechain[0].chain9.inv_chain[0] ;
 wire \thechain[0].chain9.inv_chain[100] ;
 wire \thechain[0].chain9.inv_chain[101] ;
 wire \thechain[0].chain9.inv_chain[102] ;
 wire \thechain[0].chain9.inv_chain[103] ;
 wire \thechain[0].chain9.inv_chain[104] ;
 wire \thechain[0].chain9.inv_chain[105] ;
 wire \thechain[0].chain9.inv_chain[106] ;
 wire \thechain[0].chain9.inv_chain[107] ;
 wire \thechain[0].chain9.inv_chain[108] ;
 wire \thechain[0].chain9.inv_chain[109] ;
 wire \thechain[0].chain9.inv_chain[10] ;
 wire \thechain[0].chain9.inv_chain[110] ;
 wire \thechain[0].chain9.inv_chain[111] ;
 wire \thechain[0].chain9.inv_chain[112] ;
 wire \thechain[0].chain9.inv_chain[113] ;
 wire \thechain[0].chain9.inv_chain[114] ;
 wire \thechain[0].chain9.inv_chain[115] ;
 wire \thechain[0].chain9.inv_chain[116] ;
 wire \thechain[0].chain9.inv_chain[117] ;
 wire \thechain[0].chain9.inv_chain[118] ;
 wire \thechain[0].chain9.inv_chain[119] ;
 wire \thechain[0].chain9.inv_chain[11] ;
 wire \thechain[0].chain9.inv_chain[120] ;
 wire \thechain[0].chain9.inv_chain[121] ;
 wire \thechain[0].chain9.inv_chain[122] ;
 wire \thechain[0].chain9.inv_chain[123] ;
 wire \thechain[0].chain9.inv_chain[124] ;
 wire \thechain[0].chain9.inv_chain[125] ;
 wire \thechain[0].chain9.inv_chain[126] ;
 wire \thechain[0].chain9.inv_chain[127] ;
 wire \thechain[0].chain9.inv_chain[128] ;
 wire \thechain[0].chain9.inv_chain[129] ;
 wire \thechain[0].chain9.inv_chain[12] ;
 wire \thechain[0].chain9.inv_chain[130] ;
 wire \thechain[0].chain9.inv_chain[131] ;
 wire \thechain[0].chain9.inv_chain[132] ;
 wire \thechain[0].chain9.inv_chain[133] ;
 wire \thechain[0].chain9.inv_chain[134] ;
 wire \thechain[0].chain9.inv_chain[135] ;
 wire \thechain[0].chain9.inv_chain[136] ;
 wire \thechain[0].chain9.inv_chain[137] ;
 wire \thechain[0].chain9.inv_chain[138] ;
 wire \thechain[0].chain9.inv_chain[139] ;
 wire \thechain[0].chain9.inv_chain[13] ;
 wire \thechain[0].chain9.inv_chain[140] ;
 wire \thechain[0].chain9.inv_chain[141] ;
 wire \thechain[0].chain9.inv_chain[142] ;
 wire \thechain[0].chain9.inv_chain[143] ;
 wire \thechain[0].chain9.inv_chain[144] ;
 wire \thechain[0].chain9.inv_chain[145] ;
 wire \thechain[0].chain9.inv_chain[146] ;
 wire \thechain[0].chain9.inv_chain[147] ;
 wire \thechain[0].chain9.inv_chain[148] ;
 wire \thechain[0].chain9.inv_chain[149] ;
 wire \thechain[0].chain9.inv_chain[14] ;
 wire \thechain[0].chain9.inv_chain[150] ;
 wire \thechain[0].chain9.inv_chain[151] ;
 wire \thechain[0].chain9.inv_chain[152] ;
 wire \thechain[0].chain9.inv_chain[153] ;
 wire \thechain[0].chain9.inv_chain[154] ;
 wire \thechain[0].chain9.inv_chain[155] ;
 wire \thechain[0].chain9.inv_chain[156] ;
 wire \thechain[0].chain9.inv_chain[157] ;
 wire \thechain[0].chain9.inv_chain[158] ;
 wire \thechain[0].chain9.inv_chain[159] ;
 wire \thechain[0].chain9.inv_chain[15] ;
 wire \thechain[0].chain9.inv_chain[160] ;
 wire \thechain[0].chain9.inv_chain[161] ;
 wire \thechain[0].chain9.inv_chain[162] ;
 wire \thechain[0].chain9.inv_chain[163] ;
 wire \thechain[0].chain9.inv_chain[164] ;
 wire \thechain[0].chain9.inv_chain[165] ;
 wire \thechain[0].chain9.inv_chain[166] ;
 wire \thechain[0].chain9.inv_chain[167] ;
 wire \thechain[0].chain9.inv_chain[168] ;
 wire \thechain[0].chain9.inv_chain[169] ;
 wire \thechain[0].chain9.inv_chain[16] ;
 wire \thechain[0].chain9.inv_chain[170] ;
 wire \thechain[0].chain9.inv_chain[171] ;
 wire \thechain[0].chain9.inv_chain[172] ;
 wire \thechain[0].chain9.inv_chain[173] ;
 wire \thechain[0].chain9.inv_chain[174] ;
 wire \thechain[0].chain9.inv_chain[175] ;
 wire \thechain[0].chain9.inv_chain[176] ;
 wire \thechain[0].chain9.inv_chain[177] ;
 wire \thechain[0].chain9.inv_chain[178] ;
 wire \thechain[0].chain9.inv_chain[179] ;
 wire \thechain[0].chain9.inv_chain[17] ;
 wire \thechain[0].chain9.inv_chain[180] ;
 wire \thechain[0].chain9.inv_chain[181] ;
 wire \thechain[0].chain9.inv_chain[182] ;
 wire \thechain[0].chain9.inv_chain[183] ;
 wire \thechain[0].chain9.inv_chain[184] ;
 wire \thechain[0].chain9.inv_chain[185] ;
 wire \thechain[0].chain9.inv_chain[186] ;
 wire \thechain[0].chain9.inv_chain[187] ;
 wire \thechain[0].chain9.inv_chain[188] ;
 wire \thechain[0].chain9.inv_chain[189] ;
 wire \thechain[0].chain9.inv_chain[18] ;
 wire \thechain[0].chain9.inv_chain[190] ;
 wire \thechain[0].chain9.inv_chain[191] ;
 wire \thechain[0].chain9.inv_chain[192] ;
 wire \thechain[0].chain9.inv_chain[193] ;
 wire \thechain[0].chain9.inv_chain[194] ;
 wire \thechain[0].chain9.inv_chain[195] ;
 wire \thechain[0].chain9.inv_chain[196] ;
 wire \thechain[0].chain9.inv_chain[197] ;
 wire \thechain[0].chain9.inv_chain[198] ;
 wire \thechain[0].chain9.inv_chain[199] ;
 wire \thechain[0].chain9.inv_chain[19] ;
 wire \thechain[0].chain9.inv_chain[1] ;
 wire \thechain[0].chain9.inv_chain[200] ;
 wire \thechain[0].chain9.inv_chain[201] ;
 wire \thechain[0].chain9.inv_chain[202] ;
 wire \thechain[0].chain9.inv_chain[203] ;
 wire \thechain[0].chain9.inv_chain[204] ;
 wire \thechain[0].chain9.inv_chain[205] ;
 wire \thechain[0].chain9.inv_chain[206] ;
 wire \thechain[0].chain9.inv_chain[207] ;
 wire \thechain[0].chain9.inv_chain[208] ;
 wire \thechain[0].chain9.inv_chain[209] ;
 wire \thechain[0].chain9.inv_chain[20] ;
 wire \thechain[0].chain9.inv_chain[210] ;
 wire \thechain[0].chain9.inv_chain[211] ;
 wire \thechain[0].chain9.inv_chain[212] ;
 wire \thechain[0].chain9.inv_chain[213] ;
 wire \thechain[0].chain9.inv_chain[214] ;
 wire \thechain[0].chain9.inv_chain[215] ;
 wire \thechain[0].chain9.inv_chain[216] ;
 wire \thechain[0].chain9.inv_chain[217] ;
 wire \thechain[0].chain9.inv_chain[218] ;
 wire \thechain[0].chain9.inv_chain[219] ;
 wire \thechain[0].chain9.inv_chain[21] ;
 wire \thechain[0].chain9.inv_chain[220] ;
 wire \thechain[0].chain9.inv_chain[221] ;
 wire \thechain[0].chain9.inv_chain[222] ;
 wire \thechain[0].chain9.inv_chain[223] ;
 wire \thechain[0].chain9.inv_chain[224] ;
 wire \thechain[0].chain9.inv_chain[225] ;
 wire \thechain[0].chain9.inv_chain[226] ;
 wire \thechain[0].chain9.inv_chain[227] ;
 wire \thechain[0].chain9.inv_chain[228] ;
 wire \thechain[0].chain9.inv_chain[229] ;
 wire \thechain[0].chain9.inv_chain[22] ;
 wire \thechain[0].chain9.inv_chain[230] ;
 wire \thechain[0].chain9.inv_chain[231] ;
 wire \thechain[0].chain9.inv_chain[232] ;
 wire \thechain[0].chain9.inv_chain[233] ;
 wire \thechain[0].chain9.inv_chain[234] ;
 wire \thechain[0].chain9.inv_chain[235] ;
 wire \thechain[0].chain9.inv_chain[236] ;
 wire \thechain[0].chain9.inv_chain[237] ;
 wire \thechain[0].chain9.inv_chain[238] ;
 wire \thechain[0].chain9.inv_chain[239] ;
 wire \thechain[0].chain9.inv_chain[23] ;
 wire \thechain[0].chain9.inv_chain[240] ;
 wire \thechain[0].chain9.inv_chain[241] ;
 wire \thechain[0].chain9.inv_chain[242] ;
 wire \thechain[0].chain9.inv_chain[243] ;
 wire \thechain[0].chain9.inv_chain[244] ;
 wire \thechain[0].chain9.inv_chain[245] ;
 wire \thechain[0].chain9.inv_chain[246] ;
 wire \thechain[0].chain9.inv_chain[247] ;
 wire \thechain[0].chain9.inv_chain[248] ;
 wire \thechain[0].chain9.inv_chain[249] ;
 wire \thechain[0].chain9.inv_chain[24] ;
 wire \thechain[0].chain9.inv_chain[250] ;
 wire \thechain[0].chain9.inv_chain[251] ;
 wire \thechain[0].chain9.inv_chain[252] ;
 wire \thechain[0].chain9.inv_chain[253] ;
 wire \thechain[0].chain9.inv_chain[254] ;
 wire \thechain[0].chain9.inv_chain[255] ;
 wire \thechain[0].chain9.inv_chain[256] ;
 wire \thechain[0].chain9.inv_chain[25] ;
 wire \thechain[0].chain9.inv_chain[26] ;
 wire \thechain[0].chain9.inv_chain[27] ;
 wire \thechain[0].chain9.inv_chain[28] ;
 wire \thechain[0].chain9.inv_chain[29] ;
 wire \thechain[0].chain9.inv_chain[2] ;
 wire \thechain[0].chain9.inv_chain[30] ;
 wire \thechain[0].chain9.inv_chain[31] ;
 wire \thechain[0].chain9.inv_chain[32] ;
 wire \thechain[0].chain9.inv_chain[33] ;
 wire \thechain[0].chain9.inv_chain[34] ;
 wire \thechain[0].chain9.inv_chain[35] ;
 wire \thechain[0].chain9.inv_chain[36] ;
 wire \thechain[0].chain9.inv_chain[37] ;
 wire \thechain[0].chain9.inv_chain[38] ;
 wire \thechain[0].chain9.inv_chain[39] ;
 wire \thechain[0].chain9.inv_chain[3] ;
 wire \thechain[0].chain9.inv_chain[40] ;
 wire \thechain[0].chain9.inv_chain[41] ;
 wire \thechain[0].chain9.inv_chain[42] ;
 wire \thechain[0].chain9.inv_chain[43] ;
 wire \thechain[0].chain9.inv_chain[44] ;
 wire \thechain[0].chain9.inv_chain[45] ;
 wire \thechain[0].chain9.inv_chain[46] ;
 wire \thechain[0].chain9.inv_chain[47] ;
 wire \thechain[0].chain9.inv_chain[48] ;
 wire \thechain[0].chain9.inv_chain[49] ;
 wire \thechain[0].chain9.inv_chain[4] ;
 wire \thechain[0].chain9.inv_chain[50] ;
 wire \thechain[0].chain9.inv_chain[51] ;
 wire \thechain[0].chain9.inv_chain[52] ;
 wire \thechain[0].chain9.inv_chain[53] ;
 wire \thechain[0].chain9.inv_chain[54] ;
 wire \thechain[0].chain9.inv_chain[55] ;
 wire \thechain[0].chain9.inv_chain[56] ;
 wire \thechain[0].chain9.inv_chain[57] ;
 wire \thechain[0].chain9.inv_chain[58] ;
 wire \thechain[0].chain9.inv_chain[59] ;
 wire \thechain[0].chain9.inv_chain[5] ;
 wire \thechain[0].chain9.inv_chain[60] ;
 wire \thechain[0].chain9.inv_chain[61] ;
 wire \thechain[0].chain9.inv_chain[62] ;
 wire \thechain[0].chain9.inv_chain[63] ;
 wire \thechain[0].chain9.inv_chain[64] ;
 wire \thechain[0].chain9.inv_chain[65] ;
 wire \thechain[0].chain9.inv_chain[66] ;
 wire \thechain[0].chain9.inv_chain[67] ;
 wire \thechain[0].chain9.inv_chain[68] ;
 wire \thechain[0].chain9.inv_chain[69] ;
 wire \thechain[0].chain9.inv_chain[6] ;
 wire \thechain[0].chain9.inv_chain[70] ;
 wire \thechain[0].chain9.inv_chain[71] ;
 wire \thechain[0].chain9.inv_chain[72] ;
 wire \thechain[0].chain9.inv_chain[73] ;
 wire \thechain[0].chain9.inv_chain[74] ;
 wire \thechain[0].chain9.inv_chain[75] ;
 wire \thechain[0].chain9.inv_chain[76] ;
 wire \thechain[0].chain9.inv_chain[77] ;
 wire \thechain[0].chain9.inv_chain[78] ;
 wire \thechain[0].chain9.inv_chain[79] ;
 wire \thechain[0].chain9.inv_chain[7] ;
 wire \thechain[0].chain9.inv_chain[80] ;
 wire \thechain[0].chain9.inv_chain[81] ;
 wire \thechain[0].chain9.inv_chain[82] ;
 wire \thechain[0].chain9.inv_chain[83] ;
 wire \thechain[0].chain9.inv_chain[84] ;
 wire \thechain[0].chain9.inv_chain[85] ;
 wire \thechain[0].chain9.inv_chain[86] ;
 wire \thechain[0].chain9.inv_chain[87] ;
 wire \thechain[0].chain9.inv_chain[88] ;
 wire \thechain[0].chain9.inv_chain[89] ;
 wire \thechain[0].chain9.inv_chain[8] ;
 wire \thechain[0].chain9.inv_chain[90] ;
 wire \thechain[0].chain9.inv_chain[91] ;
 wire \thechain[0].chain9.inv_chain[92] ;
 wire \thechain[0].chain9.inv_chain[93] ;
 wire \thechain[0].chain9.inv_chain[94] ;
 wire \thechain[0].chain9.inv_chain[95] ;
 wire \thechain[0].chain9.inv_chain[96] ;
 wire \thechain[0].chain9.inv_chain[97] ;
 wire \thechain[0].chain9.inv_chain[98] ;
 wire \thechain[0].chain9.inv_chain[99] ;
 wire \thechain[0].chain9.inv_chain[9] ;
 wire \thechain[1].chain1.dout ;
 wire \thechain[1].chain1.inv_chain[0] ;
 wire \thechain[1].chain1.inv_chain[1] ;
 wire \thechain[1].chain1.inv_chain[2] ;
 wire \thechain[1].chain2.dout ;
 wire \thechain[1].chain2.inv_chain[0] ;
 wire \thechain[1].chain2.inv_chain[1] ;
 wire \thechain[1].chain2.inv_chain[2] ;
 wire \thechain[1].chain2.inv_chain[3] ;
 wire \thechain[1].chain2.inv_chain[4] ;
 wire \thechain[1].chain3.dout ;
 wire \thechain[1].chain3.inv_chain[0] ;
 wire \thechain[1].chain3.inv_chain[1] ;
 wire \thechain[1].chain3.inv_chain[2] ;
 wire \thechain[1].chain3.inv_chain[3] ;
 wire \thechain[1].chain3.inv_chain[4] ;
 wire \thechain[1].chain3.inv_chain[5] ;
 wire \thechain[1].chain3.inv_chain[6] ;
 wire \thechain[1].chain3.inv_chain[7] ;
 wire \thechain[1].chain3.inv_chain[8] ;
 wire \thechain[1].chain4.dout ;
 wire \thechain[1].chain4.inv_chain[0] ;
 wire \thechain[1].chain4.inv_chain[10] ;
 wire \thechain[1].chain4.inv_chain[11] ;
 wire \thechain[1].chain4.inv_chain[12] ;
 wire \thechain[1].chain4.inv_chain[13] ;
 wire \thechain[1].chain4.inv_chain[14] ;
 wire \thechain[1].chain4.inv_chain[15] ;
 wire \thechain[1].chain4.inv_chain[16] ;
 wire \thechain[1].chain4.inv_chain[1] ;
 wire \thechain[1].chain4.inv_chain[2] ;
 wire \thechain[1].chain4.inv_chain[3] ;
 wire \thechain[1].chain4.inv_chain[4] ;
 wire \thechain[1].chain4.inv_chain[5] ;
 wire \thechain[1].chain4.inv_chain[6] ;
 wire \thechain[1].chain4.inv_chain[7] ;
 wire \thechain[1].chain4.inv_chain[8] ;
 wire \thechain[1].chain4.inv_chain[9] ;
 wire \thechain[1].chain5.dout ;
 wire \thechain[1].chain5.inv_chain[0] ;
 wire \thechain[1].chain5.inv_chain[10] ;
 wire \thechain[1].chain5.inv_chain[11] ;
 wire \thechain[1].chain5.inv_chain[12] ;
 wire \thechain[1].chain5.inv_chain[13] ;
 wire \thechain[1].chain5.inv_chain[14] ;
 wire \thechain[1].chain5.inv_chain[15] ;
 wire \thechain[1].chain5.inv_chain[16] ;
 wire \thechain[1].chain5.inv_chain[17] ;
 wire \thechain[1].chain5.inv_chain[18] ;
 wire \thechain[1].chain5.inv_chain[19] ;
 wire \thechain[1].chain5.inv_chain[1] ;
 wire \thechain[1].chain5.inv_chain[20] ;
 wire \thechain[1].chain5.inv_chain[21] ;
 wire \thechain[1].chain5.inv_chain[22] ;
 wire \thechain[1].chain5.inv_chain[23] ;
 wire \thechain[1].chain5.inv_chain[24] ;
 wire \thechain[1].chain5.inv_chain[25] ;
 wire \thechain[1].chain5.inv_chain[26] ;
 wire \thechain[1].chain5.inv_chain[27] ;
 wire \thechain[1].chain5.inv_chain[28] ;
 wire \thechain[1].chain5.inv_chain[29] ;
 wire \thechain[1].chain5.inv_chain[2] ;
 wire \thechain[1].chain5.inv_chain[30] ;
 wire \thechain[1].chain5.inv_chain[31] ;
 wire \thechain[1].chain5.inv_chain[32] ;
 wire \thechain[1].chain5.inv_chain[3] ;
 wire \thechain[1].chain5.inv_chain[4] ;
 wire \thechain[1].chain5.inv_chain[5] ;
 wire \thechain[1].chain5.inv_chain[6] ;
 wire \thechain[1].chain5.inv_chain[7] ;
 wire \thechain[1].chain5.inv_chain[8] ;
 wire \thechain[1].chain5.inv_chain[9] ;
 wire \thechain[1].chain6.dout ;
 wire \thechain[1].chain6.inv_chain[0] ;
 wire \thechain[1].chain6.inv_chain[10] ;
 wire \thechain[1].chain6.inv_chain[11] ;
 wire \thechain[1].chain6.inv_chain[12] ;
 wire \thechain[1].chain6.inv_chain[13] ;
 wire \thechain[1].chain6.inv_chain[14] ;
 wire \thechain[1].chain6.inv_chain[15] ;
 wire \thechain[1].chain6.inv_chain[16] ;
 wire \thechain[1].chain6.inv_chain[17] ;
 wire \thechain[1].chain6.inv_chain[18] ;
 wire \thechain[1].chain6.inv_chain[19] ;
 wire \thechain[1].chain6.inv_chain[1] ;
 wire \thechain[1].chain6.inv_chain[20] ;
 wire \thechain[1].chain6.inv_chain[21] ;
 wire \thechain[1].chain6.inv_chain[22] ;
 wire \thechain[1].chain6.inv_chain[23] ;
 wire \thechain[1].chain6.inv_chain[24] ;
 wire \thechain[1].chain6.inv_chain[25] ;
 wire \thechain[1].chain6.inv_chain[26] ;
 wire \thechain[1].chain6.inv_chain[27] ;
 wire \thechain[1].chain6.inv_chain[28] ;
 wire \thechain[1].chain6.inv_chain[29] ;
 wire \thechain[1].chain6.inv_chain[2] ;
 wire \thechain[1].chain6.inv_chain[30] ;
 wire \thechain[1].chain6.inv_chain[31] ;
 wire \thechain[1].chain6.inv_chain[32] ;
 wire \thechain[1].chain6.inv_chain[33] ;
 wire \thechain[1].chain6.inv_chain[34] ;
 wire \thechain[1].chain6.inv_chain[35] ;
 wire \thechain[1].chain6.inv_chain[36] ;
 wire \thechain[1].chain6.inv_chain[37] ;
 wire \thechain[1].chain6.inv_chain[38] ;
 wire \thechain[1].chain6.inv_chain[39] ;
 wire \thechain[1].chain6.inv_chain[3] ;
 wire \thechain[1].chain6.inv_chain[40] ;
 wire \thechain[1].chain6.inv_chain[41] ;
 wire \thechain[1].chain6.inv_chain[42] ;
 wire \thechain[1].chain6.inv_chain[43] ;
 wire \thechain[1].chain6.inv_chain[44] ;
 wire \thechain[1].chain6.inv_chain[45] ;
 wire \thechain[1].chain6.inv_chain[46] ;
 wire \thechain[1].chain6.inv_chain[47] ;
 wire \thechain[1].chain6.inv_chain[48] ;
 wire \thechain[1].chain6.inv_chain[49] ;
 wire \thechain[1].chain6.inv_chain[4] ;
 wire \thechain[1].chain6.inv_chain[50] ;
 wire \thechain[1].chain6.inv_chain[51] ;
 wire \thechain[1].chain6.inv_chain[52] ;
 wire \thechain[1].chain6.inv_chain[53] ;
 wire \thechain[1].chain6.inv_chain[54] ;
 wire \thechain[1].chain6.inv_chain[55] ;
 wire \thechain[1].chain6.inv_chain[56] ;
 wire \thechain[1].chain6.inv_chain[57] ;
 wire \thechain[1].chain6.inv_chain[58] ;
 wire \thechain[1].chain6.inv_chain[59] ;
 wire \thechain[1].chain6.inv_chain[5] ;
 wire \thechain[1].chain6.inv_chain[60] ;
 wire \thechain[1].chain6.inv_chain[61] ;
 wire \thechain[1].chain6.inv_chain[62] ;
 wire \thechain[1].chain6.inv_chain[63] ;
 wire \thechain[1].chain6.inv_chain[64] ;
 wire \thechain[1].chain6.inv_chain[6] ;
 wire \thechain[1].chain6.inv_chain[7] ;
 wire \thechain[1].chain6.inv_chain[8] ;
 wire \thechain[1].chain6.inv_chain[9] ;
 wire \thechain[1].chain7.dout ;
 wire \thechain[1].chain7.inv_chain[0] ;
 wire \thechain[1].chain7.inv_chain[100] ;
 wire \thechain[1].chain7.inv_chain[101] ;
 wire \thechain[1].chain7.inv_chain[102] ;
 wire \thechain[1].chain7.inv_chain[103] ;
 wire \thechain[1].chain7.inv_chain[104] ;
 wire \thechain[1].chain7.inv_chain[105] ;
 wire \thechain[1].chain7.inv_chain[106] ;
 wire \thechain[1].chain7.inv_chain[107] ;
 wire \thechain[1].chain7.inv_chain[108] ;
 wire \thechain[1].chain7.inv_chain[109] ;
 wire \thechain[1].chain7.inv_chain[10] ;
 wire \thechain[1].chain7.inv_chain[110] ;
 wire \thechain[1].chain7.inv_chain[111] ;
 wire \thechain[1].chain7.inv_chain[112] ;
 wire \thechain[1].chain7.inv_chain[113] ;
 wire \thechain[1].chain7.inv_chain[114] ;
 wire \thechain[1].chain7.inv_chain[115] ;
 wire \thechain[1].chain7.inv_chain[116] ;
 wire \thechain[1].chain7.inv_chain[117] ;
 wire \thechain[1].chain7.inv_chain[118] ;
 wire \thechain[1].chain7.inv_chain[119] ;
 wire \thechain[1].chain7.inv_chain[11] ;
 wire \thechain[1].chain7.inv_chain[120] ;
 wire \thechain[1].chain7.inv_chain[121] ;
 wire \thechain[1].chain7.inv_chain[122] ;
 wire \thechain[1].chain7.inv_chain[123] ;
 wire \thechain[1].chain7.inv_chain[124] ;
 wire \thechain[1].chain7.inv_chain[125] ;
 wire \thechain[1].chain7.inv_chain[126] ;
 wire \thechain[1].chain7.inv_chain[127] ;
 wire \thechain[1].chain7.inv_chain[128] ;
 wire \thechain[1].chain7.inv_chain[12] ;
 wire \thechain[1].chain7.inv_chain[13] ;
 wire \thechain[1].chain7.inv_chain[14] ;
 wire \thechain[1].chain7.inv_chain[15] ;
 wire \thechain[1].chain7.inv_chain[16] ;
 wire \thechain[1].chain7.inv_chain[17] ;
 wire \thechain[1].chain7.inv_chain[18] ;
 wire \thechain[1].chain7.inv_chain[19] ;
 wire \thechain[1].chain7.inv_chain[1] ;
 wire \thechain[1].chain7.inv_chain[20] ;
 wire \thechain[1].chain7.inv_chain[21] ;
 wire \thechain[1].chain7.inv_chain[22] ;
 wire \thechain[1].chain7.inv_chain[23] ;
 wire \thechain[1].chain7.inv_chain[24] ;
 wire \thechain[1].chain7.inv_chain[25] ;
 wire \thechain[1].chain7.inv_chain[26] ;
 wire \thechain[1].chain7.inv_chain[27] ;
 wire \thechain[1].chain7.inv_chain[28] ;
 wire \thechain[1].chain7.inv_chain[29] ;
 wire \thechain[1].chain7.inv_chain[2] ;
 wire \thechain[1].chain7.inv_chain[30] ;
 wire \thechain[1].chain7.inv_chain[31] ;
 wire \thechain[1].chain7.inv_chain[32] ;
 wire \thechain[1].chain7.inv_chain[33] ;
 wire \thechain[1].chain7.inv_chain[34] ;
 wire \thechain[1].chain7.inv_chain[35] ;
 wire \thechain[1].chain7.inv_chain[36] ;
 wire \thechain[1].chain7.inv_chain[37] ;
 wire \thechain[1].chain7.inv_chain[38] ;
 wire \thechain[1].chain7.inv_chain[39] ;
 wire \thechain[1].chain7.inv_chain[3] ;
 wire \thechain[1].chain7.inv_chain[40] ;
 wire \thechain[1].chain7.inv_chain[41] ;
 wire \thechain[1].chain7.inv_chain[42] ;
 wire \thechain[1].chain7.inv_chain[43] ;
 wire \thechain[1].chain7.inv_chain[44] ;
 wire \thechain[1].chain7.inv_chain[45] ;
 wire \thechain[1].chain7.inv_chain[46] ;
 wire \thechain[1].chain7.inv_chain[47] ;
 wire \thechain[1].chain7.inv_chain[48] ;
 wire \thechain[1].chain7.inv_chain[49] ;
 wire \thechain[1].chain7.inv_chain[4] ;
 wire \thechain[1].chain7.inv_chain[50] ;
 wire \thechain[1].chain7.inv_chain[51] ;
 wire \thechain[1].chain7.inv_chain[52] ;
 wire \thechain[1].chain7.inv_chain[53] ;
 wire \thechain[1].chain7.inv_chain[54] ;
 wire \thechain[1].chain7.inv_chain[55] ;
 wire \thechain[1].chain7.inv_chain[56] ;
 wire \thechain[1].chain7.inv_chain[57] ;
 wire \thechain[1].chain7.inv_chain[58] ;
 wire \thechain[1].chain7.inv_chain[59] ;
 wire \thechain[1].chain7.inv_chain[5] ;
 wire \thechain[1].chain7.inv_chain[60] ;
 wire \thechain[1].chain7.inv_chain[61] ;
 wire \thechain[1].chain7.inv_chain[62] ;
 wire \thechain[1].chain7.inv_chain[63] ;
 wire \thechain[1].chain7.inv_chain[64] ;
 wire \thechain[1].chain7.inv_chain[65] ;
 wire \thechain[1].chain7.inv_chain[66] ;
 wire \thechain[1].chain7.inv_chain[67] ;
 wire \thechain[1].chain7.inv_chain[68] ;
 wire \thechain[1].chain7.inv_chain[69] ;
 wire \thechain[1].chain7.inv_chain[6] ;
 wire \thechain[1].chain7.inv_chain[70] ;
 wire \thechain[1].chain7.inv_chain[71] ;
 wire \thechain[1].chain7.inv_chain[72] ;
 wire \thechain[1].chain7.inv_chain[73] ;
 wire \thechain[1].chain7.inv_chain[74] ;
 wire \thechain[1].chain7.inv_chain[75] ;
 wire \thechain[1].chain7.inv_chain[76] ;
 wire \thechain[1].chain7.inv_chain[77] ;
 wire \thechain[1].chain7.inv_chain[78] ;
 wire \thechain[1].chain7.inv_chain[79] ;
 wire \thechain[1].chain7.inv_chain[7] ;
 wire \thechain[1].chain7.inv_chain[80] ;
 wire \thechain[1].chain7.inv_chain[81] ;
 wire \thechain[1].chain7.inv_chain[82] ;
 wire \thechain[1].chain7.inv_chain[83] ;
 wire \thechain[1].chain7.inv_chain[84] ;
 wire \thechain[1].chain7.inv_chain[85] ;
 wire \thechain[1].chain7.inv_chain[86] ;
 wire \thechain[1].chain7.inv_chain[87] ;
 wire \thechain[1].chain7.inv_chain[88] ;
 wire \thechain[1].chain7.inv_chain[89] ;
 wire \thechain[1].chain7.inv_chain[8] ;
 wire \thechain[1].chain7.inv_chain[90] ;
 wire \thechain[1].chain7.inv_chain[91] ;
 wire \thechain[1].chain7.inv_chain[92] ;
 wire \thechain[1].chain7.inv_chain[93] ;
 wire \thechain[1].chain7.inv_chain[94] ;
 wire \thechain[1].chain7.inv_chain[95] ;
 wire \thechain[1].chain7.inv_chain[96] ;
 wire \thechain[1].chain7.inv_chain[97] ;
 wire \thechain[1].chain7.inv_chain[98] ;
 wire \thechain[1].chain7.inv_chain[99] ;
 wire \thechain[1].chain7.inv_chain[9] ;
 wire \thechain[1].chain8.dout ;
 wire \thechain[1].chain8.inv_chain[0] ;
 wire \thechain[1].chain8.inv_chain[100] ;
 wire \thechain[1].chain8.inv_chain[101] ;
 wire \thechain[1].chain8.inv_chain[102] ;
 wire \thechain[1].chain8.inv_chain[103] ;
 wire \thechain[1].chain8.inv_chain[104] ;
 wire \thechain[1].chain8.inv_chain[105] ;
 wire \thechain[1].chain8.inv_chain[106] ;
 wire \thechain[1].chain8.inv_chain[107] ;
 wire \thechain[1].chain8.inv_chain[108] ;
 wire \thechain[1].chain8.inv_chain[109] ;
 wire \thechain[1].chain8.inv_chain[10] ;
 wire \thechain[1].chain8.inv_chain[110] ;
 wire \thechain[1].chain8.inv_chain[111] ;
 wire \thechain[1].chain8.inv_chain[112] ;
 wire \thechain[1].chain8.inv_chain[113] ;
 wire \thechain[1].chain8.inv_chain[114] ;
 wire \thechain[1].chain8.inv_chain[115] ;
 wire \thechain[1].chain8.inv_chain[116] ;
 wire \thechain[1].chain8.inv_chain[117] ;
 wire \thechain[1].chain8.inv_chain[118] ;
 wire \thechain[1].chain8.inv_chain[119] ;
 wire \thechain[1].chain8.inv_chain[11] ;
 wire \thechain[1].chain8.inv_chain[120] ;
 wire \thechain[1].chain8.inv_chain[121] ;
 wire \thechain[1].chain8.inv_chain[122] ;
 wire \thechain[1].chain8.inv_chain[123] ;
 wire \thechain[1].chain8.inv_chain[124] ;
 wire \thechain[1].chain8.inv_chain[125] ;
 wire \thechain[1].chain8.inv_chain[126] ;
 wire \thechain[1].chain8.inv_chain[127] ;
 wire \thechain[1].chain8.inv_chain[128] ;
 wire \thechain[1].chain8.inv_chain[129] ;
 wire \thechain[1].chain8.inv_chain[12] ;
 wire \thechain[1].chain8.inv_chain[130] ;
 wire \thechain[1].chain8.inv_chain[131] ;
 wire \thechain[1].chain8.inv_chain[132] ;
 wire \thechain[1].chain8.inv_chain[133] ;
 wire \thechain[1].chain8.inv_chain[134] ;
 wire \thechain[1].chain8.inv_chain[135] ;
 wire \thechain[1].chain8.inv_chain[136] ;
 wire \thechain[1].chain8.inv_chain[137] ;
 wire \thechain[1].chain8.inv_chain[138] ;
 wire \thechain[1].chain8.inv_chain[139] ;
 wire \thechain[1].chain8.inv_chain[13] ;
 wire \thechain[1].chain8.inv_chain[140] ;
 wire \thechain[1].chain8.inv_chain[141] ;
 wire \thechain[1].chain8.inv_chain[142] ;
 wire \thechain[1].chain8.inv_chain[143] ;
 wire \thechain[1].chain8.inv_chain[144] ;
 wire \thechain[1].chain8.inv_chain[145] ;
 wire \thechain[1].chain8.inv_chain[146] ;
 wire \thechain[1].chain8.inv_chain[147] ;
 wire \thechain[1].chain8.inv_chain[148] ;
 wire \thechain[1].chain8.inv_chain[149] ;
 wire \thechain[1].chain8.inv_chain[14] ;
 wire \thechain[1].chain8.inv_chain[150] ;
 wire \thechain[1].chain8.inv_chain[151] ;
 wire \thechain[1].chain8.inv_chain[152] ;
 wire \thechain[1].chain8.inv_chain[153] ;
 wire \thechain[1].chain8.inv_chain[154] ;
 wire \thechain[1].chain8.inv_chain[155] ;
 wire \thechain[1].chain8.inv_chain[156] ;
 wire \thechain[1].chain8.inv_chain[157] ;
 wire \thechain[1].chain8.inv_chain[158] ;
 wire \thechain[1].chain8.inv_chain[159] ;
 wire \thechain[1].chain8.inv_chain[15] ;
 wire \thechain[1].chain8.inv_chain[160] ;
 wire \thechain[1].chain8.inv_chain[161] ;
 wire \thechain[1].chain8.inv_chain[162] ;
 wire \thechain[1].chain8.inv_chain[163] ;
 wire \thechain[1].chain8.inv_chain[164] ;
 wire \thechain[1].chain8.inv_chain[165] ;
 wire \thechain[1].chain8.inv_chain[166] ;
 wire \thechain[1].chain8.inv_chain[167] ;
 wire \thechain[1].chain8.inv_chain[168] ;
 wire \thechain[1].chain8.inv_chain[169] ;
 wire \thechain[1].chain8.inv_chain[16] ;
 wire \thechain[1].chain8.inv_chain[170] ;
 wire \thechain[1].chain8.inv_chain[171] ;
 wire \thechain[1].chain8.inv_chain[172] ;
 wire \thechain[1].chain8.inv_chain[173] ;
 wire \thechain[1].chain8.inv_chain[174] ;
 wire \thechain[1].chain8.inv_chain[175] ;
 wire \thechain[1].chain8.inv_chain[176] ;
 wire \thechain[1].chain8.inv_chain[177] ;
 wire \thechain[1].chain8.inv_chain[178] ;
 wire \thechain[1].chain8.inv_chain[179] ;
 wire \thechain[1].chain8.inv_chain[17] ;
 wire \thechain[1].chain8.inv_chain[180] ;
 wire \thechain[1].chain8.inv_chain[181] ;
 wire \thechain[1].chain8.inv_chain[182] ;
 wire \thechain[1].chain8.inv_chain[183] ;
 wire \thechain[1].chain8.inv_chain[184] ;
 wire \thechain[1].chain8.inv_chain[185] ;
 wire \thechain[1].chain8.inv_chain[186] ;
 wire \thechain[1].chain8.inv_chain[187] ;
 wire \thechain[1].chain8.inv_chain[188] ;
 wire \thechain[1].chain8.inv_chain[189] ;
 wire \thechain[1].chain8.inv_chain[18] ;
 wire \thechain[1].chain8.inv_chain[190] ;
 wire \thechain[1].chain8.inv_chain[191] ;
 wire \thechain[1].chain8.inv_chain[192] ;
 wire \thechain[1].chain8.inv_chain[19] ;
 wire \thechain[1].chain8.inv_chain[1] ;
 wire \thechain[1].chain8.inv_chain[20] ;
 wire \thechain[1].chain8.inv_chain[21] ;
 wire \thechain[1].chain8.inv_chain[22] ;
 wire \thechain[1].chain8.inv_chain[23] ;
 wire \thechain[1].chain8.inv_chain[24] ;
 wire \thechain[1].chain8.inv_chain[25] ;
 wire \thechain[1].chain8.inv_chain[26] ;
 wire \thechain[1].chain8.inv_chain[27] ;
 wire \thechain[1].chain8.inv_chain[28] ;
 wire \thechain[1].chain8.inv_chain[29] ;
 wire \thechain[1].chain8.inv_chain[2] ;
 wire \thechain[1].chain8.inv_chain[30] ;
 wire \thechain[1].chain8.inv_chain[31] ;
 wire \thechain[1].chain8.inv_chain[32] ;
 wire \thechain[1].chain8.inv_chain[33] ;
 wire \thechain[1].chain8.inv_chain[34] ;
 wire \thechain[1].chain8.inv_chain[35] ;
 wire \thechain[1].chain8.inv_chain[36] ;
 wire \thechain[1].chain8.inv_chain[37] ;
 wire \thechain[1].chain8.inv_chain[38] ;
 wire \thechain[1].chain8.inv_chain[39] ;
 wire \thechain[1].chain8.inv_chain[3] ;
 wire \thechain[1].chain8.inv_chain[40] ;
 wire \thechain[1].chain8.inv_chain[41] ;
 wire \thechain[1].chain8.inv_chain[42] ;
 wire \thechain[1].chain8.inv_chain[43] ;
 wire \thechain[1].chain8.inv_chain[44] ;
 wire \thechain[1].chain8.inv_chain[45] ;
 wire \thechain[1].chain8.inv_chain[46] ;
 wire \thechain[1].chain8.inv_chain[47] ;
 wire \thechain[1].chain8.inv_chain[48] ;
 wire \thechain[1].chain8.inv_chain[49] ;
 wire \thechain[1].chain8.inv_chain[4] ;
 wire \thechain[1].chain8.inv_chain[50] ;
 wire \thechain[1].chain8.inv_chain[51] ;
 wire \thechain[1].chain8.inv_chain[52] ;
 wire \thechain[1].chain8.inv_chain[53] ;
 wire \thechain[1].chain8.inv_chain[54] ;
 wire \thechain[1].chain8.inv_chain[55] ;
 wire \thechain[1].chain8.inv_chain[56] ;
 wire \thechain[1].chain8.inv_chain[57] ;
 wire \thechain[1].chain8.inv_chain[58] ;
 wire \thechain[1].chain8.inv_chain[59] ;
 wire \thechain[1].chain8.inv_chain[5] ;
 wire \thechain[1].chain8.inv_chain[60] ;
 wire \thechain[1].chain8.inv_chain[61] ;
 wire \thechain[1].chain8.inv_chain[62] ;
 wire \thechain[1].chain8.inv_chain[63] ;
 wire \thechain[1].chain8.inv_chain[64] ;
 wire \thechain[1].chain8.inv_chain[65] ;
 wire \thechain[1].chain8.inv_chain[66] ;
 wire \thechain[1].chain8.inv_chain[67] ;
 wire \thechain[1].chain8.inv_chain[68] ;
 wire \thechain[1].chain8.inv_chain[69] ;
 wire \thechain[1].chain8.inv_chain[6] ;
 wire \thechain[1].chain8.inv_chain[70] ;
 wire \thechain[1].chain8.inv_chain[71] ;
 wire \thechain[1].chain8.inv_chain[72] ;
 wire \thechain[1].chain8.inv_chain[73] ;
 wire \thechain[1].chain8.inv_chain[74] ;
 wire \thechain[1].chain8.inv_chain[75] ;
 wire \thechain[1].chain8.inv_chain[76] ;
 wire \thechain[1].chain8.inv_chain[77] ;
 wire \thechain[1].chain8.inv_chain[78] ;
 wire \thechain[1].chain8.inv_chain[79] ;
 wire \thechain[1].chain8.inv_chain[7] ;
 wire \thechain[1].chain8.inv_chain[80] ;
 wire \thechain[1].chain8.inv_chain[81] ;
 wire \thechain[1].chain8.inv_chain[82] ;
 wire \thechain[1].chain8.inv_chain[83] ;
 wire \thechain[1].chain8.inv_chain[84] ;
 wire \thechain[1].chain8.inv_chain[85] ;
 wire \thechain[1].chain8.inv_chain[86] ;
 wire \thechain[1].chain8.inv_chain[87] ;
 wire \thechain[1].chain8.inv_chain[88] ;
 wire \thechain[1].chain8.inv_chain[89] ;
 wire \thechain[1].chain8.inv_chain[8] ;
 wire \thechain[1].chain8.inv_chain[90] ;
 wire \thechain[1].chain8.inv_chain[91] ;
 wire \thechain[1].chain8.inv_chain[92] ;
 wire \thechain[1].chain8.inv_chain[93] ;
 wire \thechain[1].chain8.inv_chain[94] ;
 wire \thechain[1].chain8.inv_chain[95] ;
 wire \thechain[1].chain8.inv_chain[96] ;
 wire \thechain[1].chain8.inv_chain[97] ;
 wire \thechain[1].chain8.inv_chain[98] ;
 wire \thechain[1].chain8.inv_chain[99] ;
 wire \thechain[1].chain8.inv_chain[9] ;
 wire \thechain[1].chain9.dout ;
 wire \thechain[1].chain9.inv_chain[0] ;
 wire \thechain[1].chain9.inv_chain[100] ;
 wire \thechain[1].chain9.inv_chain[101] ;
 wire \thechain[1].chain9.inv_chain[102] ;
 wire \thechain[1].chain9.inv_chain[103] ;
 wire \thechain[1].chain9.inv_chain[104] ;
 wire \thechain[1].chain9.inv_chain[105] ;
 wire \thechain[1].chain9.inv_chain[106] ;
 wire \thechain[1].chain9.inv_chain[107] ;
 wire \thechain[1].chain9.inv_chain[108] ;
 wire \thechain[1].chain9.inv_chain[109] ;
 wire \thechain[1].chain9.inv_chain[10] ;
 wire \thechain[1].chain9.inv_chain[110] ;
 wire \thechain[1].chain9.inv_chain[111] ;
 wire \thechain[1].chain9.inv_chain[112] ;
 wire \thechain[1].chain9.inv_chain[113] ;
 wire \thechain[1].chain9.inv_chain[114] ;
 wire \thechain[1].chain9.inv_chain[115] ;
 wire \thechain[1].chain9.inv_chain[116] ;
 wire \thechain[1].chain9.inv_chain[117] ;
 wire \thechain[1].chain9.inv_chain[118] ;
 wire \thechain[1].chain9.inv_chain[119] ;
 wire \thechain[1].chain9.inv_chain[11] ;
 wire \thechain[1].chain9.inv_chain[120] ;
 wire \thechain[1].chain9.inv_chain[121] ;
 wire \thechain[1].chain9.inv_chain[122] ;
 wire \thechain[1].chain9.inv_chain[123] ;
 wire \thechain[1].chain9.inv_chain[124] ;
 wire \thechain[1].chain9.inv_chain[125] ;
 wire \thechain[1].chain9.inv_chain[126] ;
 wire \thechain[1].chain9.inv_chain[127] ;
 wire \thechain[1].chain9.inv_chain[128] ;
 wire \thechain[1].chain9.inv_chain[129] ;
 wire \thechain[1].chain9.inv_chain[12] ;
 wire \thechain[1].chain9.inv_chain[130] ;
 wire \thechain[1].chain9.inv_chain[131] ;
 wire \thechain[1].chain9.inv_chain[132] ;
 wire \thechain[1].chain9.inv_chain[133] ;
 wire \thechain[1].chain9.inv_chain[134] ;
 wire \thechain[1].chain9.inv_chain[135] ;
 wire \thechain[1].chain9.inv_chain[136] ;
 wire \thechain[1].chain9.inv_chain[137] ;
 wire \thechain[1].chain9.inv_chain[138] ;
 wire \thechain[1].chain9.inv_chain[139] ;
 wire \thechain[1].chain9.inv_chain[13] ;
 wire \thechain[1].chain9.inv_chain[140] ;
 wire \thechain[1].chain9.inv_chain[141] ;
 wire \thechain[1].chain9.inv_chain[142] ;
 wire \thechain[1].chain9.inv_chain[143] ;
 wire \thechain[1].chain9.inv_chain[144] ;
 wire \thechain[1].chain9.inv_chain[145] ;
 wire \thechain[1].chain9.inv_chain[146] ;
 wire \thechain[1].chain9.inv_chain[147] ;
 wire \thechain[1].chain9.inv_chain[148] ;
 wire \thechain[1].chain9.inv_chain[149] ;
 wire \thechain[1].chain9.inv_chain[14] ;
 wire \thechain[1].chain9.inv_chain[150] ;
 wire \thechain[1].chain9.inv_chain[151] ;
 wire \thechain[1].chain9.inv_chain[152] ;
 wire \thechain[1].chain9.inv_chain[153] ;
 wire \thechain[1].chain9.inv_chain[154] ;
 wire \thechain[1].chain9.inv_chain[155] ;
 wire \thechain[1].chain9.inv_chain[156] ;
 wire \thechain[1].chain9.inv_chain[157] ;
 wire \thechain[1].chain9.inv_chain[158] ;
 wire \thechain[1].chain9.inv_chain[159] ;
 wire \thechain[1].chain9.inv_chain[15] ;
 wire \thechain[1].chain9.inv_chain[160] ;
 wire \thechain[1].chain9.inv_chain[161] ;
 wire \thechain[1].chain9.inv_chain[162] ;
 wire \thechain[1].chain9.inv_chain[163] ;
 wire \thechain[1].chain9.inv_chain[164] ;
 wire \thechain[1].chain9.inv_chain[165] ;
 wire \thechain[1].chain9.inv_chain[166] ;
 wire \thechain[1].chain9.inv_chain[167] ;
 wire \thechain[1].chain9.inv_chain[168] ;
 wire \thechain[1].chain9.inv_chain[169] ;
 wire \thechain[1].chain9.inv_chain[16] ;
 wire \thechain[1].chain9.inv_chain[170] ;
 wire \thechain[1].chain9.inv_chain[171] ;
 wire \thechain[1].chain9.inv_chain[172] ;
 wire \thechain[1].chain9.inv_chain[173] ;
 wire \thechain[1].chain9.inv_chain[174] ;
 wire \thechain[1].chain9.inv_chain[175] ;
 wire \thechain[1].chain9.inv_chain[176] ;
 wire \thechain[1].chain9.inv_chain[177] ;
 wire \thechain[1].chain9.inv_chain[178] ;
 wire \thechain[1].chain9.inv_chain[179] ;
 wire \thechain[1].chain9.inv_chain[17] ;
 wire \thechain[1].chain9.inv_chain[180] ;
 wire \thechain[1].chain9.inv_chain[181] ;
 wire \thechain[1].chain9.inv_chain[182] ;
 wire \thechain[1].chain9.inv_chain[183] ;
 wire \thechain[1].chain9.inv_chain[184] ;
 wire \thechain[1].chain9.inv_chain[185] ;
 wire \thechain[1].chain9.inv_chain[186] ;
 wire \thechain[1].chain9.inv_chain[187] ;
 wire \thechain[1].chain9.inv_chain[188] ;
 wire \thechain[1].chain9.inv_chain[189] ;
 wire \thechain[1].chain9.inv_chain[18] ;
 wire \thechain[1].chain9.inv_chain[190] ;
 wire \thechain[1].chain9.inv_chain[191] ;
 wire \thechain[1].chain9.inv_chain[192] ;
 wire \thechain[1].chain9.inv_chain[193] ;
 wire \thechain[1].chain9.inv_chain[194] ;
 wire \thechain[1].chain9.inv_chain[195] ;
 wire \thechain[1].chain9.inv_chain[196] ;
 wire \thechain[1].chain9.inv_chain[197] ;
 wire \thechain[1].chain9.inv_chain[198] ;
 wire \thechain[1].chain9.inv_chain[199] ;
 wire \thechain[1].chain9.inv_chain[19] ;
 wire \thechain[1].chain9.inv_chain[1] ;
 wire \thechain[1].chain9.inv_chain[200] ;
 wire \thechain[1].chain9.inv_chain[201] ;
 wire \thechain[1].chain9.inv_chain[202] ;
 wire \thechain[1].chain9.inv_chain[203] ;
 wire \thechain[1].chain9.inv_chain[204] ;
 wire \thechain[1].chain9.inv_chain[205] ;
 wire \thechain[1].chain9.inv_chain[206] ;
 wire \thechain[1].chain9.inv_chain[207] ;
 wire \thechain[1].chain9.inv_chain[208] ;
 wire \thechain[1].chain9.inv_chain[209] ;
 wire \thechain[1].chain9.inv_chain[20] ;
 wire \thechain[1].chain9.inv_chain[210] ;
 wire \thechain[1].chain9.inv_chain[211] ;
 wire \thechain[1].chain9.inv_chain[212] ;
 wire \thechain[1].chain9.inv_chain[213] ;
 wire \thechain[1].chain9.inv_chain[214] ;
 wire \thechain[1].chain9.inv_chain[215] ;
 wire \thechain[1].chain9.inv_chain[216] ;
 wire \thechain[1].chain9.inv_chain[217] ;
 wire \thechain[1].chain9.inv_chain[218] ;
 wire \thechain[1].chain9.inv_chain[219] ;
 wire \thechain[1].chain9.inv_chain[21] ;
 wire \thechain[1].chain9.inv_chain[220] ;
 wire \thechain[1].chain9.inv_chain[221] ;
 wire \thechain[1].chain9.inv_chain[222] ;
 wire \thechain[1].chain9.inv_chain[223] ;
 wire \thechain[1].chain9.inv_chain[224] ;
 wire \thechain[1].chain9.inv_chain[225] ;
 wire \thechain[1].chain9.inv_chain[226] ;
 wire \thechain[1].chain9.inv_chain[227] ;
 wire \thechain[1].chain9.inv_chain[228] ;
 wire \thechain[1].chain9.inv_chain[229] ;
 wire \thechain[1].chain9.inv_chain[22] ;
 wire \thechain[1].chain9.inv_chain[230] ;
 wire \thechain[1].chain9.inv_chain[231] ;
 wire \thechain[1].chain9.inv_chain[232] ;
 wire \thechain[1].chain9.inv_chain[233] ;
 wire \thechain[1].chain9.inv_chain[234] ;
 wire \thechain[1].chain9.inv_chain[235] ;
 wire \thechain[1].chain9.inv_chain[236] ;
 wire \thechain[1].chain9.inv_chain[237] ;
 wire \thechain[1].chain9.inv_chain[238] ;
 wire \thechain[1].chain9.inv_chain[239] ;
 wire \thechain[1].chain9.inv_chain[23] ;
 wire \thechain[1].chain9.inv_chain[240] ;
 wire \thechain[1].chain9.inv_chain[241] ;
 wire \thechain[1].chain9.inv_chain[242] ;
 wire \thechain[1].chain9.inv_chain[243] ;
 wire \thechain[1].chain9.inv_chain[244] ;
 wire \thechain[1].chain9.inv_chain[245] ;
 wire \thechain[1].chain9.inv_chain[246] ;
 wire \thechain[1].chain9.inv_chain[247] ;
 wire \thechain[1].chain9.inv_chain[248] ;
 wire \thechain[1].chain9.inv_chain[249] ;
 wire \thechain[1].chain9.inv_chain[24] ;
 wire \thechain[1].chain9.inv_chain[250] ;
 wire \thechain[1].chain9.inv_chain[251] ;
 wire \thechain[1].chain9.inv_chain[252] ;
 wire \thechain[1].chain9.inv_chain[253] ;
 wire \thechain[1].chain9.inv_chain[254] ;
 wire \thechain[1].chain9.inv_chain[255] ;
 wire \thechain[1].chain9.inv_chain[256] ;
 wire \thechain[1].chain9.inv_chain[25] ;
 wire \thechain[1].chain9.inv_chain[26] ;
 wire \thechain[1].chain9.inv_chain[27] ;
 wire \thechain[1].chain9.inv_chain[28] ;
 wire \thechain[1].chain9.inv_chain[29] ;
 wire \thechain[1].chain9.inv_chain[2] ;
 wire \thechain[1].chain9.inv_chain[30] ;
 wire \thechain[1].chain9.inv_chain[31] ;
 wire \thechain[1].chain9.inv_chain[32] ;
 wire \thechain[1].chain9.inv_chain[33] ;
 wire \thechain[1].chain9.inv_chain[34] ;
 wire \thechain[1].chain9.inv_chain[35] ;
 wire \thechain[1].chain9.inv_chain[36] ;
 wire \thechain[1].chain9.inv_chain[37] ;
 wire \thechain[1].chain9.inv_chain[38] ;
 wire \thechain[1].chain9.inv_chain[39] ;
 wire \thechain[1].chain9.inv_chain[3] ;
 wire \thechain[1].chain9.inv_chain[40] ;
 wire \thechain[1].chain9.inv_chain[41] ;
 wire \thechain[1].chain9.inv_chain[42] ;
 wire \thechain[1].chain9.inv_chain[43] ;
 wire \thechain[1].chain9.inv_chain[44] ;
 wire \thechain[1].chain9.inv_chain[45] ;
 wire \thechain[1].chain9.inv_chain[46] ;
 wire \thechain[1].chain9.inv_chain[47] ;
 wire \thechain[1].chain9.inv_chain[48] ;
 wire \thechain[1].chain9.inv_chain[49] ;
 wire \thechain[1].chain9.inv_chain[4] ;
 wire \thechain[1].chain9.inv_chain[50] ;
 wire \thechain[1].chain9.inv_chain[51] ;
 wire \thechain[1].chain9.inv_chain[52] ;
 wire \thechain[1].chain9.inv_chain[53] ;
 wire \thechain[1].chain9.inv_chain[54] ;
 wire \thechain[1].chain9.inv_chain[55] ;
 wire \thechain[1].chain9.inv_chain[56] ;
 wire \thechain[1].chain9.inv_chain[57] ;
 wire \thechain[1].chain9.inv_chain[58] ;
 wire \thechain[1].chain9.inv_chain[59] ;
 wire \thechain[1].chain9.inv_chain[5] ;
 wire \thechain[1].chain9.inv_chain[60] ;
 wire \thechain[1].chain9.inv_chain[61] ;
 wire \thechain[1].chain9.inv_chain[62] ;
 wire \thechain[1].chain9.inv_chain[63] ;
 wire \thechain[1].chain9.inv_chain[64] ;
 wire \thechain[1].chain9.inv_chain[65] ;
 wire \thechain[1].chain9.inv_chain[66] ;
 wire \thechain[1].chain9.inv_chain[67] ;
 wire \thechain[1].chain9.inv_chain[68] ;
 wire \thechain[1].chain9.inv_chain[69] ;
 wire \thechain[1].chain9.inv_chain[6] ;
 wire \thechain[1].chain9.inv_chain[70] ;
 wire \thechain[1].chain9.inv_chain[71] ;
 wire \thechain[1].chain9.inv_chain[72] ;
 wire \thechain[1].chain9.inv_chain[73] ;
 wire \thechain[1].chain9.inv_chain[74] ;
 wire \thechain[1].chain9.inv_chain[75] ;
 wire \thechain[1].chain9.inv_chain[76] ;
 wire \thechain[1].chain9.inv_chain[77] ;
 wire \thechain[1].chain9.inv_chain[78] ;
 wire \thechain[1].chain9.inv_chain[79] ;
 wire \thechain[1].chain9.inv_chain[7] ;
 wire \thechain[1].chain9.inv_chain[80] ;
 wire \thechain[1].chain9.inv_chain[81] ;
 wire \thechain[1].chain9.inv_chain[82] ;
 wire \thechain[1].chain9.inv_chain[83] ;
 wire \thechain[1].chain9.inv_chain[84] ;
 wire \thechain[1].chain9.inv_chain[85] ;
 wire \thechain[1].chain9.inv_chain[86] ;
 wire \thechain[1].chain9.inv_chain[87] ;
 wire \thechain[1].chain9.inv_chain[88] ;
 wire \thechain[1].chain9.inv_chain[89] ;
 wire \thechain[1].chain9.inv_chain[8] ;
 wire \thechain[1].chain9.inv_chain[90] ;
 wire \thechain[1].chain9.inv_chain[91] ;
 wire \thechain[1].chain9.inv_chain[92] ;
 wire \thechain[1].chain9.inv_chain[93] ;
 wire \thechain[1].chain9.inv_chain[94] ;
 wire \thechain[1].chain9.inv_chain[95] ;
 wire \thechain[1].chain9.inv_chain[96] ;
 wire \thechain[1].chain9.inv_chain[97] ;
 wire \thechain[1].chain9.inv_chain[98] ;
 wire \thechain[1].chain9.inv_chain[99] ;
 wire \thechain[1].chain9.inv_chain[9] ;
 wire \thechain[2].chain1.dout ;
 wire \thechain[2].chain1.inv_chain[0] ;
 wire \thechain[2].chain1.inv_chain[1] ;
 wire \thechain[2].chain1.inv_chain[2] ;
 wire \thechain[2].chain2.dout ;
 wire \thechain[2].chain2.inv_chain[0] ;
 wire \thechain[2].chain2.inv_chain[1] ;
 wire \thechain[2].chain2.inv_chain[2] ;
 wire \thechain[2].chain2.inv_chain[3] ;
 wire \thechain[2].chain2.inv_chain[4] ;
 wire \thechain[2].chain3.dout ;
 wire \thechain[2].chain3.inv_chain[0] ;
 wire \thechain[2].chain3.inv_chain[1] ;
 wire \thechain[2].chain3.inv_chain[2] ;
 wire \thechain[2].chain3.inv_chain[3] ;
 wire \thechain[2].chain3.inv_chain[4] ;
 wire \thechain[2].chain3.inv_chain[5] ;
 wire \thechain[2].chain3.inv_chain[6] ;
 wire \thechain[2].chain3.inv_chain[7] ;
 wire \thechain[2].chain3.inv_chain[8] ;
 wire \thechain[2].chain4.dout ;
 wire \thechain[2].chain4.inv_chain[0] ;
 wire \thechain[2].chain4.inv_chain[10] ;
 wire \thechain[2].chain4.inv_chain[11] ;
 wire \thechain[2].chain4.inv_chain[12] ;
 wire \thechain[2].chain4.inv_chain[13] ;
 wire \thechain[2].chain4.inv_chain[14] ;
 wire \thechain[2].chain4.inv_chain[15] ;
 wire \thechain[2].chain4.inv_chain[16] ;
 wire \thechain[2].chain4.inv_chain[1] ;
 wire \thechain[2].chain4.inv_chain[2] ;
 wire \thechain[2].chain4.inv_chain[3] ;
 wire \thechain[2].chain4.inv_chain[4] ;
 wire \thechain[2].chain4.inv_chain[5] ;
 wire \thechain[2].chain4.inv_chain[6] ;
 wire \thechain[2].chain4.inv_chain[7] ;
 wire \thechain[2].chain4.inv_chain[8] ;
 wire \thechain[2].chain4.inv_chain[9] ;
 wire \thechain[2].chain5.dout ;
 wire \thechain[2].chain5.inv_chain[0] ;
 wire \thechain[2].chain5.inv_chain[10] ;
 wire \thechain[2].chain5.inv_chain[11] ;
 wire \thechain[2].chain5.inv_chain[12] ;
 wire \thechain[2].chain5.inv_chain[13] ;
 wire \thechain[2].chain5.inv_chain[14] ;
 wire \thechain[2].chain5.inv_chain[15] ;
 wire \thechain[2].chain5.inv_chain[16] ;
 wire \thechain[2].chain5.inv_chain[17] ;
 wire \thechain[2].chain5.inv_chain[18] ;
 wire \thechain[2].chain5.inv_chain[19] ;
 wire \thechain[2].chain5.inv_chain[1] ;
 wire \thechain[2].chain5.inv_chain[20] ;
 wire \thechain[2].chain5.inv_chain[21] ;
 wire \thechain[2].chain5.inv_chain[22] ;
 wire \thechain[2].chain5.inv_chain[23] ;
 wire \thechain[2].chain5.inv_chain[24] ;
 wire \thechain[2].chain5.inv_chain[25] ;
 wire \thechain[2].chain5.inv_chain[26] ;
 wire \thechain[2].chain5.inv_chain[27] ;
 wire \thechain[2].chain5.inv_chain[28] ;
 wire \thechain[2].chain5.inv_chain[29] ;
 wire \thechain[2].chain5.inv_chain[2] ;
 wire \thechain[2].chain5.inv_chain[30] ;
 wire \thechain[2].chain5.inv_chain[31] ;
 wire \thechain[2].chain5.inv_chain[32] ;
 wire \thechain[2].chain5.inv_chain[3] ;
 wire \thechain[2].chain5.inv_chain[4] ;
 wire \thechain[2].chain5.inv_chain[5] ;
 wire \thechain[2].chain5.inv_chain[6] ;
 wire \thechain[2].chain5.inv_chain[7] ;
 wire \thechain[2].chain5.inv_chain[8] ;
 wire \thechain[2].chain5.inv_chain[9] ;
 wire \thechain[2].chain6.dout ;
 wire \thechain[2].chain6.inv_chain[0] ;
 wire \thechain[2].chain6.inv_chain[10] ;
 wire \thechain[2].chain6.inv_chain[11] ;
 wire \thechain[2].chain6.inv_chain[12] ;
 wire \thechain[2].chain6.inv_chain[13] ;
 wire \thechain[2].chain6.inv_chain[14] ;
 wire \thechain[2].chain6.inv_chain[15] ;
 wire \thechain[2].chain6.inv_chain[16] ;
 wire \thechain[2].chain6.inv_chain[17] ;
 wire \thechain[2].chain6.inv_chain[18] ;
 wire \thechain[2].chain6.inv_chain[19] ;
 wire \thechain[2].chain6.inv_chain[1] ;
 wire \thechain[2].chain6.inv_chain[20] ;
 wire \thechain[2].chain6.inv_chain[21] ;
 wire \thechain[2].chain6.inv_chain[22] ;
 wire \thechain[2].chain6.inv_chain[23] ;
 wire \thechain[2].chain6.inv_chain[24] ;
 wire \thechain[2].chain6.inv_chain[25] ;
 wire \thechain[2].chain6.inv_chain[26] ;
 wire \thechain[2].chain6.inv_chain[27] ;
 wire \thechain[2].chain6.inv_chain[28] ;
 wire \thechain[2].chain6.inv_chain[29] ;
 wire \thechain[2].chain6.inv_chain[2] ;
 wire \thechain[2].chain6.inv_chain[30] ;
 wire \thechain[2].chain6.inv_chain[31] ;
 wire \thechain[2].chain6.inv_chain[32] ;
 wire \thechain[2].chain6.inv_chain[33] ;
 wire \thechain[2].chain6.inv_chain[34] ;
 wire \thechain[2].chain6.inv_chain[35] ;
 wire \thechain[2].chain6.inv_chain[36] ;
 wire \thechain[2].chain6.inv_chain[37] ;
 wire \thechain[2].chain6.inv_chain[38] ;
 wire \thechain[2].chain6.inv_chain[39] ;
 wire \thechain[2].chain6.inv_chain[3] ;
 wire \thechain[2].chain6.inv_chain[40] ;
 wire \thechain[2].chain6.inv_chain[41] ;
 wire \thechain[2].chain6.inv_chain[42] ;
 wire \thechain[2].chain6.inv_chain[43] ;
 wire \thechain[2].chain6.inv_chain[44] ;
 wire \thechain[2].chain6.inv_chain[45] ;
 wire \thechain[2].chain6.inv_chain[46] ;
 wire \thechain[2].chain6.inv_chain[47] ;
 wire \thechain[2].chain6.inv_chain[48] ;
 wire \thechain[2].chain6.inv_chain[49] ;
 wire \thechain[2].chain6.inv_chain[4] ;
 wire \thechain[2].chain6.inv_chain[50] ;
 wire \thechain[2].chain6.inv_chain[51] ;
 wire \thechain[2].chain6.inv_chain[52] ;
 wire \thechain[2].chain6.inv_chain[53] ;
 wire \thechain[2].chain6.inv_chain[54] ;
 wire \thechain[2].chain6.inv_chain[55] ;
 wire \thechain[2].chain6.inv_chain[56] ;
 wire \thechain[2].chain6.inv_chain[57] ;
 wire \thechain[2].chain6.inv_chain[58] ;
 wire \thechain[2].chain6.inv_chain[59] ;
 wire \thechain[2].chain6.inv_chain[5] ;
 wire \thechain[2].chain6.inv_chain[60] ;
 wire \thechain[2].chain6.inv_chain[61] ;
 wire \thechain[2].chain6.inv_chain[62] ;
 wire \thechain[2].chain6.inv_chain[63] ;
 wire \thechain[2].chain6.inv_chain[64] ;
 wire \thechain[2].chain6.inv_chain[6] ;
 wire \thechain[2].chain6.inv_chain[7] ;
 wire \thechain[2].chain6.inv_chain[8] ;
 wire \thechain[2].chain6.inv_chain[9] ;
 wire \thechain[2].chain7.dout ;
 wire \thechain[2].chain7.inv_chain[0] ;
 wire \thechain[2].chain7.inv_chain[100] ;
 wire \thechain[2].chain7.inv_chain[101] ;
 wire \thechain[2].chain7.inv_chain[102] ;
 wire \thechain[2].chain7.inv_chain[103] ;
 wire \thechain[2].chain7.inv_chain[104] ;
 wire \thechain[2].chain7.inv_chain[105] ;
 wire \thechain[2].chain7.inv_chain[106] ;
 wire \thechain[2].chain7.inv_chain[107] ;
 wire \thechain[2].chain7.inv_chain[108] ;
 wire \thechain[2].chain7.inv_chain[109] ;
 wire \thechain[2].chain7.inv_chain[10] ;
 wire \thechain[2].chain7.inv_chain[110] ;
 wire \thechain[2].chain7.inv_chain[111] ;
 wire \thechain[2].chain7.inv_chain[112] ;
 wire \thechain[2].chain7.inv_chain[113] ;
 wire \thechain[2].chain7.inv_chain[114] ;
 wire \thechain[2].chain7.inv_chain[115] ;
 wire \thechain[2].chain7.inv_chain[116] ;
 wire \thechain[2].chain7.inv_chain[117] ;
 wire \thechain[2].chain7.inv_chain[118] ;
 wire \thechain[2].chain7.inv_chain[119] ;
 wire \thechain[2].chain7.inv_chain[11] ;
 wire \thechain[2].chain7.inv_chain[120] ;
 wire \thechain[2].chain7.inv_chain[121] ;
 wire \thechain[2].chain7.inv_chain[122] ;
 wire \thechain[2].chain7.inv_chain[123] ;
 wire \thechain[2].chain7.inv_chain[124] ;
 wire \thechain[2].chain7.inv_chain[125] ;
 wire \thechain[2].chain7.inv_chain[126] ;
 wire \thechain[2].chain7.inv_chain[127] ;
 wire \thechain[2].chain7.inv_chain[128] ;
 wire \thechain[2].chain7.inv_chain[12] ;
 wire \thechain[2].chain7.inv_chain[13] ;
 wire \thechain[2].chain7.inv_chain[14] ;
 wire \thechain[2].chain7.inv_chain[15] ;
 wire \thechain[2].chain7.inv_chain[16] ;
 wire \thechain[2].chain7.inv_chain[17] ;
 wire \thechain[2].chain7.inv_chain[18] ;
 wire \thechain[2].chain7.inv_chain[19] ;
 wire \thechain[2].chain7.inv_chain[1] ;
 wire \thechain[2].chain7.inv_chain[20] ;
 wire \thechain[2].chain7.inv_chain[21] ;
 wire \thechain[2].chain7.inv_chain[22] ;
 wire \thechain[2].chain7.inv_chain[23] ;
 wire \thechain[2].chain7.inv_chain[24] ;
 wire \thechain[2].chain7.inv_chain[25] ;
 wire \thechain[2].chain7.inv_chain[26] ;
 wire \thechain[2].chain7.inv_chain[27] ;
 wire \thechain[2].chain7.inv_chain[28] ;
 wire \thechain[2].chain7.inv_chain[29] ;
 wire \thechain[2].chain7.inv_chain[2] ;
 wire \thechain[2].chain7.inv_chain[30] ;
 wire \thechain[2].chain7.inv_chain[31] ;
 wire \thechain[2].chain7.inv_chain[32] ;
 wire \thechain[2].chain7.inv_chain[33] ;
 wire \thechain[2].chain7.inv_chain[34] ;
 wire \thechain[2].chain7.inv_chain[35] ;
 wire \thechain[2].chain7.inv_chain[36] ;
 wire \thechain[2].chain7.inv_chain[37] ;
 wire \thechain[2].chain7.inv_chain[38] ;
 wire \thechain[2].chain7.inv_chain[39] ;
 wire \thechain[2].chain7.inv_chain[3] ;
 wire \thechain[2].chain7.inv_chain[40] ;
 wire \thechain[2].chain7.inv_chain[41] ;
 wire \thechain[2].chain7.inv_chain[42] ;
 wire \thechain[2].chain7.inv_chain[43] ;
 wire \thechain[2].chain7.inv_chain[44] ;
 wire \thechain[2].chain7.inv_chain[45] ;
 wire \thechain[2].chain7.inv_chain[46] ;
 wire \thechain[2].chain7.inv_chain[47] ;
 wire \thechain[2].chain7.inv_chain[48] ;
 wire \thechain[2].chain7.inv_chain[49] ;
 wire \thechain[2].chain7.inv_chain[4] ;
 wire \thechain[2].chain7.inv_chain[50] ;
 wire \thechain[2].chain7.inv_chain[51] ;
 wire \thechain[2].chain7.inv_chain[52] ;
 wire \thechain[2].chain7.inv_chain[53] ;
 wire \thechain[2].chain7.inv_chain[54] ;
 wire \thechain[2].chain7.inv_chain[55] ;
 wire \thechain[2].chain7.inv_chain[56] ;
 wire \thechain[2].chain7.inv_chain[57] ;
 wire \thechain[2].chain7.inv_chain[58] ;
 wire \thechain[2].chain7.inv_chain[59] ;
 wire \thechain[2].chain7.inv_chain[5] ;
 wire \thechain[2].chain7.inv_chain[60] ;
 wire \thechain[2].chain7.inv_chain[61] ;
 wire \thechain[2].chain7.inv_chain[62] ;
 wire \thechain[2].chain7.inv_chain[63] ;
 wire \thechain[2].chain7.inv_chain[64] ;
 wire \thechain[2].chain7.inv_chain[65] ;
 wire \thechain[2].chain7.inv_chain[66] ;
 wire \thechain[2].chain7.inv_chain[67] ;
 wire \thechain[2].chain7.inv_chain[68] ;
 wire \thechain[2].chain7.inv_chain[69] ;
 wire \thechain[2].chain7.inv_chain[6] ;
 wire \thechain[2].chain7.inv_chain[70] ;
 wire \thechain[2].chain7.inv_chain[71] ;
 wire \thechain[2].chain7.inv_chain[72] ;
 wire \thechain[2].chain7.inv_chain[73] ;
 wire \thechain[2].chain7.inv_chain[74] ;
 wire \thechain[2].chain7.inv_chain[75] ;
 wire \thechain[2].chain7.inv_chain[76] ;
 wire \thechain[2].chain7.inv_chain[77] ;
 wire \thechain[2].chain7.inv_chain[78] ;
 wire \thechain[2].chain7.inv_chain[79] ;
 wire \thechain[2].chain7.inv_chain[7] ;
 wire \thechain[2].chain7.inv_chain[80] ;
 wire \thechain[2].chain7.inv_chain[81] ;
 wire \thechain[2].chain7.inv_chain[82] ;
 wire \thechain[2].chain7.inv_chain[83] ;
 wire \thechain[2].chain7.inv_chain[84] ;
 wire \thechain[2].chain7.inv_chain[85] ;
 wire \thechain[2].chain7.inv_chain[86] ;
 wire \thechain[2].chain7.inv_chain[87] ;
 wire \thechain[2].chain7.inv_chain[88] ;
 wire \thechain[2].chain7.inv_chain[89] ;
 wire \thechain[2].chain7.inv_chain[8] ;
 wire \thechain[2].chain7.inv_chain[90] ;
 wire \thechain[2].chain7.inv_chain[91] ;
 wire \thechain[2].chain7.inv_chain[92] ;
 wire \thechain[2].chain7.inv_chain[93] ;
 wire \thechain[2].chain7.inv_chain[94] ;
 wire \thechain[2].chain7.inv_chain[95] ;
 wire \thechain[2].chain7.inv_chain[96] ;
 wire \thechain[2].chain7.inv_chain[97] ;
 wire \thechain[2].chain7.inv_chain[98] ;
 wire \thechain[2].chain7.inv_chain[99] ;
 wire \thechain[2].chain7.inv_chain[9] ;
 wire \thechain[2].chain8.dout ;
 wire \thechain[2].chain8.inv_chain[0] ;
 wire \thechain[2].chain8.inv_chain[100] ;
 wire \thechain[2].chain8.inv_chain[101] ;
 wire \thechain[2].chain8.inv_chain[102] ;
 wire \thechain[2].chain8.inv_chain[103] ;
 wire \thechain[2].chain8.inv_chain[104] ;
 wire \thechain[2].chain8.inv_chain[105] ;
 wire \thechain[2].chain8.inv_chain[106] ;
 wire \thechain[2].chain8.inv_chain[107] ;
 wire \thechain[2].chain8.inv_chain[108] ;
 wire \thechain[2].chain8.inv_chain[109] ;
 wire \thechain[2].chain8.inv_chain[10] ;
 wire \thechain[2].chain8.inv_chain[110] ;
 wire \thechain[2].chain8.inv_chain[111] ;
 wire \thechain[2].chain8.inv_chain[112] ;
 wire \thechain[2].chain8.inv_chain[113] ;
 wire \thechain[2].chain8.inv_chain[114] ;
 wire \thechain[2].chain8.inv_chain[115] ;
 wire \thechain[2].chain8.inv_chain[116] ;
 wire \thechain[2].chain8.inv_chain[117] ;
 wire \thechain[2].chain8.inv_chain[118] ;
 wire \thechain[2].chain8.inv_chain[119] ;
 wire \thechain[2].chain8.inv_chain[11] ;
 wire \thechain[2].chain8.inv_chain[120] ;
 wire \thechain[2].chain8.inv_chain[121] ;
 wire \thechain[2].chain8.inv_chain[122] ;
 wire \thechain[2].chain8.inv_chain[123] ;
 wire \thechain[2].chain8.inv_chain[124] ;
 wire \thechain[2].chain8.inv_chain[125] ;
 wire \thechain[2].chain8.inv_chain[126] ;
 wire \thechain[2].chain8.inv_chain[127] ;
 wire \thechain[2].chain8.inv_chain[128] ;
 wire \thechain[2].chain8.inv_chain[129] ;
 wire \thechain[2].chain8.inv_chain[12] ;
 wire \thechain[2].chain8.inv_chain[130] ;
 wire \thechain[2].chain8.inv_chain[131] ;
 wire \thechain[2].chain8.inv_chain[132] ;
 wire \thechain[2].chain8.inv_chain[133] ;
 wire \thechain[2].chain8.inv_chain[134] ;
 wire \thechain[2].chain8.inv_chain[135] ;
 wire \thechain[2].chain8.inv_chain[136] ;
 wire \thechain[2].chain8.inv_chain[137] ;
 wire \thechain[2].chain8.inv_chain[138] ;
 wire \thechain[2].chain8.inv_chain[139] ;
 wire \thechain[2].chain8.inv_chain[13] ;
 wire \thechain[2].chain8.inv_chain[140] ;
 wire \thechain[2].chain8.inv_chain[141] ;
 wire \thechain[2].chain8.inv_chain[142] ;
 wire \thechain[2].chain8.inv_chain[143] ;
 wire \thechain[2].chain8.inv_chain[144] ;
 wire \thechain[2].chain8.inv_chain[145] ;
 wire \thechain[2].chain8.inv_chain[146] ;
 wire \thechain[2].chain8.inv_chain[147] ;
 wire \thechain[2].chain8.inv_chain[148] ;
 wire \thechain[2].chain8.inv_chain[149] ;
 wire \thechain[2].chain8.inv_chain[14] ;
 wire \thechain[2].chain8.inv_chain[150] ;
 wire \thechain[2].chain8.inv_chain[151] ;
 wire \thechain[2].chain8.inv_chain[152] ;
 wire \thechain[2].chain8.inv_chain[153] ;
 wire \thechain[2].chain8.inv_chain[154] ;
 wire \thechain[2].chain8.inv_chain[155] ;
 wire \thechain[2].chain8.inv_chain[156] ;
 wire \thechain[2].chain8.inv_chain[157] ;
 wire \thechain[2].chain8.inv_chain[158] ;
 wire \thechain[2].chain8.inv_chain[159] ;
 wire \thechain[2].chain8.inv_chain[15] ;
 wire \thechain[2].chain8.inv_chain[160] ;
 wire \thechain[2].chain8.inv_chain[161] ;
 wire \thechain[2].chain8.inv_chain[162] ;
 wire \thechain[2].chain8.inv_chain[163] ;
 wire \thechain[2].chain8.inv_chain[164] ;
 wire \thechain[2].chain8.inv_chain[165] ;
 wire \thechain[2].chain8.inv_chain[166] ;
 wire \thechain[2].chain8.inv_chain[167] ;
 wire \thechain[2].chain8.inv_chain[168] ;
 wire \thechain[2].chain8.inv_chain[169] ;
 wire \thechain[2].chain8.inv_chain[16] ;
 wire \thechain[2].chain8.inv_chain[170] ;
 wire \thechain[2].chain8.inv_chain[171] ;
 wire \thechain[2].chain8.inv_chain[172] ;
 wire \thechain[2].chain8.inv_chain[173] ;
 wire \thechain[2].chain8.inv_chain[174] ;
 wire \thechain[2].chain8.inv_chain[175] ;
 wire \thechain[2].chain8.inv_chain[176] ;
 wire \thechain[2].chain8.inv_chain[177] ;
 wire \thechain[2].chain8.inv_chain[178] ;
 wire \thechain[2].chain8.inv_chain[179] ;
 wire \thechain[2].chain8.inv_chain[17] ;
 wire \thechain[2].chain8.inv_chain[180] ;
 wire \thechain[2].chain8.inv_chain[181] ;
 wire \thechain[2].chain8.inv_chain[182] ;
 wire \thechain[2].chain8.inv_chain[183] ;
 wire \thechain[2].chain8.inv_chain[184] ;
 wire \thechain[2].chain8.inv_chain[185] ;
 wire \thechain[2].chain8.inv_chain[186] ;
 wire \thechain[2].chain8.inv_chain[187] ;
 wire \thechain[2].chain8.inv_chain[188] ;
 wire \thechain[2].chain8.inv_chain[189] ;
 wire \thechain[2].chain8.inv_chain[18] ;
 wire \thechain[2].chain8.inv_chain[190] ;
 wire \thechain[2].chain8.inv_chain[191] ;
 wire \thechain[2].chain8.inv_chain[192] ;
 wire \thechain[2].chain8.inv_chain[19] ;
 wire \thechain[2].chain8.inv_chain[1] ;
 wire \thechain[2].chain8.inv_chain[20] ;
 wire \thechain[2].chain8.inv_chain[21] ;
 wire \thechain[2].chain8.inv_chain[22] ;
 wire \thechain[2].chain8.inv_chain[23] ;
 wire \thechain[2].chain8.inv_chain[24] ;
 wire \thechain[2].chain8.inv_chain[25] ;
 wire \thechain[2].chain8.inv_chain[26] ;
 wire \thechain[2].chain8.inv_chain[27] ;
 wire \thechain[2].chain8.inv_chain[28] ;
 wire \thechain[2].chain8.inv_chain[29] ;
 wire \thechain[2].chain8.inv_chain[2] ;
 wire \thechain[2].chain8.inv_chain[30] ;
 wire \thechain[2].chain8.inv_chain[31] ;
 wire \thechain[2].chain8.inv_chain[32] ;
 wire \thechain[2].chain8.inv_chain[33] ;
 wire \thechain[2].chain8.inv_chain[34] ;
 wire \thechain[2].chain8.inv_chain[35] ;
 wire \thechain[2].chain8.inv_chain[36] ;
 wire \thechain[2].chain8.inv_chain[37] ;
 wire \thechain[2].chain8.inv_chain[38] ;
 wire \thechain[2].chain8.inv_chain[39] ;
 wire \thechain[2].chain8.inv_chain[3] ;
 wire \thechain[2].chain8.inv_chain[40] ;
 wire \thechain[2].chain8.inv_chain[41] ;
 wire \thechain[2].chain8.inv_chain[42] ;
 wire \thechain[2].chain8.inv_chain[43] ;
 wire \thechain[2].chain8.inv_chain[44] ;
 wire \thechain[2].chain8.inv_chain[45] ;
 wire \thechain[2].chain8.inv_chain[46] ;
 wire \thechain[2].chain8.inv_chain[47] ;
 wire \thechain[2].chain8.inv_chain[48] ;
 wire \thechain[2].chain8.inv_chain[49] ;
 wire \thechain[2].chain8.inv_chain[4] ;
 wire \thechain[2].chain8.inv_chain[50] ;
 wire \thechain[2].chain8.inv_chain[51] ;
 wire \thechain[2].chain8.inv_chain[52] ;
 wire \thechain[2].chain8.inv_chain[53] ;
 wire \thechain[2].chain8.inv_chain[54] ;
 wire \thechain[2].chain8.inv_chain[55] ;
 wire \thechain[2].chain8.inv_chain[56] ;
 wire \thechain[2].chain8.inv_chain[57] ;
 wire \thechain[2].chain8.inv_chain[58] ;
 wire \thechain[2].chain8.inv_chain[59] ;
 wire \thechain[2].chain8.inv_chain[5] ;
 wire \thechain[2].chain8.inv_chain[60] ;
 wire \thechain[2].chain8.inv_chain[61] ;
 wire \thechain[2].chain8.inv_chain[62] ;
 wire \thechain[2].chain8.inv_chain[63] ;
 wire \thechain[2].chain8.inv_chain[64] ;
 wire \thechain[2].chain8.inv_chain[65] ;
 wire \thechain[2].chain8.inv_chain[66] ;
 wire \thechain[2].chain8.inv_chain[67] ;
 wire \thechain[2].chain8.inv_chain[68] ;
 wire \thechain[2].chain8.inv_chain[69] ;
 wire \thechain[2].chain8.inv_chain[6] ;
 wire \thechain[2].chain8.inv_chain[70] ;
 wire \thechain[2].chain8.inv_chain[71] ;
 wire \thechain[2].chain8.inv_chain[72] ;
 wire \thechain[2].chain8.inv_chain[73] ;
 wire \thechain[2].chain8.inv_chain[74] ;
 wire \thechain[2].chain8.inv_chain[75] ;
 wire \thechain[2].chain8.inv_chain[76] ;
 wire \thechain[2].chain8.inv_chain[77] ;
 wire \thechain[2].chain8.inv_chain[78] ;
 wire \thechain[2].chain8.inv_chain[79] ;
 wire \thechain[2].chain8.inv_chain[7] ;
 wire \thechain[2].chain8.inv_chain[80] ;
 wire \thechain[2].chain8.inv_chain[81] ;
 wire \thechain[2].chain8.inv_chain[82] ;
 wire \thechain[2].chain8.inv_chain[83] ;
 wire \thechain[2].chain8.inv_chain[84] ;
 wire \thechain[2].chain8.inv_chain[85] ;
 wire \thechain[2].chain8.inv_chain[86] ;
 wire \thechain[2].chain8.inv_chain[87] ;
 wire \thechain[2].chain8.inv_chain[88] ;
 wire \thechain[2].chain8.inv_chain[89] ;
 wire \thechain[2].chain8.inv_chain[8] ;
 wire \thechain[2].chain8.inv_chain[90] ;
 wire \thechain[2].chain8.inv_chain[91] ;
 wire \thechain[2].chain8.inv_chain[92] ;
 wire \thechain[2].chain8.inv_chain[93] ;
 wire \thechain[2].chain8.inv_chain[94] ;
 wire \thechain[2].chain8.inv_chain[95] ;
 wire \thechain[2].chain8.inv_chain[96] ;
 wire \thechain[2].chain8.inv_chain[97] ;
 wire \thechain[2].chain8.inv_chain[98] ;
 wire \thechain[2].chain8.inv_chain[99] ;
 wire \thechain[2].chain8.inv_chain[9] ;
 wire \thechain[2].chain9.dout ;
 wire \thechain[2].chain9.inv_chain[0] ;
 wire \thechain[2].chain9.inv_chain[100] ;
 wire \thechain[2].chain9.inv_chain[101] ;
 wire \thechain[2].chain9.inv_chain[102] ;
 wire \thechain[2].chain9.inv_chain[103] ;
 wire \thechain[2].chain9.inv_chain[104] ;
 wire \thechain[2].chain9.inv_chain[105] ;
 wire \thechain[2].chain9.inv_chain[106] ;
 wire \thechain[2].chain9.inv_chain[107] ;
 wire \thechain[2].chain9.inv_chain[108] ;
 wire \thechain[2].chain9.inv_chain[109] ;
 wire \thechain[2].chain9.inv_chain[10] ;
 wire \thechain[2].chain9.inv_chain[110] ;
 wire \thechain[2].chain9.inv_chain[111] ;
 wire \thechain[2].chain9.inv_chain[112] ;
 wire \thechain[2].chain9.inv_chain[113] ;
 wire \thechain[2].chain9.inv_chain[114] ;
 wire \thechain[2].chain9.inv_chain[115] ;
 wire \thechain[2].chain9.inv_chain[116] ;
 wire \thechain[2].chain9.inv_chain[117] ;
 wire \thechain[2].chain9.inv_chain[118] ;
 wire \thechain[2].chain9.inv_chain[119] ;
 wire \thechain[2].chain9.inv_chain[11] ;
 wire \thechain[2].chain9.inv_chain[120] ;
 wire \thechain[2].chain9.inv_chain[121] ;
 wire \thechain[2].chain9.inv_chain[122] ;
 wire \thechain[2].chain9.inv_chain[123] ;
 wire \thechain[2].chain9.inv_chain[124] ;
 wire \thechain[2].chain9.inv_chain[125] ;
 wire \thechain[2].chain9.inv_chain[126] ;
 wire \thechain[2].chain9.inv_chain[127] ;
 wire \thechain[2].chain9.inv_chain[128] ;
 wire \thechain[2].chain9.inv_chain[129] ;
 wire \thechain[2].chain9.inv_chain[12] ;
 wire \thechain[2].chain9.inv_chain[130] ;
 wire \thechain[2].chain9.inv_chain[131] ;
 wire \thechain[2].chain9.inv_chain[132] ;
 wire \thechain[2].chain9.inv_chain[133] ;
 wire \thechain[2].chain9.inv_chain[134] ;
 wire \thechain[2].chain9.inv_chain[135] ;
 wire \thechain[2].chain9.inv_chain[136] ;
 wire \thechain[2].chain9.inv_chain[137] ;
 wire \thechain[2].chain9.inv_chain[138] ;
 wire \thechain[2].chain9.inv_chain[139] ;
 wire \thechain[2].chain9.inv_chain[13] ;
 wire \thechain[2].chain9.inv_chain[140] ;
 wire \thechain[2].chain9.inv_chain[141] ;
 wire \thechain[2].chain9.inv_chain[142] ;
 wire \thechain[2].chain9.inv_chain[143] ;
 wire \thechain[2].chain9.inv_chain[144] ;
 wire \thechain[2].chain9.inv_chain[145] ;
 wire \thechain[2].chain9.inv_chain[146] ;
 wire \thechain[2].chain9.inv_chain[147] ;
 wire \thechain[2].chain9.inv_chain[148] ;
 wire \thechain[2].chain9.inv_chain[149] ;
 wire \thechain[2].chain9.inv_chain[14] ;
 wire \thechain[2].chain9.inv_chain[150] ;
 wire \thechain[2].chain9.inv_chain[151] ;
 wire \thechain[2].chain9.inv_chain[152] ;
 wire \thechain[2].chain9.inv_chain[153] ;
 wire \thechain[2].chain9.inv_chain[154] ;
 wire \thechain[2].chain9.inv_chain[155] ;
 wire \thechain[2].chain9.inv_chain[156] ;
 wire \thechain[2].chain9.inv_chain[157] ;
 wire \thechain[2].chain9.inv_chain[158] ;
 wire \thechain[2].chain9.inv_chain[159] ;
 wire \thechain[2].chain9.inv_chain[15] ;
 wire \thechain[2].chain9.inv_chain[160] ;
 wire \thechain[2].chain9.inv_chain[161] ;
 wire \thechain[2].chain9.inv_chain[162] ;
 wire \thechain[2].chain9.inv_chain[163] ;
 wire \thechain[2].chain9.inv_chain[164] ;
 wire \thechain[2].chain9.inv_chain[165] ;
 wire \thechain[2].chain9.inv_chain[166] ;
 wire \thechain[2].chain9.inv_chain[167] ;
 wire \thechain[2].chain9.inv_chain[168] ;
 wire \thechain[2].chain9.inv_chain[169] ;
 wire \thechain[2].chain9.inv_chain[16] ;
 wire \thechain[2].chain9.inv_chain[170] ;
 wire \thechain[2].chain9.inv_chain[171] ;
 wire \thechain[2].chain9.inv_chain[172] ;
 wire \thechain[2].chain9.inv_chain[173] ;
 wire \thechain[2].chain9.inv_chain[174] ;
 wire \thechain[2].chain9.inv_chain[175] ;
 wire \thechain[2].chain9.inv_chain[176] ;
 wire \thechain[2].chain9.inv_chain[177] ;
 wire \thechain[2].chain9.inv_chain[178] ;
 wire \thechain[2].chain9.inv_chain[179] ;
 wire \thechain[2].chain9.inv_chain[17] ;
 wire \thechain[2].chain9.inv_chain[180] ;
 wire \thechain[2].chain9.inv_chain[181] ;
 wire \thechain[2].chain9.inv_chain[182] ;
 wire \thechain[2].chain9.inv_chain[183] ;
 wire \thechain[2].chain9.inv_chain[184] ;
 wire \thechain[2].chain9.inv_chain[185] ;
 wire \thechain[2].chain9.inv_chain[186] ;
 wire \thechain[2].chain9.inv_chain[187] ;
 wire \thechain[2].chain9.inv_chain[188] ;
 wire \thechain[2].chain9.inv_chain[189] ;
 wire \thechain[2].chain9.inv_chain[18] ;
 wire \thechain[2].chain9.inv_chain[190] ;
 wire \thechain[2].chain9.inv_chain[191] ;
 wire \thechain[2].chain9.inv_chain[192] ;
 wire \thechain[2].chain9.inv_chain[193] ;
 wire \thechain[2].chain9.inv_chain[194] ;
 wire \thechain[2].chain9.inv_chain[195] ;
 wire \thechain[2].chain9.inv_chain[196] ;
 wire \thechain[2].chain9.inv_chain[197] ;
 wire \thechain[2].chain9.inv_chain[198] ;
 wire \thechain[2].chain9.inv_chain[199] ;
 wire \thechain[2].chain9.inv_chain[19] ;
 wire \thechain[2].chain9.inv_chain[1] ;
 wire \thechain[2].chain9.inv_chain[200] ;
 wire \thechain[2].chain9.inv_chain[201] ;
 wire \thechain[2].chain9.inv_chain[202] ;
 wire \thechain[2].chain9.inv_chain[203] ;
 wire \thechain[2].chain9.inv_chain[204] ;
 wire \thechain[2].chain9.inv_chain[205] ;
 wire \thechain[2].chain9.inv_chain[206] ;
 wire \thechain[2].chain9.inv_chain[207] ;
 wire \thechain[2].chain9.inv_chain[208] ;
 wire \thechain[2].chain9.inv_chain[209] ;
 wire \thechain[2].chain9.inv_chain[20] ;
 wire \thechain[2].chain9.inv_chain[210] ;
 wire \thechain[2].chain9.inv_chain[211] ;
 wire \thechain[2].chain9.inv_chain[212] ;
 wire \thechain[2].chain9.inv_chain[213] ;
 wire \thechain[2].chain9.inv_chain[214] ;
 wire \thechain[2].chain9.inv_chain[215] ;
 wire \thechain[2].chain9.inv_chain[216] ;
 wire \thechain[2].chain9.inv_chain[217] ;
 wire \thechain[2].chain9.inv_chain[218] ;
 wire \thechain[2].chain9.inv_chain[219] ;
 wire \thechain[2].chain9.inv_chain[21] ;
 wire \thechain[2].chain9.inv_chain[220] ;
 wire \thechain[2].chain9.inv_chain[221] ;
 wire \thechain[2].chain9.inv_chain[222] ;
 wire \thechain[2].chain9.inv_chain[223] ;
 wire \thechain[2].chain9.inv_chain[224] ;
 wire \thechain[2].chain9.inv_chain[225] ;
 wire \thechain[2].chain9.inv_chain[226] ;
 wire \thechain[2].chain9.inv_chain[227] ;
 wire \thechain[2].chain9.inv_chain[228] ;
 wire \thechain[2].chain9.inv_chain[229] ;
 wire \thechain[2].chain9.inv_chain[22] ;
 wire \thechain[2].chain9.inv_chain[230] ;
 wire \thechain[2].chain9.inv_chain[231] ;
 wire \thechain[2].chain9.inv_chain[232] ;
 wire \thechain[2].chain9.inv_chain[233] ;
 wire \thechain[2].chain9.inv_chain[234] ;
 wire \thechain[2].chain9.inv_chain[235] ;
 wire \thechain[2].chain9.inv_chain[236] ;
 wire \thechain[2].chain9.inv_chain[237] ;
 wire \thechain[2].chain9.inv_chain[238] ;
 wire \thechain[2].chain9.inv_chain[239] ;
 wire \thechain[2].chain9.inv_chain[23] ;
 wire \thechain[2].chain9.inv_chain[240] ;
 wire \thechain[2].chain9.inv_chain[241] ;
 wire \thechain[2].chain9.inv_chain[242] ;
 wire \thechain[2].chain9.inv_chain[243] ;
 wire \thechain[2].chain9.inv_chain[244] ;
 wire \thechain[2].chain9.inv_chain[245] ;
 wire \thechain[2].chain9.inv_chain[246] ;
 wire \thechain[2].chain9.inv_chain[247] ;
 wire \thechain[2].chain9.inv_chain[248] ;
 wire \thechain[2].chain9.inv_chain[249] ;
 wire \thechain[2].chain9.inv_chain[24] ;
 wire \thechain[2].chain9.inv_chain[250] ;
 wire \thechain[2].chain9.inv_chain[251] ;
 wire \thechain[2].chain9.inv_chain[252] ;
 wire \thechain[2].chain9.inv_chain[253] ;
 wire \thechain[2].chain9.inv_chain[254] ;
 wire \thechain[2].chain9.inv_chain[255] ;
 wire \thechain[2].chain9.inv_chain[256] ;
 wire \thechain[2].chain9.inv_chain[25] ;
 wire \thechain[2].chain9.inv_chain[26] ;
 wire \thechain[2].chain9.inv_chain[27] ;
 wire \thechain[2].chain9.inv_chain[28] ;
 wire \thechain[2].chain9.inv_chain[29] ;
 wire \thechain[2].chain9.inv_chain[2] ;
 wire \thechain[2].chain9.inv_chain[30] ;
 wire \thechain[2].chain9.inv_chain[31] ;
 wire \thechain[2].chain9.inv_chain[32] ;
 wire \thechain[2].chain9.inv_chain[33] ;
 wire \thechain[2].chain9.inv_chain[34] ;
 wire \thechain[2].chain9.inv_chain[35] ;
 wire \thechain[2].chain9.inv_chain[36] ;
 wire \thechain[2].chain9.inv_chain[37] ;
 wire \thechain[2].chain9.inv_chain[38] ;
 wire \thechain[2].chain9.inv_chain[39] ;
 wire \thechain[2].chain9.inv_chain[3] ;
 wire \thechain[2].chain9.inv_chain[40] ;
 wire \thechain[2].chain9.inv_chain[41] ;
 wire \thechain[2].chain9.inv_chain[42] ;
 wire \thechain[2].chain9.inv_chain[43] ;
 wire \thechain[2].chain9.inv_chain[44] ;
 wire \thechain[2].chain9.inv_chain[45] ;
 wire \thechain[2].chain9.inv_chain[46] ;
 wire \thechain[2].chain9.inv_chain[47] ;
 wire \thechain[2].chain9.inv_chain[48] ;
 wire \thechain[2].chain9.inv_chain[49] ;
 wire \thechain[2].chain9.inv_chain[4] ;
 wire \thechain[2].chain9.inv_chain[50] ;
 wire \thechain[2].chain9.inv_chain[51] ;
 wire \thechain[2].chain9.inv_chain[52] ;
 wire \thechain[2].chain9.inv_chain[53] ;
 wire \thechain[2].chain9.inv_chain[54] ;
 wire \thechain[2].chain9.inv_chain[55] ;
 wire \thechain[2].chain9.inv_chain[56] ;
 wire \thechain[2].chain9.inv_chain[57] ;
 wire \thechain[2].chain9.inv_chain[58] ;
 wire \thechain[2].chain9.inv_chain[59] ;
 wire \thechain[2].chain9.inv_chain[5] ;
 wire \thechain[2].chain9.inv_chain[60] ;
 wire \thechain[2].chain9.inv_chain[61] ;
 wire \thechain[2].chain9.inv_chain[62] ;
 wire \thechain[2].chain9.inv_chain[63] ;
 wire \thechain[2].chain9.inv_chain[64] ;
 wire \thechain[2].chain9.inv_chain[65] ;
 wire \thechain[2].chain9.inv_chain[66] ;
 wire \thechain[2].chain9.inv_chain[67] ;
 wire \thechain[2].chain9.inv_chain[68] ;
 wire \thechain[2].chain9.inv_chain[69] ;
 wire \thechain[2].chain9.inv_chain[6] ;
 wire \thechain[2].chain9.inv_chain[70] ;
 wire \thechain[2].chain9.inv_chain[71] ;
 wire \thechain[2].chain9.inv_chain[72] ;
 wire \thechain[2].chain9.inv_chain[73] ;
 wire \thechain[2].chain9.inv_chain[74] ;
 wire \thechain[2].chain9.inv_chain[75] ;
 wire \thechain[2].chain9.inv_chain[76] ;
 wire \thechain[2].chain9.inv_chain[77] ;
 wire \thechain[2].chain9.inv_chain[78] ;
 wire \thechain[2].chain9.inv_chain[79] ;
 wire \thechain[2].chain9.inv_chain[7] ;
 wire \thechain[2].chain9.inv_chain[80] ;
 wire \thechain[2].chain9.inv_chain[81] ;
 wire \thechain[2].chain9.inv_chain[82] ;
 wire \thechain[2].chain9.inv_chain[83] ;
 wire \thechain[2].chain9.inv_chain[84] ;
 wire \thechain[2].chain9.inv_chain[85] ;
 wire \thechain[2].chain9.inv_chain[86] ;
 wire \thechain[2].chain9.inv_chain[87] ;
 wire \thechain[2].chain9.inv_chain[88] ;
 wire \thechain[2].chain9.inv_chain[89] ;
 wire \thechain[2].chain9.inv_chain[8] ;
 wire \thechain[2].chain9.inv_chain[90] ;
 wire \thechain[2].chain9.inv_chain[91] ;
 wire \thechain[2].chain9.inv_chain[92] ;
 wire \thechain[2].chain9.inv_chain[93] ;
 wire \thechain[2].chain9.inv_chain[94] ;
 wire \thechain[2].chain9.inv_chain[95] ;
 wire \thechain[2].chain9.inv_chain[96] ;
 wire \thechain[2].chain9.inv_chain[97] ;
 wire \thechain[2].chain9.inv_chain[98] ;
 wire \thechain[2].chain9.inv_chain[99] ;
 wire \thechain[2].chain9.inv_chain[9] ;
 wire \thechain[3].chain1.dout ;
 wire \thechain[3].chain1.inv_chain[0] ;
 wire \thechain[3].chain1.inv_chain[1] ;
 wire \thechain[3].chain1.inv_chain[2] ;
 wire \thechain[3].chain2.dout ;
 wire \thechain[3].chain2.inv_chain[0] ;
 wire \thechain[3].chain2.inv_chain[1] ;
 wire \thechain[3].chain2.inv_chain[2] ;
 wire \thechain[3].chain2.inv_chain[3] ;
 wire \thechain[3].chain2.inv_chain[4] ;
 wire \thechain[3].chain3.dout ;
 wire \thechain[3].chain3.inv_chain[0] ;
 wire \thechain[3].chain3.inv_chain[1] ;
 wire \thechain[3].chain3.inv_chain[2] ;
 wire \thechain[3].chain3.inv_chain[3] ;
 wire \thechain[3].chain3.inv_chain[4] ;
 wire \thechain[3].chain3.inv_chain[5] ;
 wire \thechain[3].chain3.inv_chain[6] ;
 wire \thechain[3].chain3.inv_chain[7] ;
 wire \thechain[3].chain3.inv_chain[8] ;
 wire \thechain[3].chain4.dout ;
 wire \thechain[3].chain4.inv_chain[0] ;
 wire \thechain[3].chain4.inv_chain[10] ;
 wire \thechain[3].chain4.inv_chain[11] ;
 wire \thechain[3].chain4.inv_chain[12] ;
 wire \thechain[3].chain4.inv_chain[13] ;
 wire \thechain[3].chain4.inv_chain[14] ;
 wire \thechain[3].chain4.inv_chain[15] ;
 wire \thechain[3].chain4.inv_chain[16] ;
 wire \thechain[3].chain4.inv_chain[1] ;
 wire \thechain[3].chain4.inv_chain[2] ;
 wire \thechain[3].chain4.inv_chain[3] ;
 wire \thechain[3].chain4.inv_chain[4] ;
 wire \thechain[3].chain4.inv_chain[5] ;
 wire \thechain[3].chain4.inv_chain[6] ;
 wire \thechain[3].chain4.inv_chain[7] ;
 wire \thechain[3].chain4.inv_chain[8] ;
 wire \thechain[3].chain4.inv_chain[9] ;
 wire \thechain[3].chain5.dout ;
 wire \thechain[3].chain5.inv_chain[0] ;
 wire \thechain[3].chain5.inv_chain[10] ;
 wire \thechain[3].chain5.inv_chain[11] ;
 wire \thechain[3].chain5.inv_chain[12] ;
 wire \thechain[3].chain5.inv_chain[13] ;
 wire \thechain[3].chain5.inv_chain[14] ;
 wire \thechain[3].chain5.inv_chain[15] ;
 wire \thechain[3].chain5.inv_chain[16] ;
 wire \thechain[3].chain5.inv_chain[17] ;
 wire \thechain[3].chain5.inv_chain[18] ;
 wire \thechain[3].chain5.inv_chain[19] ;
 wire \thechain[3].chain5.inv_chain[1] ;
 wire \thechain[3].chain5.inv_chain[20] ;
 wire \thechain[3].chain5.inv_chain[21] ;
 wire \thechain[3].chain5.inv_chain[22] ;
 wire \thechain[3].chain5.inv_chain[23] ;
 wire \thechain[3].chain5.inv_chain[24] ;
 wire \thechain[3].chain5.inv_chain[25] ;
 wire \thechain[3].chain5.inv_chain[26] ;
 wire \thechain[3].chain5.inv_chain[27] ;
 wire \thechain[3].chain5.inv_chain[28] ;
 wire \thechain[3].chain5.inv_chain[29] ;
 wire \thechain[3].chain5.inv_chain[2] ;
 wire \thechain[3].chain5.inv_chain[30] ;
 wire \thechain[3].chain5.inv_chain[31] ;
 wire \thechain[3].chain5.inv_chain[32] ;
 wire \thechain[3].chain5.inv_chain[3] ;
 wire \thechain[3].chain5.inv_chain[4] ;
 wire \thechain[3].chain5.inv_chain[5] ;
 wire \thechain[3].chain5.inv_chain[6] ;
 wire \thechain[3].chain5.inv_chain[7] ;
 wire \thechain[3].chain5.inv_chain[8] ;
 wire \thechain[3].chain5.inv_chain[9] ;
 wire \thechain[3].chain6.dout ;
 wire \thechain[3].chain6.inv_chain[0] ;
 wire \thechain[3].chain6.inv_chain[10] ;
 wire \thechain[3].chain6.inv_chain[11] ;
 wire \thechain[3].chain6.inv_chain[12] ;
 wire \thechain[3].chain6.inv_chain[13] ;
 wire \thechain[3].chain6.inv_chain[14] ;
 wire \thechain[3].chain6.inv_chain[15] ;
 wire \thechain[3].chain6.inv_chain[16] ;
 wire \thechain[3].chain6.inv_chain[17] ;
 wire \thechain[3].chain6.inv_chain[18] ;
 wire \thechain[3].chain6.inv_chain[19] ;
 wire \thechain[3].chain6.inv_chain[1] ;
 wire \thechain[3].chain6.inv_chain[20] ;
 wire \thechain[3].chain6.inv_chain[21] ;
 wire \thechain[3].chain6.inv_chain[22] ;
 wire \thechain[3].chain6.inv_chain[23] ;
 wire \thechain[3].chain6.inv_chain[24] ;
 wire \thechain[3].chain6.inv_chain[25] ;
 wire \thechain[3].chain6.inv_chain[26] ;
 wire \thechain[3].chain6.inv_chain[27] ;
 wire \thechain[3].chain6.inv_chain[28] ;
 wire \thechain[3].chain6.inv_chain[29] ;
 wire \thechain[3].chain6.inv_chain[2] ;
 wire \thechain[3].chain6.inv_chain[30] ;
 wire \thechain[3].chain6.inv_chain[31] ;
 wire \thechain[3].chain6.inv_chain[32] ;
 wire \thechain[3].chain6.inv_chain[33] ;
 wire \thechain[3].chain6.inv_chain[34] ;
 wire \thechain[3].chain6.inv_chain[35] ;
 wire \thechain[3].chain6.inv_chain[36] ;
 wire \thechain[3].chain6.inv_chain[37] ;
 wire \thechain[3].chain6.inv_chain[38] ;
 wire \thechain[3].chain6.inv_chain[39] ;
 wire \thechain[3].chain6.inv_chain[3] ;
 wire \thechain[3].chain6.inv_chain[40] ;
 wire \thechain[3].chain6.inv_chain[41] ;
 wire \thechain[3].chain6.inv_chain[42] ;
 wire \thechain[3].chain6.inv_chain[43] ;
 wire \thechain[3].chain6.inv_chain[44] ;
 wire \thechain[3].chain6.inv_chain[45] ;
 wire \thechain[3].chain6.inv_chain[46] ;
 wire \thechain[3].chain6.inv_chain[47] ;
 wire \thechain[3].chain6.inv_chain[48] ;
 wire \thechain[3].chain6.inv_chain[49] ;
 wire \thechain[3].chain6.inv_chain[4] ;
 wire \thechain[3].chain6.inv_chain[50] ;
 wire \thechain[3].chain6.inv_chain[51] ;
 wire \thechain[3].chain6.inv_chain[52] ;
 wire \thechain[3].chain6.inv_chain[53] ;
 wire \thechain[3].chain6.inv_chain[54] ;
 wire \thechain[3].chain6.inv_chain[55] ;
 wire \thechain[3].chain6.inv_chain[56] ;
 wire \thechain[3].chain6.inv_chain[57] ;
 wire \thechain[3].chain6.inv_chain[58] ;
 wire \thechain[3].chain6.inv_chain[59] ;
 wire \thechain[3].chain6.inv_chain[5] ;
 wire \thechain[3].chain6.inv_chain[60] ;
 wire \thechain[3].chain6.inv_chain[61] ;
 wire \thechain[3].chain6.inv_chain[62] ;
 wire \thechain[3].chain6.inv_chain[63] ;
 wire \thechain[3].chain6.inv_chain[64] ;
 wire \thechain[3].chain6.inv_chain[6] ;
 wire \thechain[3].chain6.inv_chain[7] ;
 wire \thechain[3].chain6.inv_chain[8] ;
 wire \thechain[3].chain6.inv_chain[9] ;
 wire \thechain[3].chain7.dout ;
 wire \thechain[3].chain7.inv_chain[0] ;
 wire \thechain[3].chain7.inv_chain[100] ;
 wire \thechain[3].chain7.inv_chain[101] ;
 wire \thechain[3].chain7.inv_chain[102] ;
 wire \thechain[3].chain7.inv_chain[103] ;
 wire \thechain[3].chain7.inv_chain[104] ;
 wire \thechain[3].chain7.inv_chain[105] ;
 wire \thechain[3].chain7.inv_chain[106] ;
 wire \thechain[3].chain7.inv_chain[107] ;
 wire \thechain[3].chain7.inv_chain[108] ;
 wire \thechain[3].chain7.inv_chain[109] ;
 wire \thechain[3].chain7.inv_chain[10] ;
 wire \thechain[3].chain7.inv_chain[110] ;
 wire \thechain[3].chain7.inv_chain[111] ;
 wire \thechain[3].chain7.inv_chain[112] ;
 wire \thechain[3].chain7.inv_chain[113] ;
 wire \thechain[3].chain7.inv_chain[114] ;
 wire \thechain[3].chain7.inv_chain[115] ;
 wire \thechain[3].chain7.inv_chain[116] ;
 wire \thechain[3].chain7.inv_chain[117] ;
 wire \thechain[3].chain7.inv_chain[118] ;
 wire \thechain[3].chain7.inv_chain[119] ;
 wire \thechain[3].chain7.inv_chain[11] ;
 wire \thechain[3].chain7.inv_chain[120] ;
 wire \thechain[3].chain7.inv_chain[121] ;
 wire \thechain[3].chain7.inv_chain[122] ;
 wire \thechain[3].chain7.inv_chain[123] ;
 wire \thechain[3].chain7.inv_chain[124] ;
 wire \thechain[3].chain7.inv_chain[125] ;
 wire \thechain[3].chain7.inv_chain[126] ;
 wire \thechain[3].chain7.inv_chain[127] ;
 wire \thechain[3].chain7.inv_chain[128] ;
 wire \thechain[3].chain7.inv_chain[12] ;
 wire \thechain[3].chain7.inv_chain[13] ;
 wire \thechain[3].chain7.inv_chain[14] ;
 wire \thechain[3].chain7.inv_chain[15] ;
 wire \thechain[3].chain7.inv_chain[16] ;
 wire \thechain[3].chain7.inv_chain[17] ;
 wire \thechain[3].chain7.inv_chain[18] ;
 wire \thechain[3].chain7.inv_chain[19] ;
 wire \thechain[3].chain7.inv_chain[1] ;
 wire \thechain[3].chain7.inv_chain[20] ;
 wire \thechain[3].chain7.inv_chain[21] ;
 wire \thechain[3].chain7.inv_chain[22] ;
 wire \thechain[3].chain7.inv_chain[23] ;
 wire \thechain[3].chain7.inv_chain[24] ;
 wire \thechain[3].chain7.inv_chain[25] ;
 wire \thechain[3].chain7.inv_chain[26] ;
 wire \thechain[3].chain7.inv_chain[27] ;
 wire \thechain[3].chain7.inv_chain[28] ;
 wire \thechain[3].chain7.inv_chain[29] ;
 wire \thechain[3].chain7.inv_chain[2] ;
 wire \thechain[3].chain7.inv_chain[30] ;
 wire \thechain[3].chain7.inv_chain[31] ;
 wire \thechain[3].chain7.inv_chain[32] ;
 wire \thechain[3].chain7.inv_chain[33] ;
 wire \thechain[3].chain7.inv_chain[34] ;
 wire \thechain[3].chain7.inv_chain[35] ;
 wire \thechain[3].chain7.inv_chain[36] ;
 wire \thechain[3].chain7.inv_chain[37] ;
 wire \thechain[3].chain7.inv_chain[38] ;
 wire \thechain[3].chain7.inv_chain[39] ;
 wire \thechain[3].chain7.inv_chain[3] ;
 wire \thechain[3].chain7.inv_chain[40] ;
 wire \thechain[3].chain7.inv_chain[41] ;
 wire \thechain[3].chain7.inv_chain[42] ;
 wire \thechain[3].chain7.inv_chain[43] ;
 wire \thechain[3].chain7.inv_chain[44] ;
 wire \thechain[3].chain7.inv_chain[45] ;
 wire \thechain[3].chain7.inv_chain[46] ;
 wire \thechain[3].chain7.inv_chain[47] ;
 wire \thechain[3].chain7.inv_chain[48] ;
 wire \thechain[3].chain7.inv_chain[49] ;
 wire \thechain[3].chain7.inv_chain[4] ;
 wire \thechain[3].chain7.inv_chain[50] ;
 wire \thechain[3].chain7.inv_chain[51] ;
 wire \thechain[3].chain7.inv_chain[52] ;
 wire \thechain[3].chain7.inv_chain[53] ;
 wire \thechain[3].chain7.inv_chain[54] ;
 wire \thechain[3].chain7.inv_chain[55] ;
 wire \thechain[3].chain7.inv_chain[56] ;
 wire \thechain[3].chain7.inv_chain[57] ;
 wire \thechain[3].chain7.inv_chain[58] ;
 wire \thechain[3].chain7.inv_chain[59] ;
 wire \thechain[3].chain7.inv_chain[5] ;
 wire \thechain[3].chain7.inv_chain[60] ;
 wire \thechain[3].chain7.inv_chain[61] ;
 wire \thechain[3].chain7.inv_chain[62] ;
 wire \thechain[3].chain7.inv_chain[63] ;
 wire \thechain[3].chain7.inv_chain[64] ;
 wire \thechain[3].chain7.inv_chain[65] ;
 wire \thechain[3].chain7.inv_chain[66] ;
 wire \thechain[3].chain7.inv_chain[67] ;
 wire \thechain[3].chain7.inv_chain[68] ;
 wire \thechain[3].chain7.inv_chain[69] ;
 wire \thechain[3].chain7.inv_chain[6] ;
 wire \thechain[3].chain7.inv_chain[70] ;
 wire \thechain[3].chain7.inv_chain[71] ;
 wire \thechain[3].chain7.inv_chain[72] ;
 wire \thechain[3].chain7.inv_chain[73] ;
 wire \thechain[3].chain7.inv_chain[74] ;
 wire \thechain[3].chain7.inv_chain[75] ;
 wire \thechain[3].chain7.inv_chain[76] ;
 wire \thechain[3].chain7.inv_chain[77] ;
 wire \thechain[3].chain7.inv_chain[78] ;
 wire \thechain[3].chain7.inv_chain[79] ;
 wire \thechain[3].chain7.inv_chain[7] ;
 wire \thechain[3].chain7.inv_chain[80] ;
 wire \thechain[3].chain7.inv_chain[81] ;
 wire \thechain[3].chain7.inv_chain[82] ;
 wire \thechain[3].chain7.inv_chain[83] ;
 wire \thechain[3].chain7.inv_chain[84] ;
 wire \thechain[3].chain7.inv_chain[85] ;
 wire \thechain[3].chain7.inv_chain[86] ;
 wire \thechain[3].chain7.inv_chain[87] ;
 wire \thechain[3].chain7.inv_chain[88] ;
 wire \thechain[3].chain7.inv_chain[89] ;
 wire \thechain[3].chain7.inv_chain[8] ;
 wire \thechain[3].chain7.inv_chain[90] ;
 wire \thechain[3].chain7.inv_chain[91] ;
 wire \thechain[3].chain7.inv_chain[92] ;
 wire \thechain[3].chain7.inv_chain[93] ;
 wire \thechain[3].chain7.inv_chain[94] ;
 wire \thechain[3].chain7.inv_chain[95] ;
 wire \thechain[3].chain7.inv_chain[96] ;
 wire \thechain[3].chain7.inv_chain[97] ;
 wire \thechain[3].chain7.inv_chain[98] ;
 wire \thechain[3].chain7.inv_chain[99] ;
 wire \thechain[3].chain7.inv_chain[9] ;
 wire \thechain[3].chain8.dout ;
 wire \thechain[3].chain8.inv_chain[0] ;
 wire \thechain[3].chain8.inv_chain[100] ;
 wire \thechain[3].chain8.inv_chain[101] ;
 wire \thechain[3].chain8.inv_chain[102] ;
 wire \thechain[3].chain8.inv_chain[103] ;
 wire \thechain[3].chain8.inv_chain[104] ;
 wire \thechain[3].chain8.inv_chain[105] ;
 wire \thechain[3].chain8.inv_chain[106] ;
 wire \thechain[3].chain8.inv_chain[107] ;
 wire \thechain[3].chain8.inv_chain[108] ;
 wire \thechain[3].chain8.inv_chain[109] ;
 wire \thechain[3].chain8.inv_chain[10] ;
 wire \thechain[3].chain8.inv_chain[110] ;
 wire \thechain[3].chain8.inv_chain[111] ;
 wire \thechain[3].chain8.inv_chain[112] ;
 wire \thechain[3].chain8.inv_chain[113] ;
 wire \thechain[3].chain8.inv_chain[114] ;
 wire \thechain[3].chain8.inv_chain[115] ;
 wire \thechain[3].chain8.inv_chain[116] ;
 wire \thechain[3].chain8.inv_chain[117] ;
 wire \thechain[3].chain8.inv_chain[118] ;
 wire \thechain[3].chain8.inv_chain[119] ;
 wire \thechain[3].chain8.inv_chain[11] ;
 wire \thechain[3].chain8.inv_chain[120] ;
 wire \thechain[3].chain8.inv_chain[121] ;
 wire \thechain[3].chain8.inv_chain[122] ;
 wire \thechain[3].chain8.inv_chain[123] ;
 wire \thechain[3].chain8.inv_chain[124] ;
 wire \thechain[3].chain8.inv_chain[125] ;
 wire \thechain[3].chain8.inv_chain[126] ;
 wire \thechain[3].chain8.inv_chain[127] ;
 wire \thechain[3].chain8.inv_chain[128] ;
 wire \thechain[3].chain8.inv_chain[129] ;
 wire \thechain[3].chain8.inv_chain[12] ;
 wire \thechain[3].chain8.inv_chain[130] ;
 wire \thechain[3].chain8.inv_chain[131] ;
 wire \thechain[3].chain8.inv_chain[132] ;
 wire \thechain[3].chain8.inv_chain[133] ;
 wire \thechain[3].chain8.inv_chain[134] ;
 wire \thechain[3].chain8.inv_chain[135] ;
 wire \thechain[3].chain8.inv_chain[136] ;
 wire \thechain[3].chain8.inv_chain[137] ;
 wire \thechain[3].chain8.inv_chain[138] ;
 wire \thechain[3].chain8.inv_chain[139] ;
 wire \thechain[3].chain8.inv_chain[13] ;
 wire \thechain[3].chain8.inv_chain[140] ;
 wire \thechain[3].chain8.inv_chain[141] ;
 wire \thechain[3].chain8.inv_chain[142] ;
 wire \thechain[3].chain8.inv_chain[143] ;
 wire \thechain[3].chain8.inv_chain[144] ;
 wire \thechain[3].chain8.inv_chain[145] ;
 wire \thechain[3].chain8.inv_chain[146] ;
 wire \thechain[3].chain8.inv_chain[147] ;
 wire \thechain[3].chain8.inv_chain[148] ;
 wire \thechain[3].chain8.inv_chain[149] ;
 wire \thechain[3].chain8.inv_chain[14] ;
 wire \thechain[3].chain8.inv_chain[150] ;
 wire \thechain[3].chain8.inv_chain[151] ;
 wire \thechain[3].chain8.inv_chain[152] ;
 wire \thechain[3].chain8.inv_chain[153] ;
 wire \thechain[3].chain8.inv_chain[154] ;
 wire \thechain[3].chain8.inv_chain[155] ;
 wire \thechain[3].chain8.inv_chain[156] ;
 wire \thechain[3].chain8.inv_chain[157] ;
 wire \thechain[3].chain8.inv_chain[158] ;
 wire \thechain[3].chain8.inv_chain[159] ;
 wire \thechain[3].chain8.inv_chain[15] ;
 wire \thechain[3].chain8.inv_chain[160] ;
 wire \thechain[3].chain8.inv_chain[161] ;
 wire \thechain[3].chain8.inv_chain[162] ;
 wire \thechain[3].chain8.inv_chain[163] ;
 wire \thechain[3].chain8.inv_chain[164] ;
 wire \thechain[3].chain8.inv_chain[165] ;
 wire \thechain[3].chain8.inv_chain[166] ;
 wire \thechain[3].chain8.inv_chain[167] ;
 wire \thechain[3].chain8.inv_chain[168] ;
 wire \thechain[3].chain8.inv_chain[169] ;
 wire \thechain[3].chain8.inv_chain[16] ;
 wire \thechain[3].chain8.inv_chain[170] ;
 wire \thechain[3].chain8.inv_chain[171] ;
 wire \thechain[3].chain8.inv_chain[172] ;
 wire \thechain[3].chain8.inv_chain[173] ;
 wire \thechain[3].chain8.inv_chain[174] ;
 wire \thechain[3].chain8.inv_chain[175] ;
 wire \thechain[3].chain8.inv_chain[176] ;
 wire \thechain[3].chain8.inv_chain[177] ;
 wire \thechain[3].chain8.inv_chain[178] ;
 wire \thechain[3].chain8.inv_chain[179] ;
 wire \thechain[3].chain8.inv_chain[17] ;
 wire \thechain[3].chain8.inv_chain[180] ;
 wire \thechain[3].chain8.inv_chain[181] ;
 wire \thechain[3].chain8.inv_chain[182] ;
 wire \thechain[3].chain8.inv_chain[183] ;
 wire \thechain[3].chain8.inv_chain[184] ;
 wire \thechain[3].chain8.inv_chain[185] ;
 wire \thechain[3].chain8.inv_chain[186] ;
 wire \thechain[3].chain8.inv_chain[187] ;
 wire \thechain[3].chain8.inv_chain[188] ;
 wire \thechain[3].chain8.inv_chain[189] ;
 wire \thechain[3].chain8.inv_chain[18] ;
 wire \thechain[3].chain8.inv_chain[190] ;
 wire \thechain[3].chain8.inv_chain[191] ;
 wire \thechain[3].chain8.inv_chain[192] ;
 wire \thechain[3].chain8.inv_chain[19] ;
 wire \thechain[3].chain8.inv_chain[1] ;
 wire \thechain[3].chain8.inv_chain[20] ;
 wire \thechain[3].chain8.inv_chain[21] ;
 wire \thechain[3].chain8.inv_chain[22] ;
 wire \thechain[3].chain8.inv_chain[23] ;
 wire \thechain[3].chain8.inv_chain[24] ;
 wire \thechain[3].chain8.inv_chain[25] ;
 wire \thechain[3].chain8.inv_chain[26] ;
 wire \thechain[3].chain8.inv_chain[27] ;
 wire \thechain[3].chain8.inv_chain[28] ;
 wire \thechain[3].chain8.inv_chain[29] ;
 wire \thechain[3].chain8.inv_chain[2] ;
 wire \thechain[3].chain8.inv_chain[30] ;
 wire \thechain[3].chain8.inv_chain[31] ;
 wire \thechain[3].chain8.inv_chain[32] ;
 wire \thechain[3].chain8.inv_chain[33] ;
 wire \thechain[3].chain8.inv_chain[34] ;
 wire \thechain[3].chain8.inv_chain[35] ;
 wire \thechain[3].chain8.inv_chain[36] ;
 wire \thechain[3].chain8.inv_chain[37] ;
 wire \thechain[3].chain8.inv_chain[38] ;
 wire \thechain[3].chain8.inv_chain[39] ;
 wire \thechain[3].chain8.inv_chain[3] ;
 wire \thechain[3].chain8.inv_chain[40] ;
 wire \thechain[3].chain8.inv_chain[41] ;
 wire \thechain[3].chain8.inv_chain[42] ;
 wire \thechain[3].chain8.inv_chain[43] ;
 wire \thechain[3].chain8.inv_chain[44] ;
 wire \thechain[3].chain8.inv_chain[45] ;
 wire \thechain[3].chain8.inv_chain[46] ;
 wire \thechain[3].chain8.inv_chain[47] ;
 wire \thechain[3].chain8.inv_chain[48] ;
 wire \thechain[3].chain8.inv_chain[49] ;
 wire \thechain[3].chain8.inv_chain[4] ;
 wire \thechain[3].chain8.inv_chain[50] ;
 wire \thechain[3].chain8.inv_chain[51] ;
 wire \thechain[3].chain8.inv_chain[52] ;
 wire \thechain[3].chain8.inv_chain[53] ;
 wire \thechain[3].chain8.inv_chain[54] ;
 wire \thechain[3].chain8.inv_chain[55] ;
 wire \thechain[3].chain8.inv_chain[56] ;
 wire \thechain[3].chain8.inv_chain[57] ;
 wire \thechain[3].chain8.inv_chain[58] ;
 wire \thechain[3].chain8.inv_chain[59] ;
 wire \thechain[3].chain8.inv_chain[5] ;
 wire \thechain[3].chain8.inv_chain[60] ;
 wire \thechain[3].chain8.inv_chain[61] ;
 wire \thechain[3].chain8.inv_chain[62] ;
 wire \thechain[3].chain8.inv_chain[63] ;
 wire \thechain[3].chain8.inv_chain[64] ;
 wire \thechain[3].chain8.inv_chain[65] ;
 wire \thechain[3].chain8.inv_chain[66] ;
 wire \thechain[3].chain8.inv_chain[67] ;
 wire \thechain[3].chain8.inv_chain[68] ;
 wire \thechain[3].chain8.inv_chain[69] ;
 wire \thechain[3].chain8.inv_chain[6] ;
 wire \thechain[3].chain8.inv_chain[70] ;
 wire \thechain[3].chain8.inv_chain[71] ;
 wire \thechain[3].chain8.inv_chain[72] ;
 wire \thechain[3].chain8.inv_chain[73] ;
 wire \thechain[3].chain8.inv_chain[74] ;
 wire \thechain[3].chain8.inv_chain[75] ;
 wire \thechain[3].chain8.inv_chain[76] ;
 wire \thechain[3].chain8.inv_chain[77] ;
 wire \thechain[3].chain8.inv_chain[78] ;
 wire \thechain[3].chain8.inv_chain[79] ;
 wire \thechain[3].chain8.inv_chain[7] ;
 wire \thechain[3].chain8.inv_chain[80] ;
 wire \thechain[3].chain8.inv_chain[81] ;
 wire \thechain[3].chain8.inv_chain[82] ;
 wire \thechain[3].chain8.inv_chain[83] ;
 wire \thechain[3].chain8.inv_chain[84] ;
 wire \thechain[3].chain8.inv_chain[85] ;
 wire \thechain[3].chain8.inv_chain[86] ;
 wire \thechain[3].chain8.inv_chain[87] ;
 wire \thechain[3].chain8.inv_chain[88] ;
 wire \thechain[3].chain8.inv_chain[89] ;
 wire \thechain[3].chain8.inv_chain[8] ;
 wire \thechain[3].chain8.inv_chain[90] ;
 wire \thechain[3].chain8.inv_chain[91] ;
 wire \thechain[3].chain8.inv_chain[92] ;
 wire \thechain[3].chain8.inv_chain[93] ;
 wire \thechain[3].chain8.inv_chain[94] ;
 wire \thechain[3].chain8.inv_chain[95] ;
 wire \thechain[3].chain8.inv_chain[96] ;
 wire \thechain[3].chain8.inv_chain[97] ;
 wire \thechain[3].chain8.inv_chain[98] ;
 wire \thechain[3].chain8.inv_chain[99] ;
 wire \thechain[3].chain8.inv_chain[9] ;
 wire \thechain[3].chain9.dout ;
 wire \thechain[3].chain9.inv_chain[0] ;
 wire \thechain[3].chain9.inv_chain[100] ;
 wire \thechain[3].chain9.inv_chain[101] ;
 wire \thechain[3].chain9.inv_chain[102] ;
 wire \thechain[3].chain9.inv_chain[103] ;
 wire \thechain[3].chain9.inv_chain[104] ;
 wire \thechain[3].chain9.inv_chain[105] ;
 wire \thechain[3].chain9.inv_chain[106] ;
 wire \thechain[3].chain9.inv_chain[107] ;
 wire \thechain[3].chain9.inv_chain[108] ;
 wire \thechain[3].chain9.inv_chain[109] ;
 wire \thechain[3].chain9.inv_chain[10] ;
 wire \thechain[3].chain9.inv_chain[110] ;
 wire \thechain[3].chain9.inv_chain[111] ;
 wire \thechain[3].chain9.inv_chain[112] ;
 wire \thechain[3].chain9.inv_chain[113] ;
 wire \thechain[3].chain9.inv_chain[114] ;
 wire \thechain[3].chain9.inv_chain[115] ;
 wire \thechain[3].chain9.inv_chain[116] ;
 wire \thechain[3].chain9.inv_chain[117] ;
 wire \thechain[3].chain9.inv_chain[118] ;
 wire \thechain[3].chain9.inv_chain[119] ;
 wire \thechain[3].chain9.inv_chain[11] ;
 wire \thechain[3].chain9.inv_chain[120] ;
 wire \thechain[3].chain9.inv_chain[121] ;
 wire \thechain[3].chain9.inv_chain[122] ;
 wire \thechain[3].chain9.inv_chain[123] ;
 wire \thechain[3].chain9.inv_chain[124] ;
 wire \thechain[3].chain9.inv_chain[125] ;
 wire \thechain[3].chain9.inv_chain[126] ;
 wire \thechain[3].chain9.inv_chain[127] ;
 wire \thechain[3].chain9.inv_chain[128] ;
 wire \thechain[3].chain9.inv_chain[129] ;
 wire \thechain[3].chain9.inv_chain[12] ;
 wire \thechain[3].chain9.inv_chain[130] ;
 wire \thechain[3].chain9.inv_chain[131] ;
 wire \thechain[3].chain9.inv_chain[132] ;
 wire \thechain[3].chain9.inv_chain[133] ;
 wire \thechain[3].chain9.inv_chain[134] ;
 wire \thechain[3].chain9.inv_chain[135] ;
 wire \thechain[3].chain9.inv_chain[136] ;
 wire \thechain[3].chain9.inv_chain[137] ;
 wire \thechain[3].chain9.inv_chain[138] ;
 wire \thechain[3].chain9.inv_chain[139] ;
 wire \thechain[3].chain9.inv_chain[13] ;
 wire \thechain[3].chain9.inv_chain[140] ;
 wire \thechain[3].chain9.inv_chain[141] ;
 wire \thechain[3].chain9.inv_chain[142] ;
 wire \thechain[3].chain9.inv_chain[143] ;
 wire \thechain[3].chain9.inv_chain[144] ;
 wire \thechain[3].chain9.inv_chain[145] ;
 wire \thechain[3].chain9.inv_chain[146] ;
 wire \thechain[3].chain9.inv_chain[147] ;
 wire \thechain[3].chain9.inv_chain[148] ;
 wire \thechain[3].chain9.inv_chain[149] ;
 wire \thechain[3].chain9.inv_chain[14] ;
 wire \thechain[3].chain9.inv_chain[150] ;
 wire \thechain[3].chain9.inv_chain[151] ;
 wire \thechain[3].chain9.inv_chain[152] ;
 wire \thechain[3].chain9.inv_chain[153] ;
 wire \thechain[3].chain9.inv_chain[154] ;
 wire \thechain[3].chain9.inv_chain[155] ;
 wire \thechain[3].chain9.inv_chain[156] ;
 wire \thechain[3].chain9.inv_chain[157] ;
 wire \thechain[3].chain9.inv_chain[158] ;
 wire \thechain[3].chain9.inv_chain[159] ;
 wire \thechain[3].chain9.inv_chain[15] ;
 wire \thechain[3].chain9.inv_chain[160] ;
 wire \thechain[3].chain9.inv_chain[161] ;
 wire \thechain[3].chain9.inv_chain[162] ;
 wire \thechain[3].chain9.inv_chain[163] ;
 wire \thechain[3].chain9.inv_chain[164] ;
 wire \thechain[3].chain9.inv_chain[165] ;
 wire \thechain[3].chain9.inv_chain[166] ;
 wire \thechain[3].chain9.inv_chain[167] ;
 wire \thechain[3].chain9.inv_chain[168] ;
 wire \thechain[3].chain9.inv_chain[169] ;
 wire \thechain[3].chain9.inv_chain[16] ;
 wire \thechain[3].chain9.inv_chain[170] ;
 wire \thechain[3].chain9.inv_chain[171] ;
 wire \thechain[3].chain9.inv_chain[172] ;
 wire \thechain[3].chain9.inv_chain[173] ;
 wire \thechain[3].chain9.inv_chain[174] ;
 wire \thechain[3].chain9.inv_chain[175] ;
 wire \thechain[3].chain9.inv_chain[176] ;
 wire \thechain[3].chain9.inv_chain[177] ;
 wire \thechain[3].chain9.inv_chain[178] ;
 wire \thechain[3].chain9.inv_chain[179] ;
 wire \thechain[3].chain9.inv_chain[17] ;
 wire \thechain[3].chain9.inv_chain[180] ;
 wire \thechain[3].chain9.inv_chain[181] ;
 wire \thechain[3].chain9.inv_chain[182] ;
 wire \thechain[3].chain9.inv_chain[183] ;
 wire \thechain[3].chain9.inv_chain[184] ;
 wire \thechain[3].chain9.inv_chain[185] ;
 wire \thechain[3].chain9.inv_chain[186] ;
 wire \thechain[3].chain9.inv_chain[187] ;
 wire \thechain[3].chain9.inv_chain[188] ;
 wire \thechain[3].chain9.inv_chain[189] ;
 wire \thechain[3].chain9.inv_chain[18] ;
 wire \thechain[3].chain9.inv_chain[190] ;
 wire \thechain[3].chain9.inv_chain[191] ;
 wire \thechain[3].chain9.inv_chain[192] ;
 wire \thechain[3].chain9.inv_chain[193] ;
 wire \thechain[3].chain9.inv_chain[194] ;
 wire \thechain[3].chain9.inv_chain[195] ;
 wire \thechain[3].chain9.inv_chain[196] ;
 wire \thechain[3].chain9.inv_chain[197] ;
 wire \thechain[3].chain9.inv_chain[198] ;
 wire \thechain[3].chain9.inv_chain[199] ;
 wire \thechain[3].chain9.inv_chain[19] ;
 wire \thechain[3].chain9.inv_chain[1] ;
 wire \thechain[3].chain9.inv_chain[200] ;
 wire \thechain[3].chain9.inv_chain[201] ;
 wire \thechain[3].chain9.inv_chain[202] ;
 wire \thechain[3].chain9.inv_chain[203] ;
 wire \thechain[3].chain9.inv_chain[204] ;
 wire \thechain[3].chain9.inv_chain[205] ;
 wire \thechain[3].chain9.inv_chain[206] ;
 wire \thechain[3].chain9.inv_chain[207] ;
 wire \thechain[3].chain9.inv_chain[208] ;
 wire \thechain[3].chain9.inv_chain[209] ;
 wire \thechain[3].chain9.inv_chain[20] ;
 wire \thechain[3].chain9.inv_chain[210] ;
 wire \thechain[3].chain9.inv_chain[211] ;
 wire \thechain[3].chain9.inv_chain[212] ;
 wire \thechain[3].chain9.inv_chain[213] ;
 wire \thechain[3].chain9.inv_chain[214] ;
 wire \thechain[3].chain9.inv_chain[215] ;
 wire \thechain[3].chain9.inv_chain[216] ;
 wire \thechain[3].chain9.inv_chain[217] ;
 wire \thechain[3].chain9.inv_chain[218] ;
 wire \thechain[3].chain9.inv_chain[219] ;
 wire \thechain[3].chain9.inv_chain[21] ;
 wire \thechain[3].chain9.inv_chain[220] ;
 wire \thechain[3].chain9.inv_chain[221] ;
 wire \thechain[3].chain9.inv_chain[222] ;
 wire \thechain[3].chain9.inv_chain[223] ;
 wire \thechain[3].chain9.inv_chain[224] ;
 wire \thechain[3].chain9.inv_chain[225] ;
 wire \thechain[3].chain9.inv_chain[226] ;
 wire \thechain[3].chain9.inv_chain[227] ;
 wire \thechain[3].chain9.inv_chain[228] ;
 wire \thechain[3].chain9.inv_chain[229] ;
 wire \thechain[3].chain9.inv_chain[22] ;
 wire \thechain[3].chain9.inv_chain[230] ;
 wire \thechain[3].chain9.inv_chain[231] ;
 wire \thechain[3].chain9.inv_chain[232] ;
 wire \thechain[3].chain9.inv_chain[233] ;
 wire \thechain[3].chain9.inv_chain[234] ;
 wire \thechain[3].chain9.inv_chain[235] ;
 wire \thechain[3].chain9.inv_chain[236] ;
 wire \thechain[3].chain9.inv_chain[237] ;
 wire \thechain[3].chain9.inv_chain[238] ;
 wire \thechain[3].chain9.inv_chain[239] ;
 wire \thechain[3].chain9.inv_chain[23] ;
 wire \thechain[3].chain9.inv_chain[240] ;
 wire \thechain[3].chain9.inv_chain[241] ;
 wire \thechain[3].chain9.inv_chain[242] ;
 wire \thechain[3].chain9.inv_chain[243] ;
 wire \thechain[3].chain9.inv_chain[244] ;
 wire \thechain[3].chain9.inv_chain[245] ;
 wire \thechain[3].chain9.inv_chain[246] ;
 wire \thechain[3].chain9.inv_chain[247] ;
 wire \thechain[3].chain9.inv_chain[248] ;
 wire \thechain[3].chain9.inv_chain[249] ;
 wire \thechain[3].chain9.inv_chain[24] ;
 wire \thechain[3].chain9.inv_chain[250] ;
 wire \thechain[3].chain9.inv_chain[251] ;
 wire \thechain[3].chain9.inv_chain[252] ;
 wire \thechain[3].chain9.inv_chain[253] ;
 wire \thechain[3].chain9.inv_chain[254] ;
 wire \thechain[3].chain9.inv_chain[255] ;
 wire \thechain[3].chain9.inv_chain[256] ;
 wire \thechain[3].chain9.inv_chain[25] ;
 wire \thechain[3].chain9.inv_chain[26] ;
 wire \thechain[3].chain9.inv_chain[27] ;
 wire \thechain[3].chain9.inv_chain[28] ;
 wire \thechain[3].chain9.inv_chain[29] ;
 wire \thechain[3].chain9.inv_chain[2] ;
 wire \thechain[3].chain9.inv_chain[30] ;
 wire \thechain[3].chain9.inv_chain[31] ;
 wire \thechain[3].chain9.inv_chain[32] ;
 wire \thechain[3].chain9.inv_chain[33] ;
 wire \thechain[3].chain9.inv_chain[34] ;
 wire \thechain[3].chain9.inv_chain[35] ;
 wire \thechain[3].chain9.inv_chain[36] ;
 wire \thechain[3].chain9.inv_chain[37] ;
 wire \thechain[3].chain9.inv_chain[38] ;
 wire \thechain[3].chain9.inv_chain[39] ;
 wire \thechain[3].chain9.inv_chain[3] ;
 wire \thechain[3].chain9.inv_chain[40] ;
 wire \thechain[3].chain9.inv_chain[41] ;
 wire \thechain[3].chain9.inv_chain[42] ;
 wire \thechain[3].chain9.inv_chain[43] ;
 wire \thechain[3].chain9.inv_chain[44] ;
 wire \thechain[3].chain9.inv_chain[45] ;
 wire \thechain[3].chain9.inv_chain[46] ;
 wire \thechain[3].chain9.inv_chain[47] ;
 wire \thechain[3].chain9.inv_chain[48] ;
 wire \thechain[3].chain9.inv_chain[49] ;
 wire \thechain[3].chain9.inv_chain[4] ;
 wire \thechain[3].chain9.inv_chain[50] ;
 wire \thechain[3].chain9.inv_chain[51] ;
 wire \thechain[3].chain9.inv_chain[52] ;
 wire \thechain[3].chain9.inv_chain[53] ;
 wire \thechain[3].chain9.inv_chain[54] ;
 wire \thechain[3].chain9.inv_chain[55] ;
 wire \thechain[3].chain9.inv_chain[56] ;
 wire \thechain[3].chain9.inv_chain[57] ;
 wire \thechain[3].chain9.inv_chain[58] ;
 wire \thechain[3].chain9.inv_chain[59] ;
 wire \thechain[3].chain9.inv_chain[5] ;
 wire \thechain[3].chain9.inv_chain[60] ;
 wire \thechain[3].chain9.inv_chain[61] ;
 wire \thechain[3].chain9.inv_chain[62] ;
 wire \thechain[3].chain9.inv_chain[63] ;
 wire \thechain[3].chain9.inv_chain[64] ;
 wire \thechain[3].chain9.inv_chain[65] ;
 wire \thechain[3].chain9.inv_chain[66] ;
 wire \thechain[3].chain9.inv_chain[67] ;
 wire \thechain[3].chain9.inv_chain[68] ;
 wire \thechain[3].chain9.inv_chain[69] ;
 wire \thechain[3].chain9.inv_chain[6] ;
 wire \thechain[3].chain9.inv_chain[70] ;
 wire \thechain[3].chain9.inv_chain[71] ;
 wire \thechain[3].chain9.inv_chain[72] ;
 wire \thechain[3].chain9.inv_chain[73] ;
 wire \thechain[3].chain9.inv_chain[74] ;
 wire \thechain[3].chain9.inv_chain[75] ;
 wire \thechain[3].chain9.inv_chain[76] ;
 wire \thechain[3].chain9.inv_chain[77] ;
 wire \thechain[3].chain9.inv_chain[78] ;
 wire \thechain[3].chain9.inv_chain[79] ;
 wire \thechain[3].chain9.inv_chain[7] ;
 wire \thechain[3].chain9.inv_chain[80] ;
 wire \thechain[3].chain9.inv_chain[81] ;
 wire \thechain[3].chain9.inv_chain[82] ;
 wire \thechain[3].chain9.inv_chain[83] ;
 wire \thechain[3].chain9.inv_chain[84] ;
 wire \thechain[3].chain9.inv_chain[85] ;
 wire \thechain[3].chain9.inv_chain[86] ;
 wire \thechain[3].chain9.inv_chain[87] ;
 wire \thechain[3].chain9.inv_chain[88] ;
 wire \thechain[3].chain9.inv_chain[89] ;
 wire \thechain[3].chain9.inv_chain[8] ;
 wire \thechain[3].chain9.inv_chain[90] ;
 wire \thechain[3].chain9.inv_chain[91] ;
 wire \thechain[3].chain9.inv_chain[92] ;
 wire \thechain[3].chain9.inv_chain[93] ;
 wire \thechain[3].chain9.inv_chain[94] ;
 wire \thechain[3].chain9.inv_chain[95] ;
 wire \thechain[3].chain9.inv_chain[96] ;
 wire \thechain[3].chain9.inv_chain[97] ;
 wire \thechain[3].chain9.inv_chain[98] ;
 wire \thechain[3].chain9.inv_chain[99] ;
 wire \thechain[3].chain9.inv_chain[9] ;
 wire \thechain[4].chain1.dout ;
 wire \thechain[4].chain1.inv_chain[0] ;
 wire \thechain[4].chain1.inv_chain[1] ;
 wire \thechain[4].chain1.inv_chain[2] ;
 wire \thechain[4].chain2.dout ;
 wire \thechain[4].chain2.inv_chain[0] ;
 wire \thechain[4].chain2.inv_chain[1] ;
 wire \thechain[4].chain2.inv_chain[2] ;
 wire \thechain[4].chain2.inv_chain[3] ;
 wire \thechain[4].chain2.inv_chain[4] ;
 wire \thechain[4].chain3.dout ;
 wire \thechain[4].chain3.inv_chain[0] ;
 wire \thechain[4].chain3.inv_chain[1] ;
 wire \thechain[4].chain3.inv_chain[2] ;
 wire \thechain[4].chain3.inv_chain[3] ;
 wire \thechain[4].chain3.inv_chain[4] ;
 wire \thechain[4].chain3.inv_chain[5] ;
 wire \thechain[4].chain3.inv_chain[6] ;
 wire \thechain[4].chain3.inv_chain[7] ;
 wire \thechain[4].chain3.inv_chain[8] ;
 wire \thechain[4].chain4.dout ;
 wire \thechain[4].chain4.inv_chain[0] ;
 wire \thechain[4].chain4.inv_chain[10] ;
 wire \thechain[4].chain4.inv_chain[11] ;
 wire \thechain[4].chain4.inv_chain[12] ;
 wire \thechain[4].chain4.inv_chain[13] ;
 wire \thechain[4].chain4.inv_chain[14] ;
 wire \thechain[4].chain4.inv_chain[15] ;
 wire \thechain[4].chain4.inv_chain[16] ;
 wire \thechain[4].chain4.inv_chain[1] ;
 wire \thechain[4].chain4.inv_chain[2] ;
 wire \thechain[4].chain4.inv_chain[3] ;
 wire \thechain[4].chain4.inv_chain[4] ;
 wire \thechain[4].chain4.inv_chain[5] ;
 wire \thechain[4].chain4.inv_chain[6] ;
 wire \thechain[4].chain4.inv_chain[7] ;
 wire \thechain[4].chain4.inv_chain[8] ;
 wire \thechain[4].chain4.inv_chain[9] ;
 wire \thechain[4].chain5.dout ;
 wire \thechain[4].chain5.inv_chain[0] ;
 wire \thechain[4].chain5.inv_chain[10] ;
 wire \thechain[4].chain5.inv_chain[11] ;
 wire \thechain[4].chain5.inv_chain[12] ;
 wire \thechain[4].chain5.inv_chain[13] ;
 wire \thechain[4].chain5.inv_chain[14] ;
 wire \thechain[4].chain5.inv_chain[15] ;
 wire \thechain[4].chain5.inv_chain[16] ;
 wire \thechain[4].chain5.inv_chain[17] ;
 wire \thechain[4].chain5.inv_chain[18] ;
 wire \thechain[4].chain5.inv_chain[19] ;
 wire \thechain[4].chain5.inv_chain[1] ;
 wire \thechain[4].chain5.inv_chain[20] ;
 wire \thechain[4].chain5.inv_chain[21] ;
 wire \thechain[4].chain5.inv_chain[22] ;
 wire \thechain[4].chain5.inv_chain[23] ;
 wire \thechain[4].chain5.inv_chain[24] ;
 wire \thechain[4].chain5.inv_chain[25] ;
 wire \thechain[4].chain5.inv_chain[26] ;
 wire \thechain[4].chain5.inv_chain[27] ;
 wire \thechain[4].chain5.inv_chain[28] ;
 wire \thechain[4].chain5.inv_chain[29] ;
 wire \thechain[4].chain5.inv_chain[2] ;
 wire \thechain[4].chain5.inv_chain[30] ;
 wire \thechain[4].chain5.inv_chain[31] ;
 wire \thechain[4].chain5.inv_chain[32] ;
 wire \thechain[4].chain5.inv_chain[3] ;
 wire \thechain[4].chain5.inv_chain[4] ;
 wire \thechain[4].chain5.inv_chain[5] ;
 wire \thechain[4].chain5.inv_chain[6] ;
 wire \thechain[4].chain5.inv_chain[7] ;
 wire \thechain[4].chain5.inv_chain[8] ;
 wire \thechain[4].chain5.inv_chain[9] ;
 wire \thechain[4].chain6.dout ;
 wire \thechain[4].chain6.inv_chain[0] ;
 wire \thechain[4].chain6.inv_chain[10] ;
 wire \thechain[4].chain6.inv_chain[11] ;
 wire \thechain[4].chain6.inv_chain[12] ;
 wire \thechain[4].chain6.inv_chain[13] ;
 wire \thechain[4].chain6.inv_chain[14] ;
 wire \thechain[4].chain6.inv_chain[15] ;
 wire \thechain[4].chain6.inv_chain[16] ;
 wire \thechain[4].chain6.inv_chain[17] ;
 wire \thechain[4].chain6.inv_chain[18] ;
 wire \thechain[4].chain6.inv_chain[19] ;
 wire \thechain[4].chain6.inv_chain[1] ;
 wire \thechain[4].chain6.inv_chain[20] ;
 wire \thechain[4].chain6.inv_chain[21] ;
 wire \thechain[4].chain6.inv_chain[22] ;
 wire \thechain[4].chain6.inv_chain[23] ;
 wire \thechain[4].chain6.inv_chain[24] ;
 wire \thechain[4].chain6.inv_chain[25] ;
 wire \thechain[4].chain6.inv_chain[26] ;
 wire \thechain[4].chain6.inv_chain[27] ;
 wire \thechain[4].chain6.inv_chain[28] ;
 wire \thechain[4].chain6.inv_chain[29] ;
 wire \thechain[4].chain6.inv_chain[2] ;
 wire \thechain[4].chain6.inv_chain[30] ;
 wire \thechain[4].chain6.inv_chain[31] ;
 wire \thechain[4].chain6.inv_chain[32] ;
 wire \thechain[4].chain6.inv_chain[33] ;
 wire \thechain[4].chain6.inv_chain[34] ;
 wire \thechain[4].chain6.inv_chain[35] ;
 wire \thechain[4].chain6.inv_chain[36] ;
 wire \thechain[4].chain6.inv_chain[37] ;
 wire \thechain[4].chain6.inv_chain[38] ;
 wire \thechain[4].chain6.inv_chain[39] ;
 wire \thechain[4].chain6.inv_chain[3] ;
 wire \thechain[4].chain6.inv_chain[40] ;
 wire \thechain[4].chain6.inv_chain[41] ;
 wire \thechain[4].chain6.inv_chain[42] ;
 wire \thechain[4].chain6.inv_chain[43] ;
 wire \thechain[4].chain6.inv_chain[44] ;
 wire \thechain[4].chain6.inv_chain[45] ;
 wire \thechain[4].chain6.inv_chain[46] ;
 wire \thechain[4].chain6.inv_chain[47] ;
 wire \thechain[4].chain6.inv_chain[48] ;
 wire \thechain[4].chain6.inv_chain[49] ;
 wire \thechain[4].chain6.inv_chain[4] ;
 wire \thechain[4].chain6.inv_chain[50] ;
 wire \thechain[4].chain6.inv_chain[51] ;
 wire \thechain[4].chain6.inv_chain[52] ;
 wire \thechain[4].chain6.inv_chain[53] ;
 wire \thechain[4].chain6.inv_chain[54] ;
 wire \thechain[4].chain6.inv_chain[55] ;
 wire \thechain[4].chain6.inv_chain[56] ;
 wire \thechain[4].chain6.inv_chain[57] ;
 wire \thechain[4].chain6.inv_chain[58] ;
 wire \thechain[4].chain6.inv_chain[59] ;
 wire \thechain[4].chain6.inv_chain[5] ;
 wire \thechain[4].chain6.inv_chain[60] ;
 wire \thechain[4].chain6.inv_chain[61] ;
 wire \thechain[4].chain6.inv_chain[62] ;
 wire \thechain[4].chain6.inv_chain[63] ;
 wire \thechain[4].chain6.inv_chain[64] ;
 wire \thechain[4].chain6.inv_chain[6] ;
 wire \thechain[4].chain6.inv_chain[7] ;
 wire \thechain[4].chain6.inv_chain[8] ;
 wire \thechain[4].chain6.inv_chain[9] ;
 wire \thechain[4].chain7.dout ;
 wire \thechain[4].chain7.inv_chain[0] ;
 wire \thechain[4].chain7.inv_chain[100] ;
 wire \thechain[4].chain7.inv_chain[101] ;
 wire \thechain[4].chain7.inv_chain[102] ;
 wire \thechain[4].chain7.inv_chain[103] ;
 wire \thechain[4].chain7.inv_chain[104] ;
 wire \thechain[4].chain7.inv_chain[105] ;
 wire \thechain[4].chain7.inv_chain[106] ;
 wire \thechain[4].chain7.inv_chain[107] ;
 wire \thechain[4].chain7.inv_chain[108] ;
 wire \thechain[4].chain7.inv_chain[109] ;
 wire \thechain[4].chain7.inv_chain[10] ;
 wire \thechain[4].chain7.inv_chain[110] ;
 wire \thechain[4].chain7.inv_chain[111] ;
 wire \thechain[4].chain7.inv_chain[112] ;
 wire \thechain[4].chain7.inv_chain[113] ;
 wire \thechain[4].chain7.inv_chain[114] ;
 wire \thechain[4].chain7.inv_chain[115] ;
 wire \thechain[4].chain7.inv_chain[116] ;
 wire \thechain[4].chain7.inv_chain[117] ;
 wire \thechain[4].chain7.inv_chain[118] ;
 wire \thechain[4].chain7.inv_chain[119] ;
 wire \thechain[4].chain7.inv_chain[11] ;
 wire \thechain[4].chain7.inv_chain[120] ;
 wire \thechain[4].chain7.inv_chain[121] ;
 wire \thechain[4].chain7.inv_chain[122] ;
 wire \thechain[4].chain7.inv_chain[123] ;
 wire \thechain[4].chain7.inv_chain[124] ;
 wire \thechain[4].chain7.inv_chain[125] ;
 wire \thechain[4].chain7.inv_chain[126] ;
 wire \thechain[4].chain7.inv_chain[127] ;
 wire \thechain[4].chain7.inv_chain[128] ;
 wire \thechain[4].chain7.inv_chain[12] ;
 wire \thechain[4].chain7.inv_chain[13] ;
 wire \thechain[4].chain7.inv_chain[14] ;
 wire \thechain[4].chain7.inv_chain[15] ;
 wire \thechain[4].chain7.inv_chain[16] ;
 wire \thechain[4].chain7.inv_chain[17] ;
 wire \thechain[4].chain7.inv_chain[18] ;
 wire \thechain[4].chain7.inv_chain[19] ;
 wire \thechain[4].chain7.inv_chain[1] ;
 wire \thechain[4].chain7.inv_chain[20] ;
 wire \thechain[4].chain7.inv_chain[21] ;
 wire \thechain[4].chain7.inv_chain[22] ;
 wire \thechain[4].chain7.inv_chain[23] ;
 wire \thechain[4].chain7.inv_chain[24] ;
 wire \thechain[4].chain7.inv_chain[25] ;
 wire \thechain[4].chain7.inv_chain[26] ;
 wire \thechain[4].chain7.inv_chain[27] ;
 wire \thechain[4].chain7.inv_chain[28] ;
 wire \thechain[4].chain7.inv_chain[29] ;
 wire \thechain[4].chain7.inv_chain[2] ;
 wire \thechain[4].chain7.inv_chain[30] ;
 wire \thechain[4].chain7.inv_chain[31] ;
 wire \thechain[4].chain7.inv_chain[32] ;
 wire \thechain[4].chain7.inv_chain[33] ;
 wire \thechain[4].chain7.inv_chain[34] ;
 wire \thechain[4].chain7.inv_chain[35] ;
 wire \thechain[4].chain7.inv_chain[36] ;
 wire \thechain[4].chain7.inv_chain[37] ;
 wire \thechain[4].chain7.inv_chain[38] ;
 wire \thechain[4].chain7.inv_chain[39] ;
 wire \thechain[4].chain7.inv_chain[3] ;
 wire \thechain[4].chain7.inv_chain[40] ;
 wire \thechain[4].chain7.inv_chain[41] ;
 wire \thechain[4].chain7.inv_chain[42] ;
 wire \thechain[4].chain7.inv_chain[43] ;
 wire \thechain[4].chain7.inv_chain[44] ;
 wire \thechain[4].chain7.inv_chain[45] ;
 wire \thechain[4].chain7.inv_chain[46] ;
 wire \thechain[4].chain7.inv_chain[47] ;
 wire \thechain[4].chain7.inv_chain[48] ;
 wire \thechain[4].chain7.inv_chain[49] ;
 wire \thechain[4].chain7.inv_chain[4] ;
 wire \thechain[4].chain7.inv_chain[50] ;
 wire \thechain[4].chain7.inv_chain[51] ;
 wire \thechain[4].chain7.inv_chain[52] ;
 wire \thechain[4].chain7.inv_chain[53] ;
 wire \thechain[4].chain7.inv_chain[54] ;
 wire \thechain[4].chain7.inv_chain[55] ;
 wire \thechain[4].chain7.inv_chain[56] ;
 wire \thechain[4].chain7.inv_chain[57] ;
 wire \thechain[4].chain7.inv_chain[58] ;
 wire \thechain[4].chain7.inv_chain[59] ;
 wire \thechain[4].chain7.inv_chain[5] ;
 wire \thechain[4].chain7.inv_chain[60] ;
 wire \thechain[4].chain7.inv_chain[61] ;
 wire \thechain[4].chain7.inv_chain[62] ;
 wire \thechain[4].chain7.inv_chain[63] ;
 wire \thechain[4].chain7.inv_chain[64] ;
 wire \thechain[4].chain7.inv_chain[65] ;
 wire \thechain[4].chain7.inv_chain[66] ;
 wire \thechain[4].chain7.inv_chain[67] ;
 wire \thechain[4].chain7.inv_chain[68] ;
 wire \thechain[4].chain7.inv_chain[69] ;
 wire \thechain[4].chain7.inv_chain[6] ;
 wire \thechain[4].chain7.inv_chain[70] ;
 wire \thechain[4].chain7.inv_chain[71] ;
 wire \thechain[4].chain7.inv_chain[72] ;
 wire \thechain[4].chain7.inv_chain[73] ;
 wire \thechain[4].chain7.inv_chain[74] ;
 wire \thechain[4].chain7.inv_chain[75] ;
 wire \thechain[4].chain7.inv_chain[76] ;
 wire \thechain[4].chain7.inv_chain[77] ;
 wire \thechain[4].chain7.inv_chain[78] ;
 wire \thechain[4].chain7.inv_chain[79] ;
 wire \thechain[4].chain7.inv_chain[7] ;
 wire \thechain[4].chain7.inv_chain[80] ;
 wire \thechain[4].chain7.inv_chain[81] ;
 wire \thechain[4].chain7.inv_chain[82] ;
 wire \thechain[4].chain7.inv_chain[83] ;
 wire \thechain[4].chain7.inv_chain[84] ;
 wire \thechain[4].chain7.inv_chain[85] ;
 wire \thechain[4].chain7.inv_chain[86] ;
 wire \thechain[4].chain7.inv_chain[87] ;
 wire \thechain[4].chain7.inv_chain[88] ;
 wire \thechain[4].chain7.inv_chain[89] ;
 wire \thechain[4].chain7.inv_chain[8] ;
 wire \thechain[4].chain7.inv_chain[90] ;
 wire \thechain[4].chain7.inv_chain[91] ;
 wire \thechain[4].chain7.inv_chain[92] ;
 wire \thechain[4].chain7.inv_chain[93] ;
 wire \thechain[4].chain7.inv_chain[94] ;
 wire \thechain[4].chain7.inv_chain[95] ;
 wire \thechain[4].chain7.inv_chain[96] ;
 wire \thechain[4].chain7.inv_chain[97] ;
 wire \thechain[4].chain7.inv_chain[98] ;
 wire \thechain[4].chain7.inv_chain[99] ;
 wire \thechain[4].chain7.inv_chain[9] ;
 wire \thechain[4].chain8.dout ;
 wire \thechain[4].chain8.inv_chain[0] ;
 wire \thechain[4].chain8.inv_chain[100] ;
 wire \thechain[4].chain8.inv_chain[101] ;
 wire \thechain[4].chain8.inv_chain[102] ;
 wire \thechain[4].chain8.inv_chain[103] ;
 wire \thechain[4].chain8.inv_chain[104] ;
 wire \thechain[4].chain8.inv_chain[105] ;
 wire \thechain[4].chain8.inv_chain[106] ;
 wire \thechain[4].chain8.inv_chain[107] ;
 wire \thechain[4].chain8.inv_chain[108] ;
 wire \thechain[4].chain8.inv_chain[109] ;
 wire \thechain[4].chain8.inv_chain[10] ;
 wire \thechain[4].chain8.inv_chain[110] ;
 wire \thechain[4].chain8.inv_chain[111] ;
 wire \thechain[4].chain8.inv_chain[112] ;
 wire \thechain[4].chain8.inv_chain[113] ;
 wire \thechain[4].chain8.inv_chain[114] ;
 wire \thechain[4].chain8.inv_chain[115] ;
 wire \thechain[4].chain8.inv_chain[116] ;
 wire \thechain[4].chain8.inv_chain[117] ;
 wire \thechain[4].chain8.inv_chain[118] ;
 wire \thechain[4].chain8.inv_chain[119] ;
 wire \thechain[4].chain8.inv_chain[11] ;
 wire \thechain[4].chain8.inv_chain[120] ;
 wire \thechain[4].chain8.inv_chain[121] ;
 wire \thechain[4].chain8.inv_chain[122] ;
 wire \thechain[4].chain8.inv_chain[123] ;
 wire \thechain[4].chain8.inv_chain[124] ;
 wire \thechain[4].chain8.inv_chain[125] ;
 wire \thechain[4].chain8.inv_chain[126] ;
 wire \thechain[4].chain8.inv_chain[127] ;
 wire \thechain[4].chain8.inv_chain[128] ;
 wire \thechain[4].chain8.inv_chain[129] ;
 wire \thechain[4].chain8.inv_chain[12] ;
 wire \thechain[4].chain8.inv_chain[130] ;
 wire \thechain[4].chain8.inv_chain[131] ;
 wire \thechain[4].chain8.inv_chain[132] ;
 wire \thechain[4].chain8.inv_chain[133] ;
 wire \thechain[4].chain8.inv_chain[134] ;
 wire \thechain[4].chain8.inv_chain[135] ;
 wire \thechain[4].chain8.inv_chain[136] ;
 wire \thechain[4].chain8.inv_chain[137] ;
 wire \thechain[4].chain8.inv_chain[138] ;
 wire \thechain[4].chain8.inv_chain[139] ;
 wire \thechain[4].chain8.inv_chain[13] ;
 wire \thechain[4].chain8.inv_chain[140] ;
 wire \thechain[4].chain8.inv_chain[141] ;
 wire \thechain[4].chain8.inv_chain[142] ;
 wire \thechain[4].chain8.inv_chain[143] ;
 wire \thechain[4].chain8.inv_chain[144] ;
 wire \thechain[4].chain8.inv_chain[145] ;
 wire \thechain[4].chain8.inv_chain[146] ;
 wire \thechain[4].chain8.inv_chain[147] ;
 wire \thechain[4].chain8.inv_chain[148] ;
 wire \thechain[4].chain8.inv_chain[149] ;
 wire \thechain[4].chain8.inv_chain[14] ;
 wire \thechain[4].chain8.inv_chain[150] ;
 wire \thechain[4].chain8.inv_chain[151] ;
 wire \thechain[4].chain8.inv_chain[152] ;
 wire \thechain[4].chain8.inv_chain[153] ;
 wire \thechain[4].chain8.inv_chain[154] ;
 wire \thechain[4].chain8.inv_chain[155] ;
 wire \thechain[4].chain8.inv_chain[156] ;
 wire \thechain[4].chain8.inv_chain[157] ;
 wire \thechain[4].chain8.inv_chain[158] ;
 wire \thechain[4].chain8.inv_chain[159] ;
 wire \thechain[4].chain8.inv_chain[15] ;
 wire \thechain[4].chain8.inv_chain[160] ;
 wire \thechain[4].chain8.inv_chain[161] ;
 wire \thechain[4].chain8.inv_chain[162] ;
 wire \thechain[4].chain8.inv_chain[163] ;
 wire \thechain[4].chain8.inv_chain[164] ;
 wire \thechain[4].chain8.inv_chain[165] ;
 wire \thechain[4].chain8.inv_chain[166] ;
 wire \thechain[4].chain8.inv_chain[167] ;
 wire \thechain[4].chain8.inv_chain[168] ;
 wire \thechain[4].chain8.inv_chain[169] ;
 wire \thechain[4].chain8.inv_chain[16] ;
 wire \thechain[4].chain8.inv_chain[170] ;
 wire \thechain[4].chain8.inv_chain[171] ;
 wire \thechain[4].chain8.inv_chain[172] ;
 wire \thechain[4].chain8.inv_chain[173] ;
 wire \thechain[4].chain8.inv_chain[174] ;
 wire \thechain[4].chain8.inv_chain[175] ;
 wire \thechain[4].chain8.inv_chain[176] ;
 wire \thechain[4].chain8.inv_chain[177] ;
 wire \thechain[4].chain8.inv_chain[178] ;
 wire \thechain[4].chain8.inv_chain[179] ;
 wire \thechain[4].chain8.inv_chain[17] ;
 wire \thechain[4].chain8.inv_chain[180] ;
 wire \thechain[4].chain8.inv_chain[181] ;
 wire \thechain[4].chain8.inv_chain[182] ;
 wire \thechain[4].chain8.inv_chain[183] ;
 wire \thechain[4].chain8.inv_chain[184] ;
 wire \thechain[4].chain8.inv_chain[185] ;
 wire \thechain[4].chain8.inv_chain[186] ;
 wire \thechain[4].chain8.inv_chain[187] ;
 wire \thechain[4].chain8.inv_chain[188] ;
 wire \thechain[4].chain8.inv_chain[189] ;
 wire \thechain[4].chain8.inv_chain[18] ;
 wire \thechain[4].chain8.inv_chain[190] ;
 wire \thechain[4].chain8.inv_chain[191] ;
 wire \thechain[4].chain8.inv_chain[192] ;
 wire \thechain[4].chain8.inv_chain[19] ;
 wire \thechain[4].chain8.inv_chain[1] ;
 wire \thechain[4].chain8.inv_chain[20] ;
 wire \thechain[4].chain8.inv_chain[21] ;
 wire \thechain[4].chain8.inv_chain[22] ;
 wire \thechain[4].chain8.inv_chain[23] ;
 wire \thechain[4].chain8.inv_chain[24] ;
 wire \thechain[4].chain8.inv_chain[25] ;
 wire \thechain[4].chain8.inv_chain[26] ;
 wire \thechain[4].chain8.inv_chain[27] ;
 wire \thechain[4].chain8.inv_chain[28] ;
 wire \thechain[4].chain8.inv_chain[29] ;
 wire \thechain[4].chain8.inv_chain[2] ;
 wire \thechain[4].chain8.inv_chain[30] ;
 wire \thechain[4].chain8.inv_chain[31] ;
 wire \thechain[4].chain8.inv_chain[32] ;
 wire \thechain[4].chain8.inv_chain[33] ;
 wire \thechain[4].chain8.inv_chain[34] ;
 wire \thechain[4].chain8.inv_chain[35] ;
 wire \thechain[4].chain8.inv_chain[36] ;
 wire \thechain[4].chain8.inv_chain[37] ;
 wire \thechain[4].chain8.inv_chain[38] ;
 wire \thechain[4].chain8.inv_chain[39] ;
 wire \thechain[4].chain8.inv_chain[3] ;
 wire \thechain[4].chain8.inv_chain[40] ;
 wire \thechain[4].chain8.inv_chain[41] ;
 wire \thechain[4].chain8.inv_chain[42] ;
 wire \thechain[4].chain8.inv_chain[43] ;
 wire \thechain[4].chain8.inv_chain[44] ;
 wire \thechain[4].chain8.inv_chain[45] ;
 wire \thechain[4].chain8.inv_chain[46] ;
 wire \thechain[4].chain8.inv_chain[47] ;
 wire \thechain[4].chain8.inv_chain[48] ;
 wire \thechain[4].chain8.inv_chain[49] ;
 wire \thechain[4].chain8.inv_chain[4] ;
 wire \thechain[4].chain8.inv_chain[50] ;
 wire \thechain[4].chain8.inv_chain[51] ;
 wire \thechain[4].chain8.inv_chain[52] ;
 wire \thechain[4].chain8.inv_chain[53] ;
 wire \thechain[4].chain8.inv_chain[54] ;
 wire \thechain[4].chain8.inv_chain[55] ;
 wire \thechain[4].chain8.inv_chain[56] ;
 wire \thechain[4].chain8.inv_chain[57] ;
 wire \thechain[4].chain8.inv_chain[58] ;
 wire \thechain[4].chain8.inv_chain[59] ;
 wire \thechain[4].chain8.inv_chain[5] ;
 wire \thechain[4].chain8.inv_chain[60] ;
 wire \thechain[4].chain8.inv_chain[61] ;
 wire \thechain[4].chain8.inv_chain[62] ;
 wire \thechain[4].chain8.inv_chain[63] ;
 wire \thechain[4].chain8.inv_chain[64] ;
 wire \thechain[4].chain8.inv_chain[65] ;
 wire \thechain[4].chain8.inv_chain[66] ;
 wire \thechain[4].chain8.inv_chain[67] ;
 wire \thechain[4].chain8.inv_chain[68] ;
 wire \thechain[4].chain8.inv_chain[69] ;
 wire \thechain[4].chain8.inv_chain[6] ;
 wire \thechain[4].chain8.inv_chain[70] ;
 wire \thechain[4].chain8.inv_chain[71] ;
 wire \thechain[4].chain8.inv_chain[72] ;
 wire \thechain[4].chain8.inv_chain[73] ;
 wire \thechain[4].chain8.inv_chain[74] ;
 wire \thechain[4].chain8.inv_chain[75] ;
 wire \thechain[4].chain8.inv_chain[76] ;
 wire \thechain[4].chain8.inv_chain[77] ;
 wire \thechain[4].chain8.inv_chain[78] ;
 wire \thechain[4].chain8.inv_chain[79] ;
 wire \thechain[4].chain8.inv_chain[7] ;
 wire \thechain[4].chain8.inv_chain[80] ;
 wire \thechain[4].chain8.inv_chain[81] ;
 wire \thechain[4].chain8.inv_chain[82] ;
 wire \thechain[4].chain8.inv_chain[83] ;
 wire \thechain[4].chain8.inv_chain[84] ;
 wire \thechain[4].chain8.inv_chain[85] ;
 wire \thechain[4].chain8.inv_chain[86] ;
 wire \thechain[4].chain8.inv_chain[87] ;
 wire \thechain[4].chain8.inv_chain[88] ;
 wire \thechain[4].chain8.inv_chain[89] ;
 wire \thechain[4].chain8.inv_chain[8] ;
 wire \thechain[4].chain8.inv_chain[90] ;
 wire \thechain[4].chain8.inv_chain[91] ;
 wire \thechain[4].chain8.inv_chain[92] ;
 wire \thechain[4].chain8.inv_chain[93] ;
 wire \thechain[4].chain8.inv_chain[94] ;
 wire \thechain[4].chain8.inv_chain[95] ;
 wire \thechain[4].chain8.inv_chain[96] ;
 wire \thechain[4].chain8.inv_chain[97] ;
 wire \thechain[4].chain8.inv_chain[98] ;
 wire \thechain[4].chain8.inv_chain[99] ;
 wire \thechain[4].chain8.inv_chain[9] ;
 wire \thechain[4].chain9.dout ;
 wire \thechain[4].chain9.inv_chain[0] ;
 wire \thechain[4].chain9.inv_chain[100] ;
 wire \thechain[4].chain9.inv_chain[101] ;
 wire \thechain[4].chain9.inv_chain[102] ;
 wire \thechain[4].chain9.inv_chain[103] ;
 wire \thechain[4].chain9.inv_chain[104] ;
 wire \thechain[4].chain9.inv_chain[105] ;
 wire \thechain[4].chain9.inv_chain[106] ;
 wire \thechain[4].chain9.inv_chain[107] ;
 wire \thechain[4].chain9.inv_chain[108] ;
 wire \thechain[4].chain9.inv_chain[109] ;
 wire \thechain[4].chain9.inv_chain[10] ;
 wire \thechain[4].chain9.inv_chain[110] ;
 wire \thechain[4].chain9.inv_chain[111] ;
 wire \thechain[4].chain9.inv_chain[112] ;
 wire \thechain[4].chain9.inv_chain[113] ;
 wire \thechain[4].chain9.inv_chain[114] ;
 wire \thechain[4].chain9.inv_chain[115] ;
 wire \thechain[4].chain9.inv_chain[116] ;
 wire \thechain[4].chain9.inv_chain[117] ;
 wire \thechain[4].chain9.inv_chain[118] ;
 wire \thechain[4].chain9.inv_chain[119] ;
 wire \thechain[4].chain9.inv_chain[11] ;
 wire \thechain[4].chain9.inv_chain[120] ;
 wire \thechain[4].chain9.inv_chain[121] ;
 wire \thechain[4].chain9.inv_chain[122] ;
 wire \thechain[4].chain9.inv_chain[123] ;
 wire \thechain[4].chain9.inv_chain[124] ;
 wire \thechain[4].chain9.inv_chain[125] ;
 wire \thechain[4].chain9.inv_chain[126] ;
 wire \thechain[4].chain9.inv_chain[127] ;
 wire \thechain[4].chain9.inv_chain[128] ;
 wire \thechain[4].chain9.inv_chain[129] ;
 wire \thechain[4].chain9.inv_chain[12] ;
 wire \thechain[4].chain9.inv_chain[130] ;
 wire \thechain[4].chain9.inv_chain[131] ;
 wire \thechain[4].chain9.inv_chain[132] ;
 wire \thechain[4].chain9.inv_chain[133] ;
 wire \thechain[4].chain9.inv_chain[134] ;
 wire \thechain[4].chain9.inv_chain[135] ;
 wire \thechain[4].chain9.inv_chain[136] ;
 wire \thechain[4].chain9.inv_chain[137] ;
 wire \thechain[4].chain9.inv_chain[138] ;
 wire \thechain[4].chain9.inv_chain[139] ;
 wire \thechain[4].chain9.inv_chain[13] ;
 wire \thechain[4].chain9.inv_chain[140] ;
 wire \thechain[4].chain9.inv_chain[141] ;
 wire \thechain[4].chain9.inv_chain[142] ;
 wire \thechain[4].chain9.inv_chain[143] ;
 wire \thechain[4].chain9.inv_chain[144] ;
 wire \thechain[4].chain9.inv_chain[145] ;
 wire \thechain[4].chain9.inv_chain[146] ;
 wire \thechain[4].chain9.inv_chain[147] ;
 wire \thechain[4].chain9.inv_chain[148] ;
 wire \thechain[4].chain9.inv_chain[149] ;
 wire \thechain[4].chain9.inv_chain[14] ;
 wire \thechain[4].chain9.inv_chain[150] ;
 wire \thechain[4].chain9.inv_chain[151] ;
 wire \thechain[4].chain9.inv_chain[152] ;
 wire \thechain[4].chain9.inv_chain[153] ;
 wire \thechain[4].chain9.inv_chain[154] ;
 wire \thechain[4].chain9.inv_chain[155] ;
 wire \thechain[4].chain9.inv_chain[156] ;
 wire \thechain[4].chain9.inv_chain[157] ;
 wire \thechain[4].chain9.inv_chain[158] ;
 wire \thechain[4].chain9.inv_chain[159] ;
 wire \thechain[4].chain9.inv_chain[15] ;
 wire \thechain[4].chain9.inv_chain[160] ;
 wire \thechain[4].chain9.inv_chain[161] ;
 wire \thechain[4].chain9.inv_chain[162] ;
 wire \thechain[4].chain9.inv_chain[163] ;
 wire \thechain[4].chain9.inv_chain[164] ;
 wire \thechain[4].chain9.inv_chain[165] ;
 wire \thechain[4].chain9.inv_chain[166] ;
 wire \thechain[4].chain9.inv_chain[167] ;
 wire \thechain[4].chain9.inv_chain[168] ;
 wire \thechain[4].chain9.inv_chain[169] ;
 wire \thechain[4].chain9.inv_chain[16] ;
 wire \thechain[4].chain9.inv_chain[170] ;
 wire \thechain[4].chain9.inv_chain[171] ;
 wire \thechain[4].chain9.inv_chain[172] ;
 wire \thechain[4].chain9.inv_chain[173] ;
 wire \thechain[4].chain9.inv_chain[174] ;
 wire \thechain[4].chain9.inv_chain[175] ;
 wire \thechain[4].chain9.inv_chain[176] ;
 wire \thechain[4].chain9.inv_chain[177] ;
 wire \thechain[4].chain9.inv_chain[178] ;
 wire \thechain[4].chain9.inv_chain[179] ;
 wire \thechain[4].chain9.inv_chain[17] ;
 wire \thechain[4].chain9.inv_chain[180] ;
 wire \thechain[4].chain9.inv_chain[181] ;
 wire \thechain[4].chain9.inv_chain[182] ;
 wire \thechain[4].chain9.inv_chain[183] ;
 wire \thechain[4].chain9.inv_chain[184] ;
 wire \thechain[4].chain9.inv_chain[185] ;
 wire \thechain[4].chain9.inv_chain[186] ;
 wire \thechain[4].chain9.inv_chain[187] ;
 wire \thechain[4].chain9.inv_chain[188] ;
 wire \thechain[4].chain9.inv_chain[189] ;
 wire \thechain[4].chain9.inv_chain[18] ;
 wire \thechain[4].chain9.inv_chain[190] ;
 wire \thechain[4].chain9.inv_chain[191] ;
 wire \thechain[4].chain9.inv_chain[192] ;
 wire \thechain[4].chain9.inv_chain[193] ;
 wire \thechain[4].chain9.inv_chain[194] ;
 wire \thechain[4].chain9.inv_chain[195] ;
 wire \thechain[4].chain9.inv_chain[196] ;
 wire \thechain[4].chain9.inv_chain[197] ;
 wire \thechain[4].chain9.inv_chain[198] ;
 wire \thechain[4].chain9.inv_chain[199] ;
 wire \thechain[4].chain9.inv_chain[19] ;
 wire \thechain[4].chain9.inv_chain[1] ;
 wire \thechain[4].chain9.inv_chain[200] ;
 wire \thechain[4].chain9.inv_chain[201] ;
 wire \thechain[4].chain9.inv_chain[202] ;
 wire \thechain[4].chain9.inv_chain[203] ;
 wire \thechain[4].chain9.inv_chain[204] ;
 wire \thechain[4].chain9.inv_chain[205] ;
 wire \thechain[4].chain9.inv_chain[206] ;
 wire \thechain[4].chain9.inv_chain[207] ;
 wire \thechain[4].chain9.inv_chain[208] ;
 wire \thechain[4].chain9.inv_chain[209] ;
 wire \thechain[4].chain9.inv_chain[20] ;
 wire \thechain[4].chain9.inv_chain[210] ;
 wire \thechain[4].chain9.inv_chain[211] ;
 wire \thechain[4].chain9.inv_chain[212] ;
 wire \thechain[4].chain9.inv_chain[213] ;
 wire \thechain[4].chain9.inv_chain[214] ;
 wire \thechain[4].chain9.inv_chain[215] ;
 wire \thechain[4].chain9.inv_chain[216] ;
 wire \thechain[4].chain9.inv_chain[217] ;
 wire \thechain[4].chain9.inv_chain[218] ;
 wire \thechain[4].chain9.inv_chain[219] ;
 wire \thechain[4].chain9.inv_chain[21] ;
 wire \thechain[4].chain9.inv_chain[220] ;
 wire \thechain[4].chain9.inv_chain[221] ;
 wire \thechain[4].chain9.inv_chain[222] ;
 wire \thechain[4].chain9.inv_chain[223] ;
 wire \thechain[4].chain9.inv_chain[224] ;
 wire \thechain[4].chain9.inv_chain[225] ;
 wire \thechain[4].chain9.inv_chain[226] ;
 wire \thechain[4].chain9.inv_chain[227] ;
 wire \thechain[4].chain9.inv_chain[228] ;
 wire \thechain[4].chain9.inv_chain[229] ;
 wire \thechain[4].chain9.inv_chain[22] ;
 wire \thechain[4].chain9.inv_chain[230] ;
 wire \thechain[4].chain9.inv_chain[231] ;
 wire \thechain[4].chain9.inv_chain[232] ;
 wire \thechain[4].chain9.inv_chain[233] ;
 wire \thechain[4].chain9.inv_chain[234] ;
 wire \thechain[4].chain9.inv_chain[235] ;
 wire \thechain[4].chain9.inv_chain[236] ;
 wire \thechain[4].chain9.inv_chain[237] ;
 wire \thechain[4].chain9.inv_chain[238] ;
 wire \thechain[4].chain9.inv_chain[239] ;
 wire \thechain[4].chain9.inv_chain[23] ;
 wire \thechain[4].chain9.inv_chain[240] ;
 wire \thechain[4].chain9.inv_chain[241] ;
 wire \thechain[4].chain9.inv_chain[242] ;
 wire \thechain[4].chain9.inv_chain[243] ;
 wire \thechain[4].chain9.inv_chain[244] ;
 wire \thechain[4].chain9.inv_chain[245] ;
 wire \thechain[4].chain9.inv_chain[246] ;
 wire \thechain[4].chain9.inv_chain[247] ;
 wire \thechain[4].chain9.inv_chain[248] ;
 wire \thechain[4].chain9.inv_chain[249] ;
 wire \thechain[4].chain9.inv_chain[24] ;
 wire \thechain[4].chain9.inv_chain[250] ;
 wire \thechain[4].chain9.inv_chain[251] ;
 wire \thechain[4].chain9.inv_chain[252] ;
 wire \thechain[4].chain9.inv_chain[253] ;
 wire \thechain[4].chain9.inv_chain[254] ;
 wire \thechain[4].chain9.inv_chain[255] ;
 wire \thechain[4].chain9.inv_chain[256] ;
 wire \thechain[4].chain9.inv_chain[25] ;
 wire \thechain[4].chain9.inv_chain[26] ;
 wire \thechain[4].chain9.inv_chain[27] ;
 wire \thechain[4].chain9.inv_chain[28] ;
 wire \thechain[4].chain9.inv_chain[29] ;
 wire \thechain[4].chain9.inv_chain[2] ;
 wire \thechain[4].chain9.inv_chain[30] ;
 wire \thechain[4].chain9.inv_chain[31] ;
 wire \thechain[4].chain9.inv_chain[32] ;
 wire \thechain[4].chain9.inv_chain[33] ;
 wire \thechain[4].chain9.inv_chain[34] ;
 wire \thechain[4].chain9.inv_chain[35] ;
 wire \thechain[4].chain9.inv_chain[36] ;
 wire \thechain[4].chain9.inv_chain[37] ;
 wire \thechain[4].chain9.inv_chain[38] ;
 wire \thechain[4].chain9.inv_chain[39] ;
 wire \thechain[4].chain9.inv_chain[3] ;
 wire \thechain[4].chain9.inv_chain[40] ;
 wire \thechain[4].chain9.inv_chain[41] ;
 wire \thechain[4].chain9.inv_chain[42] ;
 wire \thechain[4].chain9.inv_chain[43] ;
 wire \thechain[4].chain9.inv_chain[44] ;
 wire \thechain[4].chain9.inv_chain[45] ;
 wire \thechain[4].chain9.inv_chain[46] ;
 wire \thechain[4].chain9.inv_chain[47] ;
 wire \thechain[4].chain9.inv_chain[48] ;
 wire \thechain[4].chain9.inv_chain[49] ;
 wire \thechain[4].chain9.inv_chain[4] ;
 wire \thechain[4].chain9.inv_chain[50] ;
 wire \thechain[4].chain9.inv_chain[51] ;
 wire \thechain[4].chain9.inv_chain[52] ;
 wire \thechain[4].chain9.inv_chain[53] ;
 wire \thechain[4].chain9.inv_chain[54] ;
 wire \thechain[4].chain9.inv_chain[55] ;
 wire \thechain[4].chain9.inv_chain[56] ;
 wire \thechain[4].chain9.inv_chain[57] ;
 wire \thechain[4].chain9.inv_chain[58] ;
 wire \thechain[4].chain9.inv_chain[59] ;
 wire \thechain[4].chain9.inv_chain[5] ;
 wire \thechain[4].chain9.inv_chain[60] ;
 wire \thechain[4].chain9.inv_chain[61] ;
 wire \thechain[4].chain9.inv_chain[62] ;
 wire \thechain[4].chain9.inv_chain[63] ;
 wire \thechain[4].chain9.inv_chain[64] ;
 wire \thechain[4].chain9.inv_chain[65] ;
 wire \thechain[4].chain9.inv_chain[66] ;
 wire \thechain[4].chain9.inv_chain[67] ;
 wire \thechain[4].chain9.inv_chain[68] ;
 wire \thechain[4].chain9.inv_chain[69] ;
 wire \thechain[4].chain9.inv_chain[6] ;
 wire \thechain[4].chain9.inv_chain[70] ;
 wire \thechain[4].chain9.inv_chain[71] ;
 wire \thechain[4].chain9.inv_chain[72] ;
 wire \thechain[4].chain9.inv_chain[73] ;
 wire \thechain[4].chain9.inv_chain[74] ;
 wire \thechain[4].chain9.inv_chain[75] ;
 wire \thechain[4].chain9.inv_chain[76] ;
 wire \thechain[4].chain9.inv_chain[77] ;
 wire \thechain[4].chain9.inv_chain[78] ;
 wire \thechain[4].chain9.inv_chain[79] ;
 wire \thechain[4].chain9.inv_chain[7] ;
 wire \thechain[4].chain9.inv_chain[80] ;
 wire \thechain[4].chain9.inv_chain[81] ;
 wire \thechain[4].chain9.inv_chain[82] ;
 wire \thechain[4].chain9.inv_chain[83] ;
 wire \thechain[4].chain9.inv_chain[84] ;
 wire \thechain[4].chain9.inv_chain[85] ;
 wire \thechain[4].chain9.inv_chain[86] ;
 wire \thechain[4].chain9.inv_chain[87] ;
 wire \thechain[4].chain9.inv_chain[88] ;
 wire \thechain[4].chain9.inv_chain[89] ;
 wire \thechain[4].chain9.inv_chain[8] ;
 wire \thechain[4].chain9.inv_chain[90] ;
 wire \thechain[4].chain9.inv_chain[91] ;
 wire \thechain[4].chain9.inv_chain[92] ;
 wire \thechain[4].chain9.inv_chain[93] ;
 wire \thechain[4].chain9.inv_chain[94] ;
 wire \thechain[4].chain9.inv_chain[95] ;
 wire \thechain[4].chain9.inv_chain[96] ;
 wire \thechain[4].chain9.inv_chain[97] ;
 wire \thechain[4].chain9.inv_chain[98] ;
 wire \thechain[4].chain9.inv_chain[99] ;
 wire \thechain[4].chain9.inv_chain[9] ;
 wire \thechain[5].chain1.dout ;
 wire \thechain[5].chain1.inv_chain[0] ;
 wire \thechain[5].chain1.inv_chain[1] ;
 wire \thechain[5].chain1.inv_chain[2] ;
 wire \thechain[5].chain2.dout ;
 wire \thechain[5].chain2.inv_chain[0] ;
 wire \thechain[5].chain2.inv_chain[1] ;
 wire \thechain[5].chain2.inv_chain[2] ;
 wire \thechain[5].chain2.inv_chain[3] ;
 wire \thechain[5].chain2.inv_chain[4] ;
 wire \thechain[5].chain3.dout ;
 wire \thechain[5].chain3.inv_chain[0] ;
 wire \thechain[5].chain3.inv_chain[1] ;
 wire \thechain[5].chain3.inv_chain[2] ;
 wire \thechain[5].chain3.inv_chain[3] ;
 wire \thechain[5].chain3.inv_chain[4] ;
 wire \thechain[5].chain3.inv_chain[5] ;
 wire \thechain[5].chain3.inv_chain[6] ;
 wire \thechain[5].chain3.inv_chain[7] ;
 wire \thechain[5].chain3.inv_chain[8] ;
 wire \thechain[5].chain4.dout ;
 wire \thechain[5].chain4.inv_chain[0] ;
 wire \thechain[5].chain4.inv_chain[10] ;
 wire \thechain[5].chain4.inv_chain[11] ;
 wire \thechain[5].chain4.inv_chain[12] ;
 wire \thechain[5].chain4.inv_chain[13] ;
 wire \thechain[5].chain4.inv_chain[14] ;
 wire \thechain[5].chain4.inv_chain[15] ;
 wire \thechain[5].chain4.inv_chain[16] ;
 wire \thechain[5].chain4.inv_chain[1] ;
 wire \thechain[5].chain4.inv_chain[2] ;
 wire \thechain[5].chain4.inv_chain[3] ;
 wire \thechain[5].chain4.inv_chain[4] ;
 wire \thechain[5].chain4.inv_chain[5] ;
 wire \thechain[5].chain4.inv_chain[6] ;
 wire \thechain[5].chain4.inv_chain[7] ;
 wire \thechain[5].chain4.inv_chain[8] ;
 wire \thechain[5].chain4.inv_chain[9] ;
 wire \thechain[5].chain5.dout ;
 wire \thechain[5].chain5.inv_chain[0] ;
 wire \thechain[5].chain5.inv_chain[10] ;
 wire \thechain[5].chain5.inv_chain[11] ;
 wire \thechain[5].chain5.inv_chain[12] ;
 wire \thechain[5].chain5.inv_chain[13] ;
 wire \thechain[5].chain5.inv_chain[14] ;
 wire \thechain[5].chain5.inv_chain[15] ;
 wire \thechain[5].chain5.inv_chain[16] ;
 wire \thechain[5].chain5.inv_chain[17] ;
 wire \thechain[5].chain5.inv_chain[18] ;
 wire \thechain[5].chain5.inv_chain[19] ;
 wire \thechain[5].chain5.inv_chain[1] ;
 wire \thechain[5].chain5.inv_chain[20] ;
 wire \thechain[5].chain5.inv_chain[21] ;
 wire \thechain[5].chain5.inv_chain[22] ;
 wire \thechain[5].chain5.inv_chain[23] ;
 wire \thechain[5].chain5.inv_chain[24] ;
 wire \thechain[5].chain5.inv_chain[25] ;
 wire \thechain[5].chain5.inv_chain[26] ;
 wire \thechain[5].chain5.inv_chain[27] ;
 wire \thechain[5].chain5.inv_chain[28] ;
 wire \thechain[5].chain5.inv_chain[29] ;
 wire \thechain[5].chain5.inv_chain[2] ;
 wire \thechain[5].chain5.inv_chain[30] ;
 wire \thechain[5].chain5.inv_chain[31] ;
 wire \thechain[5].chain5.inv_chain[32] ;
 wire \thechain[5].chain5.inv_chain[3] ;
 wire \thechain[5].chain5.inv_chain[4] ;
 wire \thechain[5].chain5.inv_chain[5] ;
 wire \thechain[5].chain5.inv_chain[6] ;
 wire \thechain[5].chain5.inv_chain[7] ;
 wire \thechain[5].chain5.inv_chain[8] ;
 wire \thechain[5].chain5.inv_chain[9] ;
 wire \thechain[5].chain6.dout ;
 wire \thechain[5].chain6.inv_chain[0] ;
 wire \thechain[5].chain6.inv_chain[10] ;
 wire \thechain[5].chain6.inv_chain[11] ;
 wire \thechain[5].chain6.inv_chain[12] ;
 wire \thechain[5].chain6.inv_chain[13] ;
 wire \thechain[5].chain6.inv_chain[14] ;
 wire \thechain[5].chain6.inv_chain[15] ;
 wire \thechain[5].chain6.inv_chain[16] ;
 wire \thechain[5].chain6.inv_chain[17] ;
 wire \thechain[5].chain6.inv_chain[18] ;
 wire \thechain[5].chain6.inv_chain[19] ;
 wire \thechain[5].chain6.inv_chain[1] ;
 wire \thechain[5].chain6.inv_chain[20] ;
 wire \thechain[5].chain6.inv_chain[21] ;
 wire \thechain[5].chain6.inv_chain[22] ;
 wire \thechain[5].chain6.inv_chain[23] ;
 wire \thechain[5].chain6.inv_chain[24] ;
 wire \thechain[5].chain6.inv_chain[25] ;
 wire \thechain[5].chain6.inv_chain[26] ;
 wire \thechain[5].chain6.inv_chain[27] ;
 wire \thechain[5].chain6.inv_chain[28] ;
 wire \thechain[5].chain6.inv_chain[29] ;
 wire \thechain[5].chain6.inv_chain[2] ;
 wire \thechain[5].chain6.inv_chain[30] ;
 wire \thechain[5].chain6.inv_chain[31] ;
 wire \thechain[5].chain6.inv_chain[32] ;
 wire \thechain[5].chain6.inv_chain[33] ;
 wire \thechain[5].chain6.inv_chain[34] ;
 wire \thechain[5].chain6.inv_chain[35] ;
 wire \thechain[5].chain6.inv_chain[36] ;
 wire \thechain[5].chain6.inv_chain[37] ;
 wire \thechain[5].chain6.inv_chain[38] ;
 wire \thechain[5].chain6.inv_chain[39] ;
 wire \thechain[5].chain6.inv_chain[3] ;
 wire \thechain[5].chain6.inv_chain[40] ;
 wire \thechain[5].chain6.inv_chain[41] ;
 wire \thechain[5].chain6.inv_chain[42] ;
 wire \thechain[5].chain6.inv_chain[43] ;
 wire \thechain[5].chain6.inv_chain[44] ;
 wire \thechain[5].chain6.inv_chain[45] ;
 wire \thechain[5].chain6.inv_chain[46] ;
 wire \thechain[5].chain6.inv_chain[47] ;
 wire \thechain[5].chain6.inv_chain[48] ;
 wire \thechain[5].chain6.inv_chain[49] ;
 wire \thechain[5].chain6.inv_chain[4] ;
 wire \thechain[5].chain6.inv_chain[50] ;
 wire \thechain[5].chain6.inv_chain[51] ;
 wire \thechain[5].chain6.inv_chain[52] ;
 wire \thechain[5].chain6.inv_chain[53] ;
 wire \thechain[5].chain6.inv_chain[54] ;
 wire \thechain[5].chain6.inv_chain[55] ;
 wire \thechain[5].chain6.inv_chain[56] ;
 wire \thechain[5].chain6.inv_chain[57] ;
 wire \thechain[5].chain6.inv_chain[58] ;
 wire \thechain[5].chain6.inv_chain[59] ;
 wire \thechain[5].chain6.inv_chain[5] ;
 wire \thechain[5].chain6.inv_chain[60] ;
 wire \thechain[5].chain6.inv_chain[61] ;
 wire \thechain[5].chain6.inv_chain[62] ;
 wire \thechain[5].chain6.inv_chain[63] ;
 wire \thechain[5].chain6.inv_chain[64] ;
 wire \thechain[5].chain6.inv_chain[6] ;
 wire \thechain[5].chain6.inv_chain[7] ;
 wire \thechain[5].chain6.inv_chain[8] ;
 wire \thechain[5].chain6.inv_chain[9] ;
 wire \thechain[5].chain7.dout ;
 wire \thechain[5].chain7.inv_chain[0] ;
 wire \thechain[5].chain7.inv_chain[100] ;
 wire \thechain[5].chain7.inv_chain[101] ;
 wire \thechain[5].chain7.inv_chain[102] ;
 wire \thechain[5].chain7.inv_chain[103] ;
 wire \thechain[5].chain7.inv_chain[104] ;
 wire \thechain[5].chain7.inv_chain[105] ;
 wire \thechain[5].chain7.inv_chain[106] ;
 wire \thechain[5].chain7.inv_chain[107] ;
 wire \thechain[5].chain7.inv_chain[108] ;
 wire \thechain[5].chain7.inv_chain[109] ;
 wire \thechain[5].chain7.inv_chain[10] ;
 wire \thechain[5].chain7.inv_chain[110] ;
 wire \thechain[5].chain7.inv_chain[111] ;
 wire \thechain[5].chain7.inv_chain[112] ;
 wire \thechain[5].chain7.inv_chain[113] ;
 wire \thechain[5].chain7.inv_chain[114] ;
 wire \thechain[5].chain7.inv_chain[115] ;
 wire \thechain[5].chain7.inv_chain[116] ;
 wire \thechain[5].chain7.inv_chain[117] ;
 wire \thechain[5].chain7.inv_chain[118] ;
 wire \thechain[5].chain7.inv_chain[119] ;
 wire \thechain[5].chain7.inv_chain[11] ;
 wire \thechain[5].chain7.inv_chain[120] ;
 wire \thechain[5].chain7.inv_chain[121] ;
 wire \thechain[5].chain7.inv_chain[122] ;
 wire \thechain[5].chain7.inv_chain[123] ;
 wire \thechain[5].chain7.inv_chain[124] ;
 wire \thechain[5].chain7.inv_chain[125] ;
 wire \thechain[5].chain7.inv_chain[126] ;
 wire \thechain[5].chain7.inv_chain[127] ;
 wire \thechain[5].chain7.inv_chain[128] ;
 wire \thechain[5].chain7.inv_chain[12] ;
 wire \thechain[5].chain7.inv_chain[13] ;
 wire \thechain[5].chain7.inv_chain[14] ;
 wire \thechain[5].chain7.inv_chain[15] ;
 wire \thechain[5].chain7.inv_chain[16] ;
 wire \thechain[5].chain7.inv_chain[17] ;
 wire \thechain[5].chain7.inv_chain[18] ;
 wire \thechain[5].chain7.inv_chain[19] ;
 wire \thechain[5].chain7.inv_chain[1] ;
 wire \thechain[5].chain7.inv_chain[20] ;
 wire \thechain[5].chain7.inv_chain[21] ;
 wire \thechain[5].chain7.inv_chain[22] ;
 wire \thechain[5].chain7.inv_chain[23] ;
 wire \thechain[5].chain7.inv_chain[24] ;
 wire \thechain[5].chain7.inv_chain[25] ;
 wire \thechain[5].chain7.inv_chain[26] ;
 wire \thechain[5].chain7.inv_chain[27] ;
 wire \thechain[5].chain7.inv_chain[28] ;
 wire \thechain[5].chain7.inv_chain[29] ;
 wire \thechain[5].chain7.inv_chain[2] ;
 wire \thechain[5].chain7.inv_chain[30] ;
 wire \thechain[5].chain7.inv_chain[31] ;
 wire \thechain[5].chain7.inv_chain[32] ;
 wire \thechain[5].chain7.inv_chain[33] ;
 wire \thechain[5].chain7.inv_chain[34] ;
 wire \thechain[5].chain7.inv_chain[35] ;
 wire \thechain[5].chain7.inv_chain[36] ;
 wire \thechain[5].chain7.inv_chain[37] ;
 wire \thechain[5].chain7.inv_chain[38] ;
 wire \thechain[5].chain7.inv_chain[39] ;
 wire \thechain[5].chain7.inv_chain[3] ;
 wire \thechain[5].chain7.inv_chain[40] ;
 wire \thechain[5].chain7.inv_chain[41] ;
 wire \thechain[5].chain7.inv_chain[42] ;
 wire \thechain[5].chain7.inv_chain[43] ;
 wire \thechain[5].chain7.inv_chain[44] ;
 wire \thechain[5].chain7.inv_chain[45] ;
 wire \thechain[5].chain7.inv_chain[46] ;
 wire \thechain[5].chain7.inv_chain[47] ;
 wire \thechain[5].chain7.inv_chain[48] ;
 wire \thechain[5].chain7.inv_chain[49] ;
 wire \thechain[5].chain7.inv_chain[4] ;
 wire \thechain[5].chain7.inv_chain[50] ;
 wire \thechain[5].chain7.inv_chain[51] ;
 wire \thechain[5].chain7.inv_chain[52] ;
 wire \thechain[5].chain7.inv_chain[53] ;
 wire \thechain[5].chain7.inv_chain[54] ;
 wire \thechain[5].chain7.inv_chain[55] ;
 wire \thechain[5].chain7.inv_chain[56] ;
 wire \thechain[5].chain7.inv_chain[57] ;
 wire \thechain[5].chain7.inv_chain[58] ;
 wire \thechain[5].chain7.inv_chain[59] ;
 wire \thechain[5].chain7.inv_chain[5] ;
 wire \thechain[5].chain7.inv_chain[60] ;
 wire \thechain[5].chain7.inv_chain[61] ;
 wire \thechain[5].chain7.inv_chain[62] ;
 wire \thechain[5].chain7.inv_chain[63] ;
 wire \thechain[5].chain7.inv_chain[64] ;
 wire \thechain[5].chain7.inv_chain[65] ;
 wire \thechain[5].chain7.inv_chain[66] ;
 wire \thechain[5].chain7.inv_chain[67] ;
 wire \thechain[5].chain7.inv_chain[68] ;
 wire \thechain[5].chain7.inv_chain[69] ;
 wire \thechain[5].chain7.inv_chain[6] ;
 wire \thechain[5].chain7.inv_chain[70] ;
 wire \thechain[5].chain7.inv_chain[71] ;
 wire \thechain[5].chain7.inv_chain[72] ;
 wire \thechain[5].chain7.inv_chain[73] ;
 wire \thechain[5].chain7.inv_chain[74] ;
 wire \thechain[5].chain7.inv_chain[75] ;
 wire \thechain[5].chain7.inv_chain[76] ;
 wire \thechain[5].chain7.inv_chain[77] ;
 wire \thechain[5].chain7.inv_chain[78] ;
 wire \thechain[5].chain7.inv_chain[79] ;
 wire \thechain[5].chain7.inv_chain[7] ;
 wire \thechain[5].chain7.inv_chain[80] ;
 wire \thechain[5].chain7.inv_chain[81] ;
 wire \thechain[5].chain7.inv_chain[82] ;
 wire \thechain[5].chain7.inv_chain[83] ;
 wire \thechain[5].chain7.inv_chain[84] ;
 wire \thechain[5].chain7.inv_chain[85] ;
 wire \thechain[5].chain7.inv_chain[86] ;
 wire \thechain[5].chain7.inv_chain[87] ;
 wire \thechain[5].chain7.inv_chain[88] ;
 wire \thechain[5].chain7.inv_chain[89] ;
 wire \thechain[5].chain7.inv_chain[8] ;
 wire \thechain[5].chain7.inv_chain[90] ;
 wire \thechain[5].chain7.inv_chain[91] ;
 wire \thechain[5].chain7.inv_chain[92] ;
 wire \thechain[5].chain7.inv_chain[93] ;
 wire \thechain[5].chain7.inv_chain[94] ;
 wire \thechain[5].chain7.inv_chain[95] ;
 wire \thechain[5].chain7.inv_chain[96] ;
 wire \thechain[5].chain7.inv_chain[97] ;
 wire \thechain[5].chain7.inv_chain[98] ;
 wire \thechain[5].chain7.inv_chain[99] ;
 wire \thechain[5].chain7.inv_chain[9] ;
 wire \thechain[5].chain8.dout ;
 wire \thechain[5].chain8.inv_chain[0] ;
 wire \thechain[5].chain8.inv_chain[100] ;
 wire \thechain[5].chain8.inv_chain[101] ;
 wire \thechain[5].chain8.inv_chain[102] ;
 wire \thechain[5].chain8.inv_chain[103] ;
 wire \thechain[5].chain8.inv_chain[104] ;
 wire \thechain[5].chain8.inv_chain[105] ;
 wire \thechain[5].chain8.inv_chain[106] ;
 wire \thechain[5].chain8.inv_chain[107] ;
 wire \thechain[5].chain8.inv_chain[108] ;
 wire \thechain[5].chain8.inv_chain[109] ;
 wire \thechain[5].chain8.inv_chain[10] ;
 wire \thechain[5].chain8.inv_chain[110] ;
 wire \thechain[5].chain8.inv_chain[111] ;
 wire \thechain[5].chain8.inv_chain[112] ;
 wire \thechain[5].chain8.inv_chain[113] ;
 wire \thechain[5].chain8.inv_chain[114] ;
 wire \thechain[5].chain8.inv_chain[115] ;
 wire \thechain[5].chain8.inv_chain[116] ;
 wire \thechain[5].chain8.inv_chain[117] ;
 wire \thechain[5].chain8.inv_chain[118] ;
 wire \thechain[5].chain8.inv_chain[119] ;
 wire \thechain[5].chain8.inv_chain[11] ;
 wire \thechain[5].chain8.inv_chain[120] ;
 wire \thechain[5].chain8.inv_chain[121] ;
 wire \thechain[5].chain8.inv_chain[122] ;
 wire \thechain[5].chain8.inv_chain[123] ;
 wire \thechain[5].chain8.inv_chain[124] ;
 wire \thechain[5].chain8.inv_chain[125] ;
 wire \thechain[5].chain8.inv_chain[126] ;
 wire \thechain[5].chain8.inv_chain[127] ;
 wire \thechain[5].chain8.inv_chain[128] ;
 wire \thechain[5].chain8.inv_chain[129] ;
 wire \thechain[5].chain8.inv_chain[12] ;
 wire \thechain[5].chain8.inv_chain[130] ;
 wire \thechain[5].chain8.inv_chain[131] ;
 wire \thechain[5].chain8.inv_chain[132] ;
 wire \thechain[5].chain8.inv_chain[133] ;
 wire \thechain[5].chain8.inv_chain[134] ;
 wire \thechain[5].chain8.inv_chain[135] ;
 wire \thechain[5].chain8.inv_chain[136] ;
 wire \thechain[5].chain8.inv_chain[137] ;
 wire \thechain[5].chain8.inv_chain[138] ;
 wire \thechain[5].chain8.inv_chain[139] ;
 wire \thechain[5].chain8.inv_chain[13] ;
 wire \thechain[5].chain8.inv_chain[140] ;
 wire \thechain[5].chain8.inv_chain[141] ;
 wire \thechain[5].chain8.inv_chain[142] ;
 wire \thechain[5].chain8.inv_chain[143] ;
 wire \thechain[5].chain8.inv_chain[144] ;
 wire \thechain[5].chain8.inv_chain[145] ;
 wire \thechain[5].chain8.inv_chain[146] ;
 wire \thechain[5].chain8.inv_chain[147] ;
 wire \thechain[5].chain8.inv_chain[148] ;
 wire \thechain[5].chain8.inv_chain[149] ;
 wire \thechain[5].chain8.inv_chain[14] ;
 wire \thechain[5].chain8.inv_chain[150] ;
 wire \thechain[5].chain8.inv_chain[151] ;
 wire \thechain[5].chain8.inv_chain[152] ;
 wire \thechain[5].chain8.inv_chain[153] ;
 wire \thechain[5].chain8.inv_chain[154] ;
 wire \thechain[5].chain8.inv_chain[155] ;
 wire \thechain[5].chain8.inv_chain[156] ;
 wire \thechain[5].chain8.inv_chain[157] ;
 wire \thechain[5].chain8.inv_chain[158] ;
 wire \thechain[5].chain8.inv_chain[159] ;
 wire \thechain[5].chain8.inv_chain[15] ;
 wire \thechain[5].chain8.inv_chain[160] ;
 wire \thechain[5].chain8.inv_chain[161] ;
 wire \thechain[5].chain8.inv_chain[162] ;
 wire \thechain[5].chain8.inv_chain[163] ;
 wire \thechain[5].chain8.inv_chain[164] ;
 wire \thechain[5].chain8.inv_chain[165] ;
 wire \thechain[5].chain8.inv_chain[166] ;
 wire \thechain[5].chain8.inv_chain[167] ;
 wire \thechain[5].chain8.inv_chain[168] ;
 wire \thechain[5].chain8.inv_chain[169] ;
 wire \thechain[5].chain8.inv_chain[16] ;
 wire \thechain[5].chain8.inv_chain[170] ;
 wire \thechain[5].chain8.inv_chain[171] ;
 wire \thechain[5].chain8.inv_chain[172] ;
 wire \thechain[5].chain8.inv_chain[173] ;
 wire \thechain[5].chain8.inv_chain[174] ;
 wire \thechain[5].chain8.inv_chain[175] ;
 wire \thechain[5].chain8.inv_chain[176] ;
 wire \thechain[5].chain8.inv_chain[177] ;
 wire \thechain[5].chain8.inv_chain[178] ;
 wire \thechain[5].chain8.inv_chain[179] ;
 wire \thechain[5].chain8.inv_chain[17] ;
 wire \thechain[5].chain8.inv_chain[180] ;
 wire \thechain[5].chain8.inv_chain[181] ;
 wire \thechain[5].chain8.inv_chain[182] ;
 wire \thechain[5].chain8.inv_chain[183] ;
 wire \thechain[5].chain8.inv_chain[184] ;
 wire \thechain[5].chain8.inv_chain[185] ;
 wire \thechain[5].chain8.inv_chain[186] ;
 wire \thechain[5].chain8.inv_chain[187] ;
 wire \thechain[5].chain8.inv_chain[188] ;
 wire \thechain[5].chain8.inv_chain[189] ;
 wire \thechain[5].chain8.inv_chain[18] ;
 wire \thechain[5].chain8.inv_chain[190] ;
 wire \thechain[5].chain8.inv_chain[191] ;
 wire \thechain[5].chain8.inv_chain[192] ;
 wire \thechain[5].chain8.inv_chain[19] ;
 wire \thechain[5].chain8.inv_chain[1] ;
 wire \thechain[5].chain8.inv_chain[20] ;
 wire \thechain[5].chain8.inv_chain[21] ;
 wire \thechain[5].chain8.inv_chain[22] ;
 wire \thechain[5].chain8.inv_chain[23] ;
 wire \thechain[5].chain8.inv_chain[24] ;
 wire \thechain[5].chain8.inv_chain[25] ;
 wire \thechain[5].chain8.inv_chain[26] ;
 wire \thechain[5].chain8.inv_chain[27] ;
 wire \thechain[5].chain8.inv_chain[28] ;
 wire \thechain[5].chain8.inv_chain[29] ;
 wire \thechain[5].chain8.inv_chain[2] ;
 wire \thechain[5].chain8.inv_chain[30] ;
 wire \thechain[5].chain8.inv_chain[31] ;
 wire \thechain[5].chain8.inv_chain[32] ;
 wire \thechain[5].chain8.inv_chain[33] ;
 wire \thechain[5].chain8.inv_chain[34] ;
 wire \thechain[5].chain8.inv_chain[35] ;
 wire \thechain[5].chain8.inv_chain[36] ;
 wire \thechain[5].chain8.inv_chain[37] ;
 wire \thechain[5].chain8.inv_chain[38] ;
 wire \thechain[5].chain8.inv_chain[39] ;
 wire \thechain[5].chain8.inv_chain[3] ;
 wire \thechain[5].chain8.inv_chain[40] ;
 wire \thechain[5].chain8.inv_chain[41] ;
 wire \thechain[5].chain8.inv_chain[42] ;
 wire \thechain[5].chain8.inv_chain[43] ;
 wire \thechain[5].chain8.inv_chain[44] ;
 wire \thechain[5].chain8.inv_chain[45] ;
 wire \thechain[5].chain8.inv_chain[46] ;
 wire \thechain[5].chain8.inv_chain[47] ;
 wire \thechain[5].chain8.inv_chain[48] ;
 wire \thechain[5].chain8.inv_chain[49] ;
 wire \thechain[5].chain8.inv_chain[4] ;
 wire \thechain[5].chain8.inv_chain[50] ;
 wire \thechain[5].chain8.inv_chain[51] ;
 wire \thechain[5].chain8.inv_chain[52] ;
 wire \thechain[5].chain8.inv_chain[53] ;
 wire \thechain[5].chain8.inv_chain[54] ;
 wire \thechain[5].chain8.inv_chain[55] ;
 wire \thechain[5].chain8.inv_chain[56] ;
 wire \thechain[5].chain8.inv_chain[57] ;
 wire \thechain[5].chain8.inv_chain[58] ;
 wire \thechain[5].chain8.inv_chain[59] ;
 wire \thechain[5].chain8.inv_chain[5] ;
 wire \thechain[5].chain8.inv_chain[60] ;
 wire \thechain[5].chain8.inv_chain[61] ;
 wire \thechain[5].chain8.inv_chain[62] ;
 wire \thechain[5].chain8.inv_chain[63] ;
 wire \thechain[5].chain8.inv_chain[64] ;
 wire \thechain[5].chain8.inv_chain[65] ;
 wire \thechain[5].chain8.inv_chain[66] ;
 wire \thechain[5].chain8.inv_chain[67] ;
 wire \thechain[5].chain8.inv_chain[68] ;
 wire \thechain[5].chain8.inv_chain[69] ;
 wire \thechain[5].chain8.inv_chain[6] ;
 wire \thechain[5].chain8.inv_chain[70] ;
 wire \thechain[5].chain8.inv_chain[71] ;
 wire \thechain[5].chain8.inv_chain[72] ;
 wire \thechain[5].chain8.inv_chain[73] ;
 wire \thechain[5].chain8.inv_chain[74] ;
 wire \thechain[5].chain8.inv_chain[75] ;
 wire \thechain[5].chain8.inv_chain[76] ;
 wire \thechain[5].chain8.inv_chain[77] ;
 wire \thechain[5].chain8.inv_chain[78] ;
 wire \thechain[5].chain8.inv_chain[79] ;
 wire \thechain[5].chain8.inv_chain[7] ;
 wire \thechain[5].chain8.inv_chain[80] ;
 wire \thechain[5].chain8.inv_chain[81] ;
 wire \thechain[5].chain8.inv_chain[82] ;
 wire \thechain[5].chain8.inv_chain[83] ;
 wire \thechain[5].chain8.inv_chain[84] ;
 wire \thechain[5].chain8.inv_chain[85] ;
 wire \thechain[5].chain8.inv_chain[86] ;
 wire \thechain[5].chain8.inv_chain[87] ;
 wire \thechain[5].chain8.inv_chain[88] ;
 wire \thechain[5].chain8.inv_chain[89] ;
 wire \thechain[5].chain8.inv_chain[8] ;
 wire \thechain[5].chain8.inv_chain[90] ;
 wire \thechain[5].chain8.inv_chain[91] ;
 wire \thechain[5].chain8.inv_chain[92] ;
 wire \thechain[5].chain8.inv_chain[93] ;
 wire \thechain[5].chain8.inv_chain[94] ;
 wire \thechain[5].chain8.inv_chain[95] ;
 wire \thechain[5].chain8.inv_chain[96] ;
 wire \thechain[5].chain8.inv_chain[97] ;
 wire \thechain[5].chain8.inv_chain[98] ;
 wire \thechain[5].chain8.inv_chain[99] ;
 wire \thechain[5].chain8.inv_chain[9] ;
 wire \thechain[5].chain9.dout ;
 wire \thechain[5].chain9.inv_chain[0] ;
 wire \thechain[5].chain9.inv_chain[100] ;
 wire \thechain[5].chain9.inv_chain[101] ;
 wire \thechain[5].chain9.inv_chain[102] ;
 wire \thechain[5].chain9.inv_chain[103] ;
 wire \thechain[5].chain9.inv_chain[104] ;
 wire \thechain[5].chain9.inv_chain[105] ;
 wire \thechain[5].chain9.inv_chain[106] ;
 wire \thechain[5].chain9.inv_chain[107] ;
 wire \thechain[5].chain9.inv_chain[108] ;
 wire \thechain[5].chain9.inv_chain[109] ;
 wire \thechain[5].chain9.inv_chain[10] ;
 wire \thechain[5].chain9.inv_chain[110] ;
 wire \thechain[5].chain9.inv_chain[111] ;
 wire \thechain[5].chain9.inv_chain[112] ;
 wire \thechain[5].chain9.inv_chain[113] ;
 wire \thechain[5].chain9.inv_chain[114] ;
 wire \thechain[5].chain9.inv_chain[115] ;
 wire \thechain[5].chain9.inv_chain[116] ;
 wire \thechain[5].chain9.inv_chain[117] ;
 wire \thechain[5].chain9.inv_chain[118] ;
 wire \thechain[5].chain9.inv_chain[119] ;
 wire \thechain[5].chain9.inv_chain[11] ;
 wire \thechain[5].chain9.inv_chain[120] ;
 wire \thechain[5].chain9.inv_chain[121] ;
 wire \thechain[5].chain9.inv_chain[122] ;
 wire \thechain[5].chain9.inv_chain[123] ;
 wire \thechain[5].chain9.inv_chain[124] ;
 wire \thechain[5].chain9.inv_chain[125] ;
 wire \thechain[5].chain9.inv_chain[126] ;
 wire \thechain[5].chain9.inv_chain[127] ;
 wire \thechain[5].chain9.inv_chain[128] ;
 wire \thechain[5].chain9.inv_chain[129] ;
 wire \thechain[5].chain9.inv_chain[12] ;
 wire \thechain[5].chain9.inv_chain[130] ;
 wire \thechain[5].chain9.inv_chain[131] ;
 wire \thechain[5].chain9.inv_chain[132] ;
 wire \thechain[5].chain9.inv_chain[133] ;
 wire \thechain[5].chain9.inv_chain[134] ;
 wire \thechain[5].chain9.inv_chain[135] ;
 wire \thechain[5].chain9.inv_chain[136] ;
 wire \thechain[5].chain9.inv_chain[137] ;
 wire \thechain[5].chain9.inv_chain[138] ;
 wire \thechain[5].chain9.inv_chain[139] ;
 wire \thechain[5].chain9.inv_chain[13] ;
 wire \thechain[5].chain9.inv_chain[140] ;
 wire \thechain[5].chain9.inv_chain[141] ;
 wire \thechain[5].chain9.inv_chain[142] ;
 wire \thechain[5].chain9.inv_chain[143] ;
 wire \thechain[5].chain9.inv_chain[144] ;
 wire \thechain[5].chain9.inv_chain[145] ;
 wire \thechain[5].chain9.inv_chain[146] ;
 wire \thechain[5].chain9.inv_chain[147] ;
 wire \thechain[5].chain9.inv_chain[148] ;
 wire \thechain[5].chain9.inv_chain[149] ;
 wire \thechain[5].chain9.inv_chain[14] ;
 wire \thechain[5].chain9.inv_chain[150] ;
 wire \thechain[5].chain9.inv_chain[151] ;
 wire \thechain[5].chain9.inv_chain[152] ;
 wire \thechain[5].chain9.inv_chain[153] ;
 wire \thechain[5].chain9.inv_chain[154] ;
 wire \thechain[5].chain9.inv_chain[155] ;
 wire \thechain[5].chain9.inv_chain[156] ;
 wire \thechain[5].chain9.inv_chain[157] ;
 wire \thechain[5].chain9.inv_chain[158] ;
 wire \thechain[5].chain9.inv_chain[159] ;
 wire \thechain[5].chain9.inv_chain[15] ;
 wire \thechain[5].chain9.inv_chain[160] ;
 wire \thechain[5].chain9.inv_chain[161] ;
 wire \thechain[5].chain9.inv_chain[162] ;
 wire \thechain[5].chain9.inv_chain[163] ;
 wire \thechain[5].chain9.inv_chain[164] ;
 wire \thechain[5].chain9.inv_chain[165] ;
 wire \thechain[5].chain9.inv_chain[166] ;
 wire \thechain[5].chain9.inv_chain[167] ;
 wire \thechain[5].chain9.inv_chain[168] ;
 wire \thechain[5].chain9.inv_chain[169] ;
 wire \thechain[5].chain9.inv_chain[16] ;
 wire \thechain[5].chain9.inv_chain[170] ;
 wire \thechain[5].chain9.inv_chain[171] ;
 wire \thechain[5].chain9.inv_chain[172] ;
 wire \thechain[5].chain9.inv_chain[173] ;
 wire \thechain[5].chain9.inv_chain[174] ;
 wire \thechain[5].chain9.inv_chain[175] ;
 wire \thechain[5].chain9.inv_chain[176] ;
 wire \thechain[5].chain9.inv_chain[177] ;
 wire \thechain[5].chain9.inv_chain[178] ;
 wire \thechain[5].chain9.inv_chain[179] ;
 wire \thechain[5].chain9.inv_chain[17] ;
 wire \thechain[5].chain9.inv_chain[180] ;
 wire \thechain[5].chain9.inv_chain[181] ;
 wire \thechain[5].chain9.inv_chain[182] ;
 wire \thechain[5].chain9.inv_chain[183] ;
 wire \thechain[5].chain9.inv_chain[184] ;
 wire \thechain[5].chain9.inv_chain[185] ;
 wire \thechain[5].chain9.inv_chain[186] ;
 wire \thechain[5].chain9.inv_chain[187] ;
 wire \thechain[5].chain9.inv_chain[188] ;
 wire \thechain[5].chain9.inv_chain[189] ;
 wire \thechain[5].chain9.inv_chain[18] ;
 wire \thechain[5].chain9.inv_chain[190] ;
 wire \thechain[5].chain9.inv_chain[191] ;
 wire \thechain[5].chain9.inv_chain[192] ;
 wire \thechain[5].chain9.inv_chain[193] ;
 wire \thechain[5].chain9.inv_chain[194] ;
 wire \thechain[5].chain9.inv_chain[195] ;
 wire \thechain[5].chain9.inv_chain[196] ;
 wire \thechain[5].chain9.inv_chain[197] ;
 wire \thechain[5].chain9.inv_chain[198] ;
 wire \thechain[5].chain9.inv_chain[199] ;
 wire \thechain[5].chain9.inv_chain[19] ;
 wire \thechain[5].chain9.inv_chain[1] ;
 wire \thechain[5].chain9.inv_chain[200] ;
 wire \thechain[5].chain9.inv_chain[201] ;
 wire \thechain[5].chain9.inv_chain[202] ;
 wire \thechain[5].chain9.inv_chain[203] ;
 wire \thechain[5].chain9.inv_chain[204] ;
 wire \thechain[5].chain9.inv_chain[205] ;
 wire \thechain[5].chain9.inv_chain[206] ;
 wire \thechain[5].chain9.inv_chain[207] ;
 wire \thechain[5].chain9.inv_chain[208] ;
 wire \thechain[5].chain9.inv_chain[209] ;
 wire \thechain[5].chain9.inv_chain[20] ;
 wire \thechain[5].chain9.inv_chain[210] ;
 wire \thechain[5].chain9.inv_chain[211] ;
 wire \thechain[5].chain9.inv_chain[212] ;
 wire \thechain[5].chain9.inv_chain[213] ;
 wire \thechain[5].chain9.inv_chain[214] ;
 wire \thechain[5].chain9.inv_chain[215] ;
 wire \thechain[5].chain9.inv_chain[216] ;
 wire \thechain[5].chain9.inv_chain[217] ;
 wire \thechain[5].chain9.inv_chain[218] ;
 wire \thechain[5].chain9.inv_chain[219] ;
 wire \thechain[5].chain9.inv_chain[21] ;
 wire \thechain[5].chain9.inv_chain[220] ;
 wire \thechain[5].chain9.inv_chain[221] ;
 wire \thechain[5].chain9.inv_chain[222] ;
 wire \thechain[5].chain9.inv_chain[223] ;
 wire \thechain[5].chain9.inv_chain[224] ;
 wire \thechain[5].chain9.inv_chain[225] ;
 wire \thechain[5].chain9.inv_chain[226] ;
 wire \thechain[5].chain9.inv_chain[227] ;
 wire \thechain[5].chain9.inv_chain[228] ;
 wire \thechain[5].chain9.inv_chain[229] ;
 wire \thechain[5].chain9.inv_chain[22] ;
 wire \thechain[5].chain9.inv_chain[230] ;
 wire \thechain[5].chain9.inv_chain[231] ;
 wire \thechain[5].chain9.inv_chain[232] ;
 wire \thechain[5].chain9.inv_chain[233] ;
 wire \thechain[5].chain9.inv_chain[234] ;
 wire \thechain[5].chain9.inv_chain[235] ;
 wire \thechain[5].chain9.inv_chain[236] ;
 wire \thechain[5].chain9.inv_chain[237] ;
 wire \thechain[5].chain9.inv_chain[238] ;
 wire \thechain[5].chain9.inv_chain[239] ;
 wire \thechain[5].chain9.inv_chain[23] ;
 wire \thechain[5].chain9.inv_chain[240] ;
 wire \thechain[5].chain9.inv_chain[241] ;
 wire \thechain[5].chain9.inv_chain[242] ;
 wire \thechain[5].chain9.inv_chain[243] ;
 wire \thechain[5].chain9.inv_chain[244] ;
 wire \thechain[5].chain9.inv_chain[245] ;
 wire \thechain[5].chain9.inv_chain[246] ;
 wire \thechain[5].chain9.inv_chain[247] ;
 wire \thechain[5].chain9.inv_chain[248] ;
 wire \thechain[5].chain9.inv_chain[249] ;
 wire \thechain[5].chain9.inv_chain[24] ;
 wire \thechain[5].chain9.inv_chain[250] ;
 wire \thechain[5].chain9.inv_chain[251] ;
 wire \thechain[5].chain9.inv_chain[252] ;
 wire \thechain[5].chain9.inv_chain[253] ;
 wire \thechain[5].chain9.inv_chain[254] ;
 wire \thechain[5].chain9.inv_chain[255] ;
 wire \thechain[5].chain9.inv_chain[256] ;
 wire \thechain[5].chain9.inv_chain[25] ;
 wire \thechain[5].chain9.inv_chain[26] ;
 wire \thechain[5].chain9.inv_chain[27] ;
 wire \thechain[5].chain9.inv_chain[28] ;
 wire \thechain[5].chain9.inv_chain[29] ;
 wire \thechain[5].chain9.inv_chain[2] ;
 wire \thechain[5].chain9.inv_chain[30] ;
 wire \thechain[5].chain9.inv_chain[31] ;
 wire \thechain[5].chain9.inv_chain[32] ;
 wire \thechain[5].chain9.inv_chain[33] ;
 wire \thechain[5].chain9.inv_chain[34] ;
 wire \thechain[5].chain9.inv_chain[35] ;
 wire \thechain[5].chain9.inv_chain[36] ;
 wire \thechain[5].chain9.inv_chain[37] ;
 wire \thechain[5].chain9.inv_chain[38] ;
 wire \thechain[5].chain9.inv_chain[39] ;
 wire \thechain[5].chain9.inv_chain[3] ;
 wire \thechain[5].chain9.inv_chain[40] ;
 wire \thechain[5].chain9.inv_chain[41] ;
 wire \thechain[5].chain9.inv_chain[42] ;
 wire \thechain[5].chain9.inv_chain[43] ;
 wire \thechain[5].chain9.inv_chain[44] ;
 wire \thechain[5].chain9.inv_chain[45] ;
 wire \thechain[5].chain9.inv_chain[46] ;
 wire \thechain[5].chain9.inv_chain[47] ;
 wire \thechain[5].chain9.inv_chain[48] ;
 wire \thechain[5].chain9.inv_chain[49] ;
 wire \thechain[5].chain9.inv_chain[4] ;
 wire \thechain[5].chain9.inv_chain[50] ;
 wire \thechain[5].chain9.inv_chain[51] ;
 wire \thechain[5].chain9.inv_chain[52] ;
 wire \thechain[5].chain9.inv_chain[53] ;
 wire \thechain[5].chain9.inv_chain[54] ;
 wire \thechain[5].chain9.inv_chain[55] ;
 wire \thechain[5].chain9.inv_chain[56] ;
 wire \thechain[5].chain9.inv_chain[57] ;
 wire \thechain[5].chain9.inv_chain[58] ;
 wire \thechain[5].chain9.inv_chain[59] ;
 wire \thechain[5].chain9.inv_chain[5] ;
 wire \thechain[5].chain9.inv_chain[60] ;
 wire \thechain[5].chain9.inv_chain[61] ;
 wire \thechain[5].chain9.inv_chain[62] ;
 wire \thechain[5].chain9.inv_chain[63] ;
 wire \thechain[5].chain9.inv_chain[64] ;
 wire \thechain[5].chain9.inv_chain[65] ;
 wire \thechain[5].chain9.inv_chain[66] ;
 wire \thechain[5].chain9.inv_chain[67] ;
 wire \thechain[5].chain9.inv_chain[68] ;
 wire \thechain[5].chain9.inv_chain[69] ;
 wire \thechain[5].chain9.inv_chain[6] ;
 wire \thechain[5].chain9.inv_chain[70] ;
 wire \thechain[5].chain9.inv_chain[71] ;
 wire \thechain[5].chain9.inv_chain[72] ;
 wire \thechain[5].chain9.inv_chain[73] ;
 wire \thechain[5].chain9.inv_chain[74] ;
 wire \thechain[5].chain9.inv_chain[75] ;
 wire \thechain[5].chain9.inv_chain[76] ;
 wire \thechain[5].chain9.inv_chain[77] ;
 wire \thechain[5].chain9.inv_chain[78] ;
 wire \thechain[5].chain9.inv_chain[79] ;
 wire \thechain[5].chain9.inv_chain[7] ;
 wire \thechain[5].chain9.inv_chain[80] ;
 wire \thechain[5].chain9.inv_chain[81] ;
 wire \thechain[5].chain9.inv_chain[82] ;
 wire \thechain[5].chain9.inv_chain[83] ;
 wire \thechain[5].chain9.inv_chain[84] ;
 wire \thechain[5].chain9.inv_chain[85] ;
 wire \thechain[5].chain9.inv_chain[86] ;
 wire \thechain[5].chain9.inv_chain[87] ;
 wire \thechain[5].chain9.inv_chain[88] ;
 wire \thechain[5].chain9.inv_chain[89] ;
 wire \thechain[5].chain9.inv_chain[8] ;
 wire \thechain[5].chain9.inv_chain[90] ;
 wire \thechain[5].chain9.inv_chain[91] ;
 wire \thechain[5].chain9.inv_chain[92] ;
 wire \thechain[5].chain9.inv_chain[93] ;
 wire \thechain[5].chain9.inv_chain[94] ;
 wire \thechain[5].chain9.inv_chain[95] ;
 wire \thechain[5].chain9.inv_chain[96] ;
 wire \thechain[5].chain9.inv_chain[97] ;
 wire \thechain[5].chain9.inv_chain[98] ;
 wire \thechain[5].chain9.inv_chain[99] ;
 wire \thechain[5].chain9.inv_chain[9] ;
 wire \thechain[6].chain1.dout ;
 wire \thechain[6].chain1.inv_chain[0] ;
 wire \thechain[6].chain1.inv_chain[1] ;
 wire \thechain[6].chain1.inv_chain[2] ;
 wire \thechain[6].chain2.dout ;
 wire \thechain[6].chain2.inv_chain[0] ;
 wire \thechain[6].chain2.inv_chain[1] ;
 wire \thechain[6].chain2.inv_chain[2] ;
 wire \thechain[6].chain2.inv_chain[3] ;
 wire \thechain[6].chain2.inv_chain[4] ;
 wire \thechain[6].chain3.dout ;
 wire \thechain[6].chain3.inv_chain[0] ;
 wire \thechain[6].chain3.inv_chain[1] ;
 wire \thechain[6].chain3.inv_chain[2] ;
 wire \thechain[6].chain3.inv_chain[3] ;
 wire \thechain[6].chain3.inv_chain[4] ;
 wire \thechain[6].chain3.inv_chain[5] ;
 wire \thechain[6].chain3.inv_chain[6] ;
 wire \thechain[6].chain3.inv_chain[7] ;
 wire \thechain[6].chain3.inv_chain[8] ;
 wire \thechain[6].chain4.dout ;
 wire \thechain[6].chain4.inv_chain[0] ;
 wire \thechain[6].chain4.inv_chain[10] ;
 wire \thechain[6].chain4.inv_chain[11] ;
 wire \thechain[6].chain4.inv_chain[12] ;
 wire \thechain[6].chain4.inv_chain[13] ;
 wire \thechain[6].chain4.inv_chain[14] ;
 wire \thechain[6].chain4.inv_chain[15] ;
 wire \thechain[6].chain4.inv_chain[16] ;
 wire \thechain[6].chain4.inv_chain[1] ;
 wire \thechain[6].chain4.inv_chain[2] ;
 wire \thechain[6].chain4.inv_chain[3] ;
 wire \thechain[6].chain4.inv_chain[4] ;
 wire \thechain[6].chain4.inv_chain[5] ;
 wire \thechain[6].chain4.inv_chain[6] ;
 wire \thechain[6].chain4.inv_chain[7] ;
 wire \thechain[6].chain4.inv_chain[8] ;
 wire \thechain[6].chain4.inv_chain[9] ;
 wire \thechain[6].chain5.dout ;
 wire \thechain[6].chain5.inv_chain[0] ;
 wire \thechain[6].chain5.inv_chain[10] ;
 wire \thechain[6].chain5.inv_chain[11] ;
 wire \thechain[6].chain5.inv_chain[12] ;
 wire \thechain[6].chain5.inv_chain[13] ;
 wire \thechain[6].chain5.inv_chain[14] ;
 wire \thechain[6].chain5.inv_chain[15] ;
 wire \thechain[6].chain5.inv_chain[16] ;
 wire \thechain[6].chain5.inv_chain[17] ;
 wire \thechain[6].chain5.inv_chain[18] ;
 wire \thechain[6].chain5.inv_chain[19] ;
 wire \thechain[6].chain5.inv_chain[1] ;
 wire \thechain[6].chain5.inv_chain[20] ;
 wire \thechain[6].chain5.inv_chain[21] ;
 wire \thechain[6].chain5.inv_chain[22] ;
 wire \thechain[6].chain5.inv_chain[23] ;
 wire \thechain[6].chain5.inv_chain[24] ;
 wire \thechain[6].chain5.inv_chain[25] ;
 wire \thechain[6].chain5.inv_chain[26] ;
 wire \thechain[6].chain5.inv_chain[27] ;
 wire \thechain[6].chain5.inv_chain[28] ;
 wire \thechain[6].chain5.inv_chain[29] ;
 wire \thechain[6].chain5.inv_chain[2] ;
 wire \thechain[6].chain5.inv_chain[30] ;
 wire \thechain[6].chain5.inv_chain[31] ;
 wire \thechain[6].chain5.inv_chain[32] ;
 wire \thechain[6].chain5.inv_chain[3] ;
 wire \thechain[6].chain5.inv_chain[4] ;
 wire \thechain[6].chain5.inv_chain[5] ;
 wire \thechain[6].chain5.inv_chain[6] ;
 wire \thechain[6].chain5.inv_chain[7] ;
 wire \thechain[6].chain5.inv_chain[8] ;
 wire \thechain[6].chain5.inv_chain[9] ;
 wire \thechain[6].chain6.dout ;
 wire \thechain[6].chain6.inv_chain[0] ;
 wire \thechain[6].chain6.inv_chain[10] ;
 wire \thechain[6].chain6.inv_chain[11] ;
 wire \thechain[6].chain6.inv_chain[12] ;
 wire \thechain[6].chain6.inv_chain[13] ;
 wire \thechain[6].chain6.inv_chain[14] ;
 wire \thechain[6].chain6.inv_chain[15] ;
 wire \thechain[6].chain6.inv_chain[16] ;
 wire \thechain[6].chain6.inv_chain[17] ;
 wire \thechain[6].chain6.inv_chain[18] ;
 wire \thechain[6].chain6.inv_chain[19] ;
 wire \thechain[6].chain6.inv_chain[1] ;
 wire \thechain[6].chain6.inv_chain[20] ;
 wire \thechain[6].chain6.inv_chain[21] ;
 wire \thechain[6].chain6.inv_chain[22] ;
 wire \thechain[6].chain6.inv_chain[23] ;
 wire \thechain[6].chain6.inv_chain[24] ;
 wire \thechain[6].chain6.inv_chain[25] ;
 wire \thechain[6].chain6.inv_chain[26] ;
 wire \thechain[6].chain6.inv_chain[27] ;
 wire \thechain[6].chain6.inv_chain[28] ;
 wire \thechain[6].chain6.inv_chain[29] ;
 wire \thechain[6].chain6.inv_chain[2] ;
 wire \thechain[6].chain6.inv_chain[30] ;
 wire \thechain[6].chain6.inv_chain[31] ;
 wire \thechain[6].chain6.inv_chain[32] ;
 wire \thechain[6].chain6.inv_chain[33] ;
 wire \thechain[6].chain6.inv_chain[34] ;
 wire \thechain[6].chain6.inv_chain[35] ;
 wire \thechain[6].chain6.inv_chain[36] ;
 wire \thechain[6].chain6.inv_chain[37] ;
 wire \thechain[6].chain6.inv_chain[38] ;
 wire \thechain[6].chain6.inv_chain[39] ;
 wire \thechain[6].chain6.inv_chain[3] ;
 wire \thechain[6].chain6.inv_chain[40] ;
 wire \thechain[6].chain6.inv_chain[41] ;
 wire \thechain[6].chain6.inv_chain[42] ;
 wire \thechain[6].chain6.inv_chain[43] ;
 wire \thechain[6].chain6.inv_chain[44] ;
 wire \thechain[6].chain6.inv_chain[45] ;
 wire \thechain[6].chain6.inv_chain[46] ;
 wire \thechain[6].chain6.inv_chain[47] ;
 wire \thechain[6].chain6.inv_chain[48] ;
 wire \thechain[6].chain6.inv_chain[49] ;
 wire \thechain[6].chain6.inv_chain[4] ;
 wire \thechain[6].chain6.inv_chain[50] ;
 wire \thechain[6].chain6.inv_chain[51] ;
 wire \thechain[6].chain6.inv_chain[52] ;
 wire \thechain[6].chain6.inv_chain[53] ;
 wire \thechain[6].chain6.inv_chain[54] ;
 wire \thechain[6].chain6.inv_chain[55] ;
 wire \thechain[6].chain6.inv_chain[56] ;
 wire \thechain[6].chain6.inv_chain[57] ;
 wire \thechain[6].chain6.inv_chain[58] ;
 wire \thechain[6].chain6.inv_chain[59] ;
 wire \thechain[6].chain6.inv_chain[5] ;
 wire \thechain[6].chain6.inv_chain[60] ;
 wire \thechain[6].chain6.inv_chain[61] ;
 wire \thechain[6].chain6.inv_chain[62] ;
 wire \thechain[6].chain6.inv_chain[63] ;
 wire \thechain[6].chain6.inv_chain[64] ;
 wire \thechain[6].chain6.inv_chain[6] ;
 wire \thechain[6].chain6.inv_chain[7] ;
 wire \thechain[6].chain6.inv_chain[8] ;
 wire \thechain[6].chain6.inv_chain[9] ;
 wire \thechain[6].chain7.dout ;
 wire \thechain[6].chain7.inv_chain[0] ;
 wire \thechain[6].chain7.inv_chain[100] ;
 wire \thechain[6].chain7.inv_chain[101] ;
 wire \thechain[6].chain7.inv_chain[102] ;
 wire \thechain[6].chain7.inv_chain[103] ;
 wire \thechain[6].chain7.inv_chain[104] ;
 wire \thechain[6].chain7.inv_chain[105] ;
 wire \thechain[6].chain7.inv_chain[106] ;
 wire \thechain[6].chain7.inv_chain[107] ;
 wire \thechain[6].chain7.inv_chain[108] ;
 wire \thechain[6].chain7.inv_chain[109] ;
 wire \thechain[6].chain7.inv_chain[10] ;
 wire \thechain[6].chain7.inv_chain[110] ;
 wire \thechain[6].chain7.inv_chain[111] ;
 wire \thechain[6].chain7.inv_chain[112] ;
 wire \thechain[6].chain7.inv_chain[113] ;
 wire \thechain[6].chain7.inv_chain[114] ;
 wire \thechain[6].chain7.inv_chain[115] ;
 wire \thechain[6].chain7.inv_chain[116] ;
 wire \thechain[6].chain7.inv_chain[117] ;
 wire \thechain[6].chain7.inv_chain[118] ;
 wire \thechain[6].chain7.inv_chain[119] ;
 wire \thechain[6].chain7.inv_chain[11] ;
 wire \thechain[6].chain7.inv_chain[120] ;
 wire \thechain[6].chain7.inv_chain[121] ;
 wire \thechain[6].chain7.inv_chain[122] ;
 wire \thechain[6].chain7.inv_chain[123] ;
 wire \thechain[6].chain7.inv_chain[124] ;
 wire \thechain[6].chain7.inv_chain[125] ;
 wire \thechain[6].chain7.inv_chain[126] ;
 wire \thechain[6].chain7.inv_chain[127] ;
 wire \thechain[6].chain7.inv_chain[128] ;
 wire \thechain[6].chain7.inv_chain[12] ;
 wire \thechain[6].chain7.inv_chain[13] ;
 wire \thechain[6].chain7.inv_chain[14] ;
 wire \thechain[6].chain7.inv_chain[15] ;
 wire \thechain[6].chain7.inv_chain[16] ;
 wire \thechain[6].chain7.inv_chain[17] ;
 wire \thechain[6].chain7.inv_chain[18] ;
 wire \thechain[6].chain7.inv_chain[19] ;
 wire \thechain[6].chain7.inv_chain[1] ;
 wire \thechain[6].chain7.inv_chain[20] ;
 wire \thechain[6].chain7.inv_chain[21] ;
 wire \thechain[6].chain7.inv_chain[22] ;
 wire \thechain[6].chain7.inv_chain[23] ;
 wire \thechain[6].chain7.inv_chain[24] ;
 wire \thechain[6].chain7.inv_chain[25] ;
 wire \thechain[6].chain7.inv_chain[26] ;
 wire \thechain[6].chain7.inv_chain[27] ;
 wire \thechain[6].chain7.inv_chain[28] ;
 wire \thechain[6].chain7.inv_chain[29] ;
 wire \thechain[6].chain7.inv_chain[2] ;
 wire \thechain[6].chain7.inv_chain[30] ;
 wire \thechain[6].chain7.inv_chain[31] ;
 wire \thechain[6].chain7.inv_chain[32] ;
 wire \thechain[6].chain7.inv_chain[33] ;
 wire \thechain[6].chain7.inv_chain[34] ;
 wire \thechain[6].chain7.inv_chain[35] ;
 wire \thechain[6].chain7.inv_chain[36] ;
 wire \thechain[6].chain7.inv_chain[37] ;
 wire \thechain[6].chain7.inv_chain[38] ;
 wire \thechain[6].chain7.inv_chain[39] ;
 wire \thechain[6].chain7.inv_chain[3] ;
 wire \thechain[6].chain7.inv_chain[40] ;
 wire \thechain[6].chain7.inv_chain[41] ;
 wire \thechain[6].chain7.inv_chain[42] ;
 wire \thechain[6].chain7.inv_chain[43] ;
 wire \thechain[6].chain7.inv_chain[44] ;
 wire \thechain[6].chain7.inv_chain[45] ;
 wire \thechain[6].chain7.inv_chain[46] ;
 wire \thechain[6].chain7.inv_chain[47] ;
 wire \thechain[6].chain7.inv_chain[48] ;
 wire \thechain[6].chain7.inv_chain[49] ;
 wire \thechain[6].chain7.inv_chain[4] ;
 wire \thechain[6].chain7.inv_chain[50] ;
 wire \thechain[6].chain7.inv_chain[51] ;
 wire \thechain[6].chain7.inv_chain[52] ;
 wire \thechain[6].chain7.inv_chain[53] ;
 wire \thechain[6].chain7.inv_chain[54] ;
 wire \thechain[6].chain7.inv_chain[55] ;
 wire \thechain[6].chain7.inv_chain[56] ;
 wire \thechain[6].chain7.inv_chain[57] ;
 wire \thechain[6].chain7.inv_chain[58] ;
 wire \thechain[6].chain7.inv_chain[59] ;
 wire \thechain[6].chain7.inv_chain[5] ;
 wire \thechain[6].chain7.inv_chain[60] ;
 wire \thechain[6].chain7.inv_chain[61] ;
 wire \thechain[6].chain7.inv_chain[62] ;
 wire \thechain[6].chain7.inv_chain[63] ;
 wire \thechain[6].chain7.inv_chain[64] ;
 wire \thechain[6].chain7.inv_chain[65] ;
 wire \thechain[6].chain7.inv_chain[66] ;
 wire \thechain[6].chain7.inv_chain[67] ;
 wire \thechain[6].chain7.inv_chain[68] ;
 wire \thechain[6].chain7.inv_chain[69] ;
 wire \thechain[6].chain7.inv_chain[6] ;
 wire \thechain[6].chain7.inv_chain[70] ;
 wire \thechain[6].chain7.inv_chain[71] ;
 wire \thechain[6].chain7.inv_chain[72] ;
 wire \thechain[6].chain7.inv_chain[73] ;
 wire \thechain[6].chain7.inv_chain[74] ;
 wire \thechain[6].chain7.inv_chain[75] ;
 wire \thechain[6].chain7.inv_chain[76] ;
 wire \thechain[6].chain7.inv_chain[77] ;
 wire \thechain[6].chain7.inv_chain[78] ;
 wire \thechain[6].chain7.inv_chain[79] ;
 wire \thechain[6].chain7.inv_chain[7] ;
 wire \thechain[6].chain7.inv_chain[80] ;
 wire \thechain[6].chain7.inv_chain[81] ;
 wire \thechain[6].chain7.inv_chain[82] ;
 wire \thechain[6].chain7.inv_chain[83] ;
 wire \thechain[6].chain7.inv_chain[84] ;
 wire \thechain[6].chain7.inv_chain[85] ;
 wire \thechain[6].chain7.inv_chain[86] ;
 wire \thechain[6].chain7.inv_chain[87] ;
 wire \thechain[6].chain7.inv_chain[88] ;
 wire \thechain[6].chain7.inv_chain[89] ;
 wire \thechain[6].chain7.inv_chain[8] ;
 wire \thechain[6].chain7.inv_chain[90] ;
 wire \thechain[6].chain7.inv_chain[91] ;
 wire \thechain[6].chain7.inv_chain[92] ;
 wire \thechain[6].chain7.inv_chain[93] ;
 wire \thechain[6].chain7.inv_chain[94] ;
 wire \thechain[6].chain7.inv_chain[95] ;
 wire \thechain[6].chain7.inv_chain[96] ;
 wire \thechain[6].chain7.inv_chain[97] ;
 wire \thechain[6].chain7.inv_chain[98] ;
 wire \thechain[6].chain7.inv_chain[99] ;
 wire \thechain[6].chain7.inv_chain[9] ;
 wire \thechain[6].chain8.dout ;
 wire \thechain[6].chain8.inv_chain[0] ;
 wire \thechain[6].chain8.inv_chain[100] ;
 wire \thechain[6].chain8.inv_chain[101] ;
 wire \thechain[6].chain8.inv_chain[102] ;
 wire \thechain[6].chain8.inv_chain[103] ;
 wire \thechain[6].chain8.inv_chain[104] ;
 wire \thechain[6].chain8.inv_chain[105] ;
 wire \thechain[6].chain8.inv_chain[106] ;
 wire \thechain[6].chain8.inv_chain[107] ;
 wire \thechain[6].chain8.inv_chain[108] ;
 wire \thechain[6].chain8.inv_chain[109] ;
 wire \thechain[6].chain8.inv_chain[10] ;
 wire \thechain[6].chain8.inv_chain[110] ;
 wire \thechain[6].chain8.inv_chain[111] ;
 wire \thechain[6].chain8.inv_chain[112] ;
 wire \thechain[6].chain8.inv_chain[113] ;
 wire \thechain[6].chain8.inv_chain[114] ;
 wire \thechain[6].chain8.inv_chain[115] ;
 wire \thechain[6].chain8.inv_chain[116] ;
 wire \thechain[6].chain8.inv_chain[117] ;
 wire \thechain[6].chain8.inv_chain[118] ;
 wire \thechain[6].chain8.inv_chain[119] ;
 wire \thechain[6].chain8.inv_chain[11] ;
 wire \thechain[6].chain8.inv_chain[120] ;
 wire \thechain[6].chain8.inv_chain[121] ;
 wire \thechain[6].chain8.inv_chain[122] ;
 wire \thechain[6].chain8.inv_chain[123] ;
 wire \thechain[6].chain8.inv_chain[124] ;
 wire \thechain[6].chain8.inv_chain[125] ;
 wire \thechain[6].chain8.inv_chain[126] ;
 wire \thechain[6].chain8.inv_chain[127] ;
 wire \thechain[6].chain8.inv_chain[128] ;
 wire \thechain[6].chain8.inv_chain[129] ;
 wire \thechain[6].chain8.inv_chain[12] ;
 wire \thechain[6].chain8.inv_chain[130] ;
 wire \thechain[6].chain8.inv_chain[131] ;
 wire \thechain[6].chain8.inv_chain[132] ;
 wire \thechain[6].chain8.inv_chain[133] ;
 wire \thechain[6].chain8.inv_chain[134] ;
 wire \thechain[6].chain8.inv_chain[135] ;
 wire \thechain[6].chain8.inv_chain[136] ;
 wire \thechain[6].chain8.inv_chain[137] ;
 wire \thechain[6].chain8.inv_chain[138] ;
 wire \thechain[6].chain8.inv_chain[139] ;
 wire \thechain[6].chain8.inv_chain[13] ;
 wire \thechain[6].chain8.inv_chain[140] ;
 wire \thechain[6].chain8.inv_chain[141] ;
 wire \thechain[6].chain8.inv_chain[142] ;
 wire \thechain[6].chain8.inv_chain[143] ;
 wire \thechain[6].chain8.inv_chain[144] ;
 wire \thechain[6].chain8.inv_chain[145] ;
 wire \thechain[6].chain8.inv_chain[146] ;
 wire \thechain[6].chain8.inv_chain[147] ;
 wire \thechain[6].chain8.inv_chain[148] ;
 wire \thechain[6].chain8.inv_chain[149] ;
 wire \thechain[6].chain8.inv_chain[14] ;
 wire \thechain[6].chain8.inv_chain[150] ;
 wire \thechain[6].chain8.inv_chain[151] ;
 wire \thechain[6].chain8.inv_chain[152] ;
 wire \thechain[6].chain8.inv_chain[153] ;
 wire \thechain[6].chain8.inv_chain[154] ;
 wire \thechain[6].chain8.inv_chain[155] ;
 wire \thechain[6].chain8.inv_chain[156] ;
 wire \thechain[6].chain8.inv_chain[157] ;
 wire \thechain[6].chain8.inv_chain[158] ;
 wire \thechain[6].chain8.inv_chain[159] ;
 wire \thechain[6].chain8.inv_chain[15] ;
 wire \thechain[6].chain8.inv_chain[160] ;
 wire \thechain[6].chain8.inv_chain[161] ;
 wire \thechain[6].chain8.inv_chain[162] ;
 wire \thechain[6].chain8.inv_chain[163] ;
 wire \thechain[6].chain8.inv_chain[164] ;
 wire \thechain[6].chain8.inv_chain[165] ;
 wire \thechain[6].chain8.inv_chain[166] ;
 wire \thechain[6].chain8.inv_chain[167] ;
 wire \thechain[6].chain8.inv_chain[168] ;
 wire \thechain[6].chain8.inv_chain[169] ;
 wire \thechain[6].chain8.inv_chain[16] ;
 wire \thechain[6].chain8.inv_chain[170] ;
 wire \thechain[6].chain8.inv_chain[171] ;
 wire \thechain[6].chain8.inv_chain[172] ;
 wire \thechain[6].chain8.inv_chain[173] ;
 wire \thechain[6].chain8.inv_chain[174] ;
 wire \thechain[6].chain8.inv_chain[175] ;
 wire \thechain[6].chain8.inv_chain[176] ;
 wire \thechain[6].chain8.inv_chain[177] ;
 wire \thechain[6].chain8.inv_chain[178] ;
 wire \thechain[6].chain8.inv_chain[179] ;
 wire \thechain[6].chain8.inv_chain[17] ;
 wire \thechain[6].chain8.inv_chain[180] ;
 wire \thechain[6].chain8.inv_chain[181] ;
 wire \thechain[6].chain8.inv_chain[182] ;
 wire \thechain[6].chain8.inv_chain[183] ;
 wire \thechain[6].chain8.inv_chain[184] ;
 wire \thechain[6].chain8.inv_chain[185] ;
 wire \thechain[6].chain8.inv_chain[186] ;
 wire \thechain[6].chain8.inv_chain[187] ;
 wire \thechain[6].chain8.inv_chain[188] ;
 wire \thechain[6].chain8.inv_chain[189] ;
 wire \thechain[6].chain8.inv_chain[18] ;
 wire \thechain[6].chain8.inv_chain[190] ;
 wire \thechain[6].chain8.inv_chain[191] ;
 wire \thechain[6].chain8.inv_chain[192] ;
 wire \thechain[6].chain8.inv_chain[19] ;
 wire \thechain[6].chain8.inv_chain[1] ;
 wire \thechain[6].chain8.inv_chain[20] ;
 wire \thechain[6].chain8.inv_chain[21] ;
 wire \thechain[6].chain8.inv_chain[22] ;
 wire \thechain[6].chain8.inv_chain[23] ;
 wire \thechain[6].chain8.inv_chain[24] ;
 wire \thechain[6].chain8.inv_chain[25] ;
 wire \thechain[6].chain8.inv_chain[26] ;
 wire \thechain[6].chain8.inv_chain[27] ;
 wire \thechain[6].chain8.inv_chain[28] ;
 wire \thechain[6].chain8.inv_chain[29] ;
 wire \thechain[6].chain8.inv_chain[2] ;
 wire \thechain[6].chain8.inv_chain[30] ;
 wire \thechain[6].chain8.inv_chain[31] ;
 wire \thechain[6].chain8.inv_chain[32] ;
 wire \thechain[6].chain8.inv_chain[33] ;
 wire \thechain[6].chain8.inv_chain[34] ;
 wire \thechain[6].chain8.inv_chain[35] ;
 wire \thechain[6].chain8.inv_chain[36] ;
 wire \thechain[6].chain8.inv_chain[37] ;
 wire \thechain[6].chain8.inv_chain[38] ;
 wire \thechain[6].chain8.inv_chain[39] ;
 wire \thechain[6].chain8.inv_chain[3] ;
 wire \thechain[6].chain8.inv_chain[40] ;
 wire \thechain[6].chain8.inv_chain[41] ;
 wire \thechain[6].chain8.inv_chain[42] ;
 wire \thechain[6].chain8.inv_chain[43] ;
 wire \thechain[6].chain8.inv_chain[44] ;
 wire \thechain[6].chain8.inv_chain[45] ;
 wire \thechain[6].chain8.inv_chain[46] ;
 wire \thechain[6].chain8.inv_chain[47] ;
 wire \thechain[6].chain8.inv_chain[48] ;
 wire \thechain[6].chain8.inv_chain[49] ;
 wire \thechain[6].chain8.inv_chain[4] ;
 wire \thechain[6].chain8.inv_chain[50] ;
 wire \thechain[6].chain8.inv_chain[51] ;
 wire \thechain[6].chain8.inv_chain[52] ;
 wire \thechain[6].chain8.inv_chain[53] ;
 wire \thechain[6].chain8.inv_chain[54] ;
 wire \thechain[6].chain8.inv_chain[55] ;
 wire \thechain[6].chain8.inv_chain[56] ;
 wire \thechain[6].chain8.inv_chain[57] ;
 wire \thechain[6].chain8.inv_chain[58] ;
 wire \thechain[6].chain8.inv_chain[59] ;
 wire \thechain[6].chain8.inv_chain[5] ;
 wire \thechain[6].chain8.inv_chain[60] ;
 wire \thechain[6].chain8.inv_chain[61] ;
 wire \thechain[6].chain8.inv_chain[62] ;
 wire \thechain[6].chain8.inv_chain[63] ;
 wire \thechain[6].chain8.inv_chain[64] ;
 wire \thechain[6].chain8.inv_chain[65] ;
 wire \thechain[6].chain8.inv_chain[66] ;
 wire \thechain[6].chain8.inv_chain[67] ;
 wire \thechain[6].chain8.inv_chain[68] ;
 wire \thechain[6].chain8.inv_chain[69] ;
 wire \thechain[6].chain8.inv_chain[6] ;
 wire \thechain[6].chain8.inv_chain[70] ;
 wire \thechain[6].chain8.inv_chain[71] ;
 wire \thechain[6].chain8.inv_chain[72] ;
 wire \thechain[6].chain8.inv_chain[73] ;
 wire \thechain[6].chain8.inv_chain[74] ;
 wire \thechain[6].chain8.inv_chain[75] ;
 wire \thechain[6].chain8.inv_chain[76] ;
 wire \thechain[6].chain8.inv_chain[77] ;
 wire \thechain[6].chain8.inv_chain[78] ;
 wire \thechain[6].chain8.inv_chain[79] ;
 wire \thechain[6].chain8.inv_chain[7] ;
 wire \thechain[6].chain8.inv_chain[80] ;
 wire \thechain[6].chain8.inv_chain[81] ;
 wire \thechain[6].chain8.inv_chain[82] ;
 wire \thechain[6].chain8.inv_chain[83] ;
 wire \thechain[6].chain8.inv_chain[84] ;
 wire \thechain[6].chain8.inv_chain[85] ;
 wire \thechain[6].chain8.inv_chain[86] ;
 wire \thechain[6].chain8.inv_chain[87] ;
 wire \thechain[6].chain8.inv_chain[88] ;
 wire \thechain[6].chain8.inv_chain[89] ;
 wire \thechain[6].chain8.inv_chain[8] ;
 wire \thechain[6].chain8.inv_chain[90] ;
 wire \thechain[6].chain8.inv_chain[91] ;
 wire \thechain[6].chain8.inv_chain[92] ;
 wire \thechain[6].chain8.inv_chain[93] ;
 wire \thechain[6].chain8.inv_chain[94] ;
 wire \thechain[6].chain8.inv_chain[95] ;
 wire \thechain[6].chain8.inv_chain[96] ;
 wire \thechain[6].chain8.inv_chain[97] ;
 wire \thechain[6].chain8.inv_chain[98] ;
 wire \thechain[6].chain8.inv_chain[99] ;
 wire \thechain[6].chain8.inv_chain[9] ;
 wire \thechain[6].chain9.dout ;
 wire \thechain[6].chain9.inv_chain[0] ;
 wire \thechain[6].chain9.inv_chain[100] ;
 wire \thechain[6].chain9.inv_chain[101] ;
 wire \thechain[6].chain9.inv_chain[102] ;
 wire \thechain[6].chain9.inv_chain[103] ;
 wire \thechain[6].chain9.inv_chain[104] ;
 wire \thechain[6].chain9.inv_chain[105] ;
 wire \thechain[6].chain9.inv_chain[106] ;
 wire \thechain[6].chain9.inv_chain[107] ;
 wire \thechain[6].chain9.inv_chain[108] ;
 wire \thechain[6].chain9.inv_chain[109] ;
 wire \thechain[6].chain9.inv_chain[10] ;
 wire \thechain[6].chain9.inv_chain[110] ;
 wire \thechain[6].chain9.inv_chain[111] ;
 wire \thechain[6].chain9.inv_chain[112] ;
 wire \thechain[6].chain9.inv_chain[113] ;
 wire \thechain[6].chain9.inv_chain[114] ;
 wire \thechain[6].chain9.inv_chain[115] ;
 wire \thechain[6].chain9.inv_chain[116] ;
 wire \thechain[6].chain9.inv_chain[117] ;
 wire \thechain[6].chain9.inv_chain[118] ;
 wire \thechain[6].chain9.inv_chain[119] ;
 wire \thechain[6].chain9.inv_chain[11] ;
 wire \thechain[6].chain9.inv_chain[120] ;
 wire \thechain[6].chain9.inv_chain[121] ;
 wire \thechain[6].chain9.inv_chain[122] ;
 wire \thechain[6].chain9.inv_chain[123] ;
 wire \thechain[6].chain9.inv_chain[124] ;
 wire \thechain[6].chain9.inv_chain[125] ;
 wire \thechain[6].chain9.inv_chain[126] ;
 wire \thechain[6].chain9.inv_chain[127] ;
 wire \thechain[6].chain9.inv_chain[128] ;
 wire \thechain[6].chain9.inv_chain[129] ;
 wire \thechain[6].chain9.inv_chain[12] ;
 wire \thechain[6].chain9.inv_chain[130] ;
 wire \thechain[6].chain9.inv_chain[131] ;
 wire \thechain[6].chain9.inv_chain[132] ;
 wire \thechain[6].chain9.inv_chain[133] ;
 wire \thechain[6].chain9.inv_chain[134] ;
 wire \thechain[6].chain9.inv_chain[135] ;
 wire \thechain[6].chain9.inv_chain[136] ;
 wire \thechain[6].chain9.inv_chain[137] ;
 wire \thechain[6].chain9.inv_chain[138] ;
 wire \thechain[6].chain9.inv_chain[139] ;
 wire \thechain[6].chain9.inv_chain[13] ;
 wire \thechain[6].chain9.inv_chain[140] ;
 wire \thechain[6].chain9.inv_chain[141] ;
 wire \thechain[6].chain9.inv_chain[142] ;
 wire \thechain[6].chain9.inv_chain[143] ;
 wire \thechain[6].chain9.inv_chain[144] ;
 wire \thechain[6].chain9.inv_chain[145] ;
 wire \thechain[6].chain9.inv_chain[146] ;
 wire \thechain[6].chain9.inv_chain[147] ;
 wire \thechain[6].chain9.inv_chain[148] ;
 wire \thechain[6].chain9.inv_chain[149] ;
 wire \thechain[6].chain9.inv_chain[14] ;
 wire \thechain[6].chain9.inv_chain[150] ;
 wire \thechain[6].chain9.inv_chain[151] ;
 wire \thechain[6].chain9.inv_chain[152] ;
 wire \thechain[6].chain9.inv_chain[153] ;
 wire \thechain[6].chain9.inv_chain[154] ;
 wire \thechain[6].chain9.inv_chain[155] ;
 wire \thechain[6].chain9.inv_chain[156] ;
 wire \thechain[6].chain9.inv_chain[157] ;
 wire \thechain[6].chain9.inv_chain[158] ;
 wire \thechain[6].chain9.inv_chain[159] ;
 wire \thechain[6].chain9.inv_chain[15] ;
 wire \thechain[6].chain9.inv_chain[160] ;
 wire \thechain[6].chain9.inv_chain[161] ;
 wire \thechain[6].chain9.inv_chain[162] ;
 wire \thechain[6].chain9.inv_chain[163] ;
 wire \thechain[6].chain9.inv_chain[164] ;
 wire \thechain[6].chain9.inv_chain[165] ;
 wire \thechain[6].chain9.inv_chain[166] ;
 wire \thechain[6].chain9.inv_chain[167] ;
 wire \thechain[6].chain9.inv_chain[168] ;
 wire \thechain[6].chain9.inv_chain[169] ;
 wire \thechain[6].chain9.inv_chain[16] ;
 wire \thechain[6].chain9.inv_chain[170] ;
 wire \thechain[6].chain9.inv_chain[171] ;
 wire \thechain[6].chain9.inv_chain[172] ;
 wire \thechain[6].chain9.inv_chain[173] ;
 wire \thechain[6].chain9.inv_chain[174] ;
 wire \thechain[6].chain9.inv_chain[175] ;
 wire \thechain[6].chain9.inv_chain[176] ;
 wire \thechain[6].chain9.inv_chain[177] ;
 wire \thechain[6].chain9.inv_chain[178] ;
 wire \thechain[6].chain9.inv_chain[179] ;
 wire \thechain[6].chain9.inv_chain[17] ;
 wire \thechain[6].chain9.inv_chain[180] ;
 wire \thechain[6].chain9.inv_chain[181] ;
 wire \thechain[6].chain9.inv_chain[182] ;
 wire \thechain[6].chain9.inv_chain[183] ;
 wire \thechain[6].chain9.inv_chain[184] ;
 wire \thechain[6].chain9.inv_chain[185] ;
 wire \thechain[6].chain9.inv_chain[186] ;
 wire \thechain[6].chain9.inv_chain[187] ;
 wire \thechain[6].chain9.inv_chain[188] ;
 wire \thechain[6].chain9.inv_chain[189] ;
 wire \thechain[6].chain9.inv_chain[18] ;
 wire \thechain[6].chain9.inv_chain[190] ;
 wire \thechain[6].chain9.inv_chain[191] ;
 wire \thechain[6].chain9.inv_chain[192] ;
 wire \thechain[6].chain9.inv_chain[193] ;
 wire \thechain[6].chain9.inv_chain[194] ;
 wire \thechain[6].chain9.inv_chain[195] ;
 wire \thechain[6].chain9.inv_chain[196] ;
 wire \thechain[6].chain9.inv_chain[197] ;
 wire \thechain[6].chain9.inv_chain[198] ;
 wire \thechain[6].chain9.inv_chain[199] ;
 wire \thechain[6].chain9.inv_chain[19] ;
 wire \thechain[6].chain9.inv_chain[1] ;
 wire \thechain[6].chain9.inv_chain[200] ;
 wire \thechain[6].chain9.inv_chain[201] ;
 wire \thechain[6].chain9.inv_chain[202] ;
 wire \thechain[6].chain9.inv_chain[203] ;
 wire \thechain[6].chain9.inv_chain[204] ;
 wire \thechain[6].chain9.inv_chain[205] ;
 wire \thechain[6].chain9.inv_chain[206] ;
 wire \thechain[6].chain9.inv_chain[207] ;
 wire \thechain[6].chain9.inv_chain[208] ;
 wire \thechain[6].chain9.inv_chain[209] ;
 wire \thechain[6].chain9.inv_chain[20] ;
 wire \thechain[6].chain9.inv_chain[210] ;
 wire \thechain[6].chain9.inv_chain[211] ;
 wire \thechain[6].chain9.inv_chain[212] ;
 wire \thechain[6].chain9.inv_chain[213] ;
 wire \thechain[6].chain9.inv_chain[214] ;
 wire \thechain[6].chain9.inv_chain[215] ;
 wire \thechain[6].chain9.inv_chain[216] ;
 wire \thechain[6].chain9.inv_chain[217] ;
 wire \thechain[6].chain9.inv_chain[218] ;
 wire \thechain[6].chain9.inv_chain[219] ;
 wire \thechain[6].chain9.inv_chain[21] ;
 wire \thechain[6].chain9.inv_chain[220] ;
 wire \thechain[6].chain9.inv_chain[221] ;
 wire \thechain[6].chain9.inv_chain[222] ;
 wire \thechain[6].chain9.inv_chain[223] ;
 wire \thechain[6].chain9.inv_chain[224] ;
 wire \thechain[6].chain9.inv_chain[225] ;
 wire \thechain[6].chain9.inv_chain[226] ;
 wire \thechain[6].chain9.inv_chain[227] ;
 wire \thechain[6].chain9.inv_chain[228] ;
 wire \thechain[6].chain9.inv_chain[229] ;
 wire \thechain[6].chain9.inv_chain[22] ;
 wire \thechain[6].chain9.inv_chain[230] ;
 wire \thechain[6].chain9.inv_chain[231] ;
 wire \thechain[6].chain9.inv_chain[232] ;
 wire \thechain[6].chain9.inv_chain[233] ;
 wire \thechain[6].chain9.inv_chain[234] ;
 wire \thechain[6].chain9.inv_chain[235] ;
 wire \thechain[6].chain9.inv_chain[236] ;
 wire \thechain[6].chain9.inv_chain[237] ;
 wire \thechain[6].chain9.inv_chain[238] ;
 wire \thechain[6].chain9.inv_chain[239] ;
 wire \thechain[6].chain9.inv_chain[23] ;
 wire \thechain[6].chain9.inv_chain[240] ;
 wire \thechain[6].chain9.inv_chain[241] ;
 wire \thechain[6].chain9.inv_chain[242] ;
 wire \thechain[6].chain9.inv_chain[243] ;
 wire \thechain[6].chain9.inv_chain[244] ;
 wire \thechain[6].chain9.inv_chain[245] ;
 wire \thechain[6].chain9.inv_chain[246] ;
 wire \thechain[6].chain9.inv_chain[247] ;
 wire \thechain[6].chain9.inv_chain[248] ;
 wire \thechain[6].chain9.inv_chain[249] ;
 wire \thechain[6].chain9.inv_chain[24] ;
 wire \thechain[6].chain9.inv_chain[250] ;
 wire \thechain[6].chain9.inv_chain[251] ;
 wire \thechain[6].chain9.inv_chain[252] ;
 wire \thechain[6].chain9.inv_chain[253] ;
 wire \thechain[6].chain9.inv_chain[254] ;
 wire \thechain[6].chain9.inv_chain[255] ;
 wire \thechain[6].chain9.inv_chain[256] ;
 wire \thechain[6].chain9.inv_chain[25] ;
 wire \thechain[6].chain9.inv_chain[26] ;
 wire \thechain[6].chain9.inv_chain[27] ;
 wire \thechain[6].chain9.inv_chain[28] ;
 wire \thechain[6].chain9.inv_chain[29] ;
 wire \thechain[6].chain9.inv_chain[2] ;
 wire \thechain[6].chain9.inv_chain[30] ;
 wire \thechain[6].chain9.inv_chain[31] ;
 wire \thechain[6].chain9.inv_chain[32] ;
 wire \thechain[6].chain9.inv_chain[33] ;
 wire \thechain[6].chain9.inv_chain[34] ;
 wire \thechain[6].chain9.inv_chain[35] ;
 wire \thechain[6].chain9.inv_chain[36] ;
 wire \thechain[6].chain9.inv_chain[37] ;
 wire \thechain[6].chain9.inv_chain[38] ;
 wire \thechain[6].chain9.inv_chain[39] ;
 wire \thechain[6].chain9.inv_chain[3] ;
 wire \thechain[6].chain9.inv_chain[40] ;
 wire \thechain[6].chain9.inv_chain[41] ;
 wire \thechain[6].chain9.inv_chain[42] ;
 wire \thechain[6].chain9.inv_chain[43] ;
 wire \thechain[6].chain9.inv_chain[44] ;
 wire \thechain[6].chain9.inv_chain[45] ;
 wire \thechain[6].chain9.inv_chain[46] ;
 wire \thechain[6].chain9.inv_chain[47] ;
 wire \thechain[6].chain9.inv_chain[48] ;
 wire \thechain[6].chain9.inv_chain[49] ;
 wire \thechain[6].chain9.inv_chain[4] ;
 wire \thechain[6].chain9.inv_chain[50] ;
 wire \thechain[6].chain9.inv_chain[51] ;
 wire \thechain[6].chain9.inv_chain[52] ;
 wire \thechain[6].chain9.inv_chain[53] ;
 wire \thechain[6].chain9.inv_chain[54] ;
 wire \thechain[6].chain9.inv_chain[55] ;
 wire \thechain[6].chain9.inv_chain[56] ;
 wire \thechain[6].chain9.inv_chain[57] ;
 wire \thechain[6].chain9.inv_chain[58] ;
 wire \thechain[6].chain9.inv_chain[59] ;
 wire \thechain[6].chain9.inv_chain[5] ;
 wire \thechain[6].chain9.inv_chain[60] ;
 wire \thechain[6].chain9.inv_chain[61] ;
 wire \thechain[6].chain9.inv_chain[62] ;
 wire \thechain[6].chain9.inv_chain[63] ;
 wire \thechain[6].chain9.inv_chain[64] ;
 wire \thechain[6].chain9.inv_chain[65] ;
 wire \thechain[6].chain9.inv_chain[66] ;
 wire \thechain[6].chain9.inv_chain[67] ;
 wire \thechain[6].chain9.inv_chain[68] ;
 wire \thechain[6].chain9.inv_chain[69] ;
 wire \thechain[6].chain9.inv_chain[6] ;
 wire \thechain[6].chain9.inv_chain[70] ;
 wire \thechain[6].chain9.inv_chain[71] ;
 wire \thechain[6].chain9.inv_chain[72] ;
 wire \thechain[6].chain9.inv_chain[73] ;
 wire \thechain[6].chain9.inv_chain[74] ;
 wire \thechain[6].chain9.inv_chain[75] ;
 wire \thechain[6].chain9.inv_chain[76] ;
 wire \thechain[6].chain9.inv_chain[77] ;
 wire \thechain[6].chain9.inv_chain[78] ;
 wire \thechain[6].chain9.inv_chain[79] ;
 wire \thechain[6].chain9.inv_chain[7] ;
 wire \thechain[6].chain9.inv_chain[80] ;
 wire \thechain[6].chain9.inv_chain[81] ;
 wire \thechain[6].chain9.inv_chain[82] ;
 wire \thechain[6].chain9.inv_chain[83] ;
 wire \thechain[6].chain9.inv_chain[84] ;
 wire \thechain[6].chain9.inv_chain[85] ;
 wire \thechain[6].chain9.inv_chain[86] ;
 wire \thechain[6].chain9.inv_chain[87] ;
 wire \thechain[6].chain9.inv_chain[88] ;
 wire \thechain[6].chain9.inv_chain[89] ;
 wire \thechain[6].chain9.inv_chain[8] ;
 wire \thechain[6].chain9.inv_chain[90] ;
 wire \thechain[6].chain9.inv_chain[91] ;
 wire \thechain[6].chain9.inv_chain[92] ;
 wire \thechain[6].chain9.inv_chain[93] ;
 wire \thechain[6].chain9.inv_chain[94] ;
 wire \thechain[6].chain9.inv_chain[95] ;
 wire \thechain[6].chain9.inv_chain[96] ;
 wire \thechain[6].chain9.inv_chain[97] ;
 wire \thechain[6].chain9.inv_chain[98] ;
 wire \thechain[6].chain9.inv_chain[99] ;
 wire \thechain[6].chain9.inv_chain[9] ;
 wire \thechain[7].chain1.dout ;
 wire \thechain[7].chain1.inv_chain[0] ;
 wire \thechain[7].chain1.inv_chain[1] ;
 wire \thechain[7].chain1.inv_chain[2] ;
 wire \thechain[7].chain2.dout ;
 wire \thechain[7].chain2.inv_chain[0] ;
 wire \thechain[7].chain2.inv_chain[1] ;
 wire \thechain[7].chain2.inv_chain[2] ;
 wire \thechain[7].chain2.inv_chain[3] ;
 wire \thechain[7].chain2.inv_chain[4] ;
 wire \thechain[7].chain3.dout ;
 wire \thechain[7].chain3.inv_chain[0] ;
 wire \thechain[7].chain3.inv_chain[1] ;
 wire \thechain[7].chain3.inv_chain[2] ;
 wire \thechain[7].chain3.inv_chain[3] ;
 wire \thechain[7].chain3.inv_chain[4] ;
 wire \thechain[7].chain3.inv_chain[5] ;
 wire \thechain[7].chain3.inv_chain[6] ;
 wire \thechain[7].chain3.inv_chain[7] ;
 wire \thechain[7].chain3.inv_chain[8] ;
 wire \thechain[7].chain4.dout ;
 wire \thechain[7].chain4.inv_chain[0] ;
 wire \thechain[7].chain4.inv_chain[10] ;
 wire \thechain[7].chain4.inv_chain[11] ;
 wire \thechain[7].chain4.inv_chain[12] ;
 wire \thechain[7].chain4.inv_chain[13] ;
 wire \thechain[7].chain4.inv_chain[14] ;
 wire \thechain[7].chain4.inv_chain[15] ;
 wire \thechain[7].chain4.inv_chain[16] ;
 wire \thechain[7].chain4.inv_chain[1] ;
 wire \thechain[7].chain4.inv_chain[2] ;
 wire \thechain[7].chain4.inv_chain[3] ;
 wire \thechain[7].chain4.inv_chain[4] ;
 wire \thechain[7].chain4.inv_chain[5] ;
 wire \thechain[7].chain4.inv_chain[6] ;
 wire \thechain[7].chain4.inv_chain[7] ;
 wire \thechain[7].chain4.inv_chain[8] ;
 wire \thechain[7].chain4.inv_chain[9] ;
 wire \thechain[7].chain5.dout ;
 wire \thechain[7].chain5.inv_chain[0] ;
 wire \thechain[7].chain5.inv_chain[10] ;
 wire \thechain[7].chain5.inv_chain[11] ;
 wire \thechain[7].chain5.inv_chain[12] ;
 wire \thechain[7].chain5.inv_chain[13] ;
 wire \thechain[7].chain5.inv_chain[14] ;
 wire \thechain[7].chain5.inv_chain[15] ;
 wire \thechain[7].chain5.inv_chain[16] ;
 wire \thechain[7].chain5.inv_chain[17] ;
 wire \thechain[7].chain5.inv_chain[18] ;
 wire \thechain[7].chain5.inv_chain[19] ;
 wire \thechain[7].chain5.inv_chain[1] ;
 wire \thechain[7].chain5.inv_chain[20] ;
 wire \thechain[7].chain5.inv_chain[21] ;
 wire \thechain[7].chain5.inv_chain[22] ;
 wire \thechain[7].chain5.inv_chain[23] ;
 wire \thechain[7].chain5.inv_chain[24] ;
 wire \thechain[7].chain5.inv_chain[25] ;
 wire \thechain[7].chain5.inv_chain[26] ;
 wire \thechain[7].chain5.inv_chain[27] ;
 wire \thechain[7].chain5.inv_chain[28] ;
 wire \thechain[7].chain5.inv_chain[29] ;
 wire \thechain[7].chain5.inv_chain[2] ;
 wire \thechain[7].chain5.inv_chain[30] ;
 wire \thechain[7].chain5.inv_chain[31] ;
 wire \thechain[7].chain5.inv_chain[32] ;
 wire \thechain[7].chain5.inv_chain[3] ;
 wire \thechain[7].chain5.inv_chain[4] ;
 wire \thechain[7].chain5.inv_chain[5] ;
 wire \thechain[7].chain5.inv_chain[6] ;
 wire \thechain[7].chain5.inv_chain[7] ;
 wire \thechain[7].chain5.inv_chain[8] ;
 wire \thechain[7].chain5.inv_chain[9] ;
 wire \thechain[7].chain6.dout ;
 wire \thechain[7].chain6.inv_chain[0] ;
 wire \thechain[7].chain6.inv_chain[10] ;
 wire \thechain[7].chain6.inv_chain[11] ;
 wire \thechain[7].chain6.inv_chain[12] ;
 wire \thechain[7].chain6.inv_chain[13] ;
 wire \thechain[7].chain6.inv_chain[14] ;
 wire \thechain[7].chain6.inv_chain[15] ;
 wire \thechain[7].chain6.inv_chain[16] ;
 wire \thechain[7].chain6.inv_chain[17] ;
 wire \thechain[7].chain6.inv_chain[18] ;
 wire \thechain[7].chain6.inv_chain[19] ;
 wire \thechain[7].chain6.inv_chain[1] ;
 wire \thechain[7].chain6.inv_chain[20] ;
 wire \thechain[7].chain6.inv_chain[21] ;
 wire \thechain[7].chain6.inv_chain[22] ;
 wire \thechain[7].chain6.inv_chain[23] ;
 wire \thechain[7].chain6.inv_chain[24] ;
 wire \thechain[7].chain6.inv_chain[25] ;
 wire \thechain[7].chain6.inv_chain[26] ;
 wire \thechain[7].chain6.inv_chain[27] ;
 wire \thechain[7].chain6.inv_chain[28] ;
 wire \thechain[7].chain6.inv_chain[29] ;
 wire \thechain[7].chain6.inv_chain[2] ;
 wire \thechain[7].chain6.inv_chain[30] ;
 wire \thechain[7].chain6.inv_chain[31] ;
 wire \thechain[7].chain6.inv_chain[32] ;
 wire \thechain[7].chain6.inv_chain[33] ;
 wire \thechain[7].chain6.inv_chain[34] ;
 wire \thechain[7].chain6.inv_chain[35] ;
 wire \thechain[7].chain6.inv_chain[36] ;
 wire \thechain[7].chain6.inv_chain[37] ;
 wire \thechain[7].chain6.inv_chain[38] ;
 wire \thechain[7].chain6.inv_chain[39] ;
 wire \thechain[7].chain6.inv_chain[3] ;
 wire \thechain[7].chain6.inv_chain[40] ;
 wire \thechain[7].chain6.inv_chain[41] ;
 wire \thechain[7].chain6.inv_chain[42] ;
 wire \thechain[7].chain6.inv_chain[43] ;
 wire \thechain[7].chain6.inv_chain[44] ;
 wire \thechain[7].chain6.inv_chain[45] ;
 wire \thechain[7].chain6.inv_chain[46] ;
 wire \thechain[7].chain6.inv_chain[47] ;
 wire \thechain[7].chain6.inv_chain[48] ;
 wire \thechain[7].chain6.inv_chain[49] ;
 wire \thechain[7].chain6.inv_chain[4] ;
 wire \thechain[7].chain6.inv_chain[50] ;
 wire \thechain[7].chain6.inv_chain[51] ;
 wire \thechain[7].chain6.inv_chain[52] ;
 wire \thechain[7].chain6.inv_chain[53] ;
 wire \thechain[7].chain6.inv_chain[54] ;
 wire \thechain[7].chain6.inv_chain[55] ;
 wire \thechain[7].chain6.inv_chain[56] ;
 wire \thechain[7].chain6.inv_chain[57] ;
 wire \thechain[7].chain6.inv_chain[58] ;
 wire \thechain[7].chain6.inv_chain[59] ;
 wire \thechain[7].chain6.inv_chain[5] ;
 wire \thechain[7].chain6.inv_chain[60] ;
 wire \thechain[7].chain6.inv_chain[61] ;
 wire \thechain[7].chain6.inv_chain[62] ;
 wire \thechain[7].chain6.inv_chain[63] ;
 wire \thechain[7].chain6.inv_chain[64] ;
 wire \thechain[7].chain6.inv_chain[6] ;
 wire \thechain[7].chain6.inv_chain[7] ;
 wire \thechain[7].chain6.inv_chain[8] ;
 wire \thechain[7].chain6.inv_chain[9] ;
 wire \thechain[7].chain7.dout ;
 wire \thechain[7].chain7.inv_chain[0] ;
 wire \thechain[7].chain7.inv_chain[100] ;
 wire \thechain[7].chain7.inv_chain[101] ;
 wire \thechain[7].chain7.inv_chain[102] ;
 wire \thechain[7].chain7.inv_chain[103] ;
 wire \thechain[7].chain7.inv_chain[104] ;
 wire \thechain[7].chain7.inv_chain[105] ;
 wire \thechain[7].chain7.inv_chain[106] ;
 wire \thechain[7].chain7.inv_chain[107] ;
 wire \thechain[7].chain7.inv_chain[108] ;
 wire \thechain[7].chain7.inv_chain[109] ;
 wire \thechain[7].chain7.inv_chain[10] ;
 wire \thechain[7].chain7.inv_chain[110] ;
 wire \thechain[7].chain7.inv_chain[111] ;
 wire \thechain[7].chain7.inv_chain[112] ;
 wire \thechain[7].chain7.inv_chain[113] ;
 wire \thechain[7].chain7.inv_chain[114] ;
 wire \thechain[7].chain7.inv_chain[115] ;
 wire \thechain[7].chain7.inv_chain[116] ;
 wire \thechain[7].chain7.inv_chain[117] ;
 wire \thechain[7].chain7.inv_chain[118] ;
 wire \thechain[7].chain7.inv_chain[119] ;
 wire \thechain[7].chain7.inv_chain[11] ;
 wire \thechain[7].chain7.inv_chain[120] ;
 wire \thechain[7].chain7.inv_chain[121] ;
 wire \thechain[7].chain7.inv_chain[122] ;
 wire \thechain[7].chain7.inv_chain[123] ;
 wire \thechain[7].chain7.inv_chain[124] ;
 wire \thechain[7].chain7.inv_chain[125] ;
 wire \thechain[7].chain7.inv_chain[126] ;
 wire \thechain[7].chain7.inv_chain[127] ;
 wire \thechain[7].chain7.inv_chain[128] ;
 wire \thechain[7].chain7.inv_chain[12] ;
 wire \thechain[7].chain7.inv_chain[13] ;
 wire \thechain[7].chain7.inv_chain[14] ;
 wire \thechain[7].chain7.inv_chain[15] ;
 wire \thechain[7].chain7.inv_chain[16] ;
 wire \thechain[7].chain7.inv_chain[17] ;
 wire \thechain[7].chain7.inv_chain[18] ;
 wire \thechain[7].chain7.inv_chain[19] ;
 wire \thechain[7].chain7.inv_chain[1] ;
 wire \thechain[7].chain7.inv_chain[20] ;
 wire \thechain[7].chain7.inv_chain[21] ;
 wire \thechain[7].chain7.inv_chain[22] ;
 wire \thechain[7].chain7.inv_chain[23] ;
 wire \thechain[7].chain7.inv_chain[24] ;
 wire \thechain[7].chain7.inv_chain[25] ;
 wire \thechain[7].chain7.inv_chain[26] ;
 wire \thechain[7].chain7.inv_chain[27] ;
 wire \thechain[7].chain7.inv_chain[28] ;
 wire \thechain[7].chain7.inv_chain[29] ;
 wire \thechain[7].chain7.inv_chain[2] ;
 wire \thechain[7].chain7.inv_chain[30] ;
 wire \thechain[7].chain7.inv_chain[31] ;
 wire \thechain[7].chain7.inv_chain[32] ;
 wire \thechain[7].chain7.inv_chain[33] ;
 wire \thechain[7].chain7.inv_chain[34] ;
 wire \thechain[7].chain7.inv_chain[35] ;
 wire \thechain[7].chain7.inv_chain[36] ;
 wire \thechain[7].chain7.inv_chain[37] ;
 wire \thechain[7].chain7.inv_chain[38] ;
 wire \thechain[7].chain7.inv_chain[39] ;
 wire \thechain[7].chain7.inv_chain[3] ;
 wire \thechain[7].chain7.inv_chain[40] ;
 wire \thechain[7].chain7.inv_chain[41] ;
 wire \thechain[7].chain7.inv_chain[42] ;
 wire \thechain[7].chain7.inv_chain[43] ;
 wire \thechain[7].chain7.inv_chain[44] ;
 wire \thechain[7].chain7.inv_chain[45] ;
 wire \thechain[7].chain7.inv_chain[46] ;
 wire \thechain[7].chain7.inv_chain[47] ;
 wire \thechain[7].chain7.inv_chain[48] ;
 wire \thechain[7].chain7.inv_chain[49] ;
 wire \thechain[7].chain7.inv_chain[4] ;
 wire \thechain[7].chain7.inv_chain[50] ;
 wire \thechain[7].chain7.inv_chain[51] ;
 wire \thechain[7].chain7.inv_chain[52] ;
 wire \thechain[7].chain7.inv_chain[53] ;
 wire \thechain[7].chain7.inv_chain[54] ;
 wire \thechain[7].chain7.inv_chain[55] ;
 wire \thechain[7].chain7.inv_chain[56] ;
 wire \thechain[7].chain7.inv_chain[57] ;
 wire \thechain[7].chain7.inv_chain[58] ;
 wire \thechain[7].chain7.inv_chain[59] ;
 wire \thechain[7].chain7.inv_chain[5] ;
 wire \thechain[7].chain7.inv_chain[60] ;
 wire \thechain[7].chain7.inv_chain[61] ;
 wire \thechain[7].chain7.inv_chain[62] ;
 wire \thechain[7].chain7.inv_chain[63] ;
 wire \thechain[7].chain7.inv_chain[64] ;
 wire \thechain[7].chain7.inv_chain[65] ;
 wire \thechain[7].chain7.inv_chain[66] ;
 wire \thechain[7].chain7.inv_chain[67] ;
 wire \thechain[7].chain7.inv_chain[68] ;
 wire \thechain[7].chain7.inv_chain[69] ;
 wire \thechain[7].chain7.inv_chain[6] ;
 wire \thechain[7].chain7.inv_chain[70] ;
 wire \thechain[7].chain7.inv_chain[71] ;
 wire \thechain[7].chain7.inv_chain[72] ;
 wire \thechain[7].chain7.inv_chain[73] ;
 wire \thechain[7].chain7.inv_chain[74] ;
 wire \thechain[7].chain7.inv_chain[75] ;
 wire \thechain[7].chain7.inv_chain[76] ;
 wire \thechain[7].chain7.inv_chain[77] ;
 wire \thechain[7].chain7.inv_chain[78] ;
 wire \thechain[7].chain7.inv_chain[79] ;
 wire \thechain[7].chain7.inv_chain[7] ;
 wire \thechain[7].chain7.inv_chain[80] ;
 wire \thechain[7].chain7.inv_chain[81] ;
 wire \thechain[7].chain7.inv_chain[82] ;
 wire \thechain[7].chain7.inv_chain[83] ;
 wire \thechain[7].chain7.inv_chain[84] ;
 wire \thechain[7].chain7.inv_chain[85] ;
 wire \thechain[7].chain7.inv_chain[86] ;
 wire \thechain[7].chain7.inv_chain[87] ;
 wire \thechain[7].chain7.inv_chain[88] ;
 wire \thechain[7].chain7.inv_chain[89] ;
 wire \thechain[7].chain7.inv_chain[8] ;
 wire \thechain[7].chain7.inv_chain[90] ;
 wire \thechain[7].chain7.inv_chain[91] ;
 wire \thechain[7].chain7.inv_chain[92] ;
 wire \thechain[7].chain7.inv_chain[93] ;
 wire \thechain[7].chain7.inv_chain[94] ;
 wire \thechain[7].chain7.inv_chain[95] ;
 wire \thechain[7].chain7.inv_chain[96] ;
 wire \thechain[7].chain7.inv_chain[97] ;
 wire \thechain[7].chain7.inv_chain[98] ;
 wire \thechain[7].chain7.inv_chain[99] ;
 wire \thechain[7].chain7.inv_chain[9] ;
 wire \thechain[7].chain8.dout ;
 wire \thechain[7].chain8.inv_chain[0] ;
 wire \thechain[7].chain8.inv_chain[100] ;
 wire \thechain[7].chain8.inv_chain[101] ;
 wire \thechain[7].chain8.inv_chain[102] ;
 wire \thechain[7].chain8.inv_chain[103] ;
 wire \thechain[7].chain8.inv_chain[104] ;
 wire \thechain[7].chain8.inv_chain[105] ;
 wire \thechain[7].chain8.inv_chain[106] ;
 wire \thechain[7].chain8.inv_chain[107] ;
 wire \thechain[7].chain8.inv_chain[108] ;
 wire \thechain[7].chain8.inv_chain[109] ;
 wire \thechain[7].chain8.inv_chain[10] ;
 wire \thechain[7].chain8.inv_chain[110] ;
 wire \thechain[7].chain8.inv_chain[111] ;
 wire \thechain[7].chain8.inv_chain[112] ;
 wire \thechain[7].chain8.inv_chain[113] ;
 wire \thechain[7].chain8.inv_chain[114] ;
 wire \thechain[7].chain8.inv_chain[115] ;
 wire \thechain[7].chain8.inv_chain[116] ;
 wire \thechain[7].chain8.inv_chain[117] ;
 wire \thechain[7].chain8.inv_chain[118] ;
 wire \thechain[7].chain8.inv_chain[119] ;
 wire \thechain[7].chain8.inv_chain[11] ;
 wire \thechain[7].chain8.inv_chain[120] ;
 wire \thechain[7].chain8.inv_chain[121] ;
 wire \thechain[7].chain8.inv_chain[122] ;
 wire \thechain[7].chain8.inv_chain[123] ;
 wire \thechain[7].chain8.inv_chain[124] ;
 wire \thechain[7].chain8.inv_chain[125] ;
 wire \thechain[7].chain8.inv_chain[126] ;
 wire \thechain[7].chain8.inv_chain[127] ;
 wire \thechain[7].chain8.inv_chain[128] ;
 wire \thechain[7].chain8.inv_chain[129] ;
 wire \thechain[7].chain8.inv_chain[12] ;
 wire \thechain[7].chain8.inv_chain[130] ;
 wire \thechain[7].chain8.inv_chain[131] ;
 wire \thechain[7].chain8.inv_chain[132] ;
 wire \thechain[7].chain8.inv_chain[133] ;
 wire \thechain[7].chain8.inv_chain[134] ;
 wire \thechain[7].chain8.inv_chain[135] ;
 wire \thechain[7].chain8.inv_chain[136] ;
 wire \thechain[7].chain8.inv_chain[137] ;
 wire \thechain[7].chain8.inv_chain[138] ;
 wire \thechain[7].chain8.inv_chain[139] ;
 wire \thechain[7].chain8.inv_chain[13] ;
 wire \thechain[7].chain8.inv_chain[140] ;
 wire \thechain[7].chain8.inv_chain[141] ;
 wire \thechain[7].chain8.inv_chain[142] ;
 wire \thechain[7].chain8.inv_chain[143] ;
 wire \thechain[7].chain8.inv_chain[144] ;
 wire \thechain[7].chain8.inv_chain[145] ;
 wire \thechain[7].chain8.inv_chain[146] ;
 wire \thechain[7].chain8.inv_chain[147] ;
 wire \thechain[7].chain8.inv_chain[148] ;
 wire \thechain[7].chain8.inv_chain[149] ;
 wire \thechain[7].chain8.inv_chain[14] ;
 wire \thechain[7].chain8.inv_chain[150] ;
 wire \thechain[7].chain8.inv_chain[151] ;
 wire \thechain[7].chain8.inv_chain[152] ;
 wire \thechain[7].chain8.inv_chain[153] ;
 wire \thechain[7].chain8.inv_chain[154] ;
 wire \thechain[7].chain8.inv_chain[155] ;
 wire \thechain[7].chain8.inv_chain[156] ;
 wire \thechain[7].chain8.inv_chain[157] ;
 wire \thechain[7].chain8.inv_chain[158] ;
 wire \thechain[7].chain8.inv_chain[159] ;
 wire \thechain[7].chain8.inv_chain[15] ;
 wire \thechain[7].chain8.inv_chain[160] ;
 wire \thechain[7].chain8.inv_chain[161] ;
 wire \thechain[7].chain8.inv_chain[162] ;
 wire \thechain[7].chain8.inv_chain[163] ;
 wire \thechain[7].chain8.inv_chain[164] ;
 wire \thechain[7].chain8.inv_chain[165] ;
 wire \thechain[7].chain8.inv_chain[166] ;
 wire \thechain[7].chain8.inv_chain[167] ;
 wire \thechain[7].chain8.inv_chain[168] ;
 wire \thechain[7].chain8.inv_chain[169] ;
 wire \thechain[7].chain8.inv_chain[16] ;
 wire \thechain[7].chain8.inv_chain[170] ;
 wire \thechain[7].chain8.inv_chain[171] ;
 wire \thechain[7].chain8.inv_chain[172] ;
 wire \thechain[7].chain8.inv_chain[173] ;
 wire \thechain[7].chain8.inv_chain[174] ;
 wire \thechain[7].chain8.inv_chain[175] ;
 wire \thechain[7].chain8.inv_chain[176] ;
 wire \thechain[7].chain8.inv_chain[177] ;
 wire \thechain[7].chain8.inv_chain[178] ;
 wire \thechain[7].chain8.inv_chain[179] ;
 wire \thechain[7].chain8.inv_chain[17] ;
 wire \thechain[7].chain8.inv_chain[180] ;
 wire \thechain[7].chain8.inv_chain[181] ;
 wire \thechain[7].chain8.inv_chain[182] ;
 wire \thechain[7].chain8.inv_chain[183] ;
 wire \thechain[7].chain8.inv_chain[184] ;
 wire \thechain[7].chain8.inv_chain[185] ;
 wire \thechain[7].chain8.inv_chain[186] ;
 wire \thechain[7].chain8.inv_chain[187] ;
 wire \thechain[7].chain8.inv_chain[188] ;
 wire \thechain[7].chain8.inv_chain[189] ;
 wire \thechain[7].chain8.inv_chain[18] ;
 wire \thechain[7].chain8.inv_chain[190] ;
 wire \thechain[7].chain8.inv_chain[191] ;
 wire \thechain[7].chain8.inv_chain[192] ;
 wire \thechain[7].chain8.inv_chain[19] ;
 wire \thechain[7].chain8.inv_chain[1] ;
 wire \thechain[7].chain8.inv_chain[20] ;
 wire \thechain[7].chain8.inv_chain[21] ;
 wire \thechain[7].chain8.inv_chain[22] ;
 wire \thechain[7].chain8.inv_chain[23] ;
 wire \thechain[7].chain8.inv_chain[24] ;
 wire \thechain[7].chain8.inv_chain[25] ;
 wire \thechain[7].chain8.inv_chain[26] ;
 wire \thechain[7].chain8.inv_chain[27] ;
 wire \thechain[7].chain8.inv_chain[28] ;
 wire \thechain[7].chain8.inv_chain[29] ;
 wire \thechain[7].chain8.inv_chain[2] ;
 wire \thechain[7].chain8.inv_chain[30] ;
 wire \thechain[7].chain8.inv_chain[31] ;
 wire \thechain[7].chain8.inv_chain[32] ;
 wire \thechain[7].chain8.inv_chain[33] ;
 wire \thechain[7].chain8.inv_chain[34] ;
 wire \thechain[7].chain8.inv_chain[35] ;
 wire \thechain[7].chain8.inv_chain[36] ;
 wire \thechain[7].chain8.inv_chain[37] ;
 wire \thechain[7].chain8.inv_chain[38] ;
 wire \thechain[7].chain8.inv_chain[39] ;
 wire \thechain[7].chain8.inv_chain[3] ;
 wire \thechain[7].chain8.inv_chain[40] ;
 wire \thechain[7].chain8.inv_chain[41] ;
 wire \thechain[7].chain8.inv_chain[42] ;
 wire \thechain[7].chain8.inv_chain[43] ;
 wire \thechain[7].chain8.inv_chain[44] ;
 wire \thechain[7].chain8.inv_chain[45] ;
 wire \thechain[7].chain8.inv_chain[46] ;
 wire \thechain[7].chain8.inv_chain[47] ;
 wire \thechain[7].chain8.inv_chain[48] ;
 wire \thechain[7].chain8.inv_chain[49] ;
 wire \thechain[7].chain8.inv_chain[4] ;
 wire \thechain[7].chain8.inv_chain[50] ;
 wire \thechain[7].chain8.inv_chain[51] ;
 wire \thechain[7].chain8.inv_chain[52] ;
 wire \thechain[7].chain8.inv_chain[53] ;
 wire \thechain[7].chain8.inv_chain[54] ;
 wire \thechain[7].chain8.inv_chain[55] ;
 wire \thechain[7].chain8.inv_chain[56] ;
 wire \thechain[7].chain8.inv_chain[57] ;
 wire \thechain[7].chain8.inv_chain[58] ;
 wire \thechain[7].chain8.inv_chain[59] ;
 wire \thechain[7].chain8.inv_chain[5] ;
 wire \thechain[7].chain8.inv_chain[60] ;
 wire \thechain[7].chain8.inv_chain[61] ;
 wire \thechain[7].chain8.inv_chain[62] ;
 wire \thechain[7].chain8.inv_chain[63] ;
 wire \thechain[7].chain8.inv_chain[64] ;
 wire \thechain[7].chain8.inv_chain[65] ;
 wire \thechain[7].chain8.inv_chain[66] ;
 wire \thechain[7].chain8.inv_chain[67] ;
 wire \thechain[7].chain8.inv_chain[68] ;
 wire \thechain[7].chain8.inv_chain[69] ;
 wire \thechain[7].chain8.inv_chain[6] ;
 wire \thechain[7].chain8.inv_chain[70] ;
 wire \thechain[7].chain8.inv_chain[71] ;
 wire \thechain[7].chain8.inv_chain[72] ;
 wire \thechain[7].chain8.inv_chain[73] ;
 wire \thechain[7].chain8.inv_chain[74] ;
 wire \thechain[7].chain8.inv_chain[75] ;
 wire \thechain[7].chain8.inv_chain[76] ;
 wire \thechain[7].chain8.inv_chain[77] ;
 wire \thechain[7].chain8.inv_chain[78] ;
 wire \thechain[7].chain8.inv_chain[79] ;
 wire \thechain[7].chain8.inv_chain[7] ;
 wire \thechain[7].chain8.inv_chain[80] ;
 wire \thechain[7].chain8.inv_chain[81] ;
 wire \thechain[7].chain8.inv_chain[82] ;
 wire \thechain[7].chain8.inv_chain[83] ;
 wire \thechain[7].chain8.inv_chain[84] ;
 wire \thechain[7].chain8.inv_chain[85] ;
 wire \thechain[7].chain8.inv_chain[86] ;
 wire \thechain[7].chain8.inv_chain[87] ;
 wire \thechain[7].chain8.inv_chain[88] ;
 wire \thechain[7].chain8.inv_chain[89] ;
 wire \thechain[7].chain8.inv_chain[8] ;
 wire \thechain[7].chain8.inv_chain[90] ;
 wire \thechain[7].chain8.inv_chain[91] ;
 wire \thechain[7].chain8.inv_chain[92] ;
 wire \thechain[7].chain8.inv_chain[93] ;
 wire \thechain[7].chain8.inv_chain[94] ;
 wire \thechain[7].chain8.inv_chain[95] ;
 wire \thechain[7].chain8.inv_chain[96] ;
 wire \thechain[7].chain8.inv_chain[97] ;
 wire \thechain[7].chain8.inv_chain[98] ;
 wire \thechain[7].chain8.inv_chain[99] ;
 wire \thechain[7].chain8.inv_chain[9] ;
 wire \thechain[7].chain9.dout ;
 wire \thechain[7].chain9.inv_chain[0] ;
 wire \thechain[7].chain9.inv_chain[100] ;
 wire \thechain[7].chain9.inv_chain[101] ;
 wire \thechain[7].chain9.inv_chain[102] ;
 wire \thechain[7].chain9.inv_chain[103] ;
 wire \thechain[7].chain9.inv_chain[104] ;
 wire \thechain[7].chain9.inv_chain[105] ;
 wire \thechain[7].chain9.inv_chain[106] ;
 wire \thechain[7].chain9.inv_chain[107] ;
 wire \thechain[7].chain9.inv_chain[108] ;
 wire \thechain[7].chain9.inv_chain[109] ;
 wire \thechain[7].chain9.inv_chain[10] ;
 wire \thechain[7].chain9.inv_chain[110] ;
 wire \thechain[7].chain9.inv_chain[111] ;
 wire \thechain[7].chain9.inv_chain[112] ;
 wire \thechain[7].chain9.inv_chain[113] ;
 wire \thechain[7].chain9.inv_chain[114] ;
 wire \thechain[7].chain9.inv_chain[115] ;
 wire \thechain[7].chain9.inv_chain[116] ;
 wire \thechain[7].chain9.inv_chain[117] ;
 wire \thechain[7].chain9.inv_chain[118] ;
 wire \thechain[7].chain9.inv_chain[119] ;
 wire \thechain[7].chain9.inv_chain[11] ;
 wire \thechain[7].chain9.inv_chain[120] ;
 wire \thechain[7].chain9.inv_chain[121] ;
 wire \thechain[7].chain9.inv_chain[122] ;
 wire \thechain[7].chain9.inv_chain[123] ;
 wire \thechain[7].chain9.inv_chain[124] ;
 wire \thechain[7].chain9.inv_chain[125] ;
 wire \thechain[7].chain9.inv_chain[126] ;
 wire \thechain[7].chain9.inv_chain[127] ;
 wire \thechain[7].chain9.inv_chain[128] ;
 wire \thechain[7].chain9.inv_chain[129] ;
 wire \thechain[7].chain9.inv_chain[12] ;
 wire \thechain[7].chain9.inv_chain[130] ;
 wire \thechain[7].chain9.inv_chain[131] ;
 wire \thechain[7].chain9.inv_chain[132] ;
 wire \thechain[7].chain9.inv_chain[133] ;
 wire \thechain[7].chain9.inv_chain[134] ;
 wire \thechain[7].chain9.inv_chain[135] ;
 wire \thechain[7].chain9.inv_chain[136] ;
 wire \thechain[7].chain9.inv_chain[137] ;
 wire \thechain[7].chain9.inv_chain[138] ;
 wire \thechain[7].chain9.inv_chain[139] ;
 wire \thechain[7].chain9.inv_chain[13] ;
 wire \thechain[7].chain9.inv_chain[140] ;
 wire \thechain[7].chain9.inv_chain[141] ;
 wire \thechain[7].chain9.inv_chain[142] ;
 wire \thechain[7].chain9.inv_chain[143] ;
 wire \thechain[7].chain9.inv_chain[144] ;
 wire \thechain[7].chain9.inv_chain[145] ;
 wire \thechain[7].chain9.inv_chain[146] ;
 wire \thechain[7].chain9.inv_chain[147] ;
 wire \thechain[7].chain9.inv_chain[148] ;
 wire \thechain[7].chain9.inv_chain[149] ;
 wire \thechain[7].chain9.inv_chain[14] ;
 wire \thechain[7].chain9.inv_chain[150] ;
 wire \thechain[7].chain9.inv_chain[151] ;
 wire \thechain[7].chain9.inv_chain[152] ;
 wire \thechain[7].chain9.inv_chain[153] ;
 wire \thechain[7].chain9.inv_chain[154] ;
 wire \thechain[7].chain9.inv_chain[155] ;
 wire \thechain[7].chain9.inv_chain[156] ;
 wire \thechain[7].chain9.inv_chain[157] ;
 wire \thechain[7].chain9.inv_chain[158] ;
 wire \thechain[7].chain9.inv_chain[159] ;
 wire \thechain[7].chain9.inv_chain[15] ;
 wire \thechain[7].chain9.inv_chain[160] ;
 wire \thechain[7].chain9.inv_chain[161] ;
 wire \thechain[7].chain9.inv_chain[162] ;
 wire \thechain[7].chain9.inv_chain[163] ;
 wire \thechain[7].chain9.inv_chain[164] ;
 wire \thechain[7].chain9.inv_chain[165] ;
 wire \thechain[7].chain9.inv_chain[166] ;
 wire \thechain[7].chain9.inv_chain[167] ;
 wire \thechain[7].chain9.inv_chain[168] ;
 wire \thechain[7].chain9.inv_chain[169] ;
 wire \thechain[7].chain9.inv_chain[16] ;
 wire \thechain[7].chain9.inv_chain[170] ;
 wire \thechain[7].chain9.inv_chain[171] ;
 wire \thechain[7].chain9.inv_chain[172] ;
 wire \thechain[7].chain9.inv_chain[173] ;
 wire \thechain[7].chain9.inv_chain[174] ;
 wire \thechain[7].chain9.inv_chain[175] ;
 wire \thechain[7].chain9.inv_chain[176] ;
 wire \thechain[7].chain9.inv_chain[177] ;
 wire \thechain[7].chain9.inv_chain[178] ;
 wire \thechain[7].chain9.inv_chain[179] ;
 wire \thechain[7].chain9.inv_chain[17] ;
 wire \thechain[7].chain9.inv_chain[180] ;
 wire \thechain[7].chain9.inv_chain[181] ;
 wire \thechain[7].chain9.inv_chain[182] ;
 wire \thechain[7].chain9.inv_chain[183] ;
 wire \thechain[7].chain9.inv_chain[184] ;
 wire \thechain[7].chain9.inv_chain[185] ;
 wire \thechain[7].chain9.inv_chain[186] ;
 wire \thechain[7].chain9.inv_chain[187] ;
 wire \thechain[7].chain9.inv_chain[188] ;
 wire \thechain[7].chain9.inv_chain[189] ;
 wire \thechain[7].chain9.inv_chain[18] ;
 wire \thechain[7].chain9.inv_chain[190] ;
 wire \thechain[7].chain9.inv_chain[191] ;
 wire \thechain[7].chain9.inv_chain[192] ;
 wire \thechain[7].chain9.inv_chain[193] ;
 wire \thechain[7].chain9.inv_chain[194] ;
 wire \thechain[7].chain9.inv_chain[195] ;
 wire \thechain[7].chain9.inv_chain[196] ;
 wire \thechain[7].chain9.inv_chain[197] ;
 wire \thechain[7].chain9.inv_chain[198] ;
 wire \thechain[7].chain9.inv_chain[199] ;
 wire \thechain[7].chain9.inv_chain[19] ;
 wire \thechain[7].chain9.inv_chain[1] ;
 wire \thechain[7].chain9.inv_chain[200] ;
 wire \thechain[7].chain9.inv_chain[201] ;
 wire \thechain[7].chain9.inv_chain[202] ;
 wire \thechain[7].chain9.inv_chain[203] ;
 wire \thechain[7].chain9.inv_chain[204] ;
 wire \thechain[7].chain9.inv_chain[205] ;
 wire \thechain[7].chain9.inv_chain[206] ;
 wire \thechain[7].chain9.inv_chain[207] ;
 wire \thechain[7].chain9.inv_chain[208] ;
 wire \thechain[7].chain9.inv_chain[209] ;
 wire \thechain[7].chain9.inv_chain[20] ;
 wire \thechain[7].chain9.inv_chain[210] ;
 wire \thechain[7].chain9.inv_chain[211] ;
 wire \thechain[7].chain9.inv_chain[212] ;
 wire \thechain[7].chain9.inv_chain[213] ;
 wire \thechain[7].chain9.inv_chain[214] ;
 wire \thechain[7].chain9.inv_chain[215] ;
 wire \thechain[7].chain9.inv_chain[216] ;
 wire \thechain[7].chain9.inv_chain[217] ;
 wire \thechain[7].chain9.inv_chain[218] ;
 wire \thechain[7].chain9.inv_chain[219] ;
 wire \thechain[7].chain9.inv_chain[21] ;
 wire \thechain[7].chain9.inv_chain[220] ;
 wire \thechain[7].chain9.inv_chain[221] ;
 wire \thechain[7].chain9.inv_chain[222] ;
 wire \thechain[7].chain9.inv_chain[223] ;
 wire \thechain[7].chain9.inv_chain[224] ;
 wire \thechain[7].chain9.inv_chain[225] ;
 wire \thechain[7].chain9.inv_chain[226] ;
 wire \thechain[7].chain9.inv_chain[227] ;
 wire \thechain[7].chain9.inv_chain[228] ;
 wire \thechain[7].chain9.inv_chain[229] ;
 wire \thechain[7].chain9.inv_chain[22] ;
 wire \thechain[7].chain9.inv_chain[230] ;
 wire \thechain[7].chain9.inv_chain[231] ;
 wire \thechain[7].chain9.inv_chain[232] ;
 wire \thechain[7].chain9.inv_chain[233] ;
 wire \thechain[7].chain9.inv_chain[234] ;
 wire \thechain[7].chain9.inv_chain[235] ;
 wire \thechain[7].chain9.inv_chain[236] ;
 wire \thechain[7].chain9.inv_chain[237] ;
 wire \thechain[7].chain9.inv_chain[238] ;
 wire \thechain[7].chain9.inv_chain[239] ;
 wire \thechain[7].chain9.inv_chain[23] ;
 wire \thechain[7].chain9.inv_chain[240] ;
 wire \thechain[7].chain9.inv_chain[241] ;
 wire \thechain[7].chain9.inv_chain[242] ;
 wire \thechain[7].chain9.inv_chain[243] ;
 wire \thechain[7].chain9.inv_chain[244] ;
 wire \thechain[7].chain9.inv_chain[245] ;
 wire \thechain[7].chain9.inv_chain[246] ;
 wire \thechain[7].chain9.inv_chain[247] ;
 wire \thechain[7].chain9.inv_chain[248] ;
 wire \thechain[7].chain9.inv_chain[249] ;
 wire \thechain[7].chain9.inv_chain[24] ;
 wire \thechain[7].chain9.inv_chain[250] ;
 wire \thechain[7].chain9.inv_chain[251] ;
 wire \thechain[7].chain9.inv_chain[252] ;
 wire \thechain[7].chain9.inv_chain[253] ;
 wire \thechain[7].chain9.inv_chain[254] ;
 wire \thechain[7].chain9.inv_chain[255] ;
 wire \thechain[7].chain9.inv_chain[256] ;
 wire \thechain[7].chain9.inv_chain[25] ;
 wire \thechain[7].chain9.inv_chain[26] ;
 wire \thechain[7].chain9.inv_chain[27] ;
 wire \thechain[7].chain9.inv_chain[28] ;
 wire \thechain[7].chain9.inv_chain[29] ;
 wire \thechain[7].chain9.inv_chain[2] ;
 wire \thechain[7].chain9.inv_chain[30] ;
 wire \thechain[7].chain9.inv_chain[31] ;
 wire \thechain[7].chain9.inv_chain[32] ;
 wire \thechain[7].chain9.inv_chain[33] ;
 wire \thechain[7].chain9.inv_chain[34] ;
 wire \thechain[7].chain9.inv_chain[35] ;
 wire \thechain[7].chain9.inv_chain[36] ;
 wire \thechain[7].chain9.inv_chain[37] ;
 wire \thechain[7].chain9.inv_chain[38] ;
 wire \thechain[7].chain9.inv_chain[39] ;
 wire \thechain[7].chain9.inv_chain[3] ;
 wire \thechain[7].chain9.inv_chain[40] ;
 wire \thechain[7].chain9.inv_chain[41] ;
 wire \thechain[7].chain9.inv_chain[42] ;
 wire \thechain[7].chain9.inv_chain[43] ;
 wire \thechain[7].chain9.inv_chain[44] ;
 wire \thechain[7].chain9.inv_chain[45] ;
 wire \thechain[7].chain9.inv_chain[46] ;
 wire \thechain[7].chain9.inv_chain[47] ;
 wire \thechain[7].chain9.inv_chain[48] ;
 wire \thechain[7].chain9.inv_chain[49] ;
 wire \thechain[7].chain9.inv_chain[4] ;
 wire \thechain[7].chain9.inv_chain[50] ;
 wire \thechain[7].chain9.inv_chain[51] ;
 wire \thechain[7].chain9.inv_chain[52] ;
 wire \thechain[7].chain9.inv_chain[53] ;
 wire \thechain[7].chain9.inv_chain[54] ;
 wire \thechain[7].chain9.inv_chain[55] ;
 wire \thechain[7].chain9.inv_chain[56] ;
 wire \thechain[7].chain9.inv_chain[57] ;
 wire \thechain[7].chain9.inv_chain[58] ;
 wire \thechain[7].chain9.inv_chain[59] ;
 wire \thechain[7].chain9.inv_chain[5] ;
 wire \thechain[7].chain9.inv_chain[60] ;
 wire \thechain[7].chain9.inv_chain[61] ;
 wire \thechain[7].chain9.inv_chain[62] ;
 wire \thechain[7].chain9.inv_chain[63] ;
 wire \thechain[7].chain9.inv_chain[64] ;
 wire \thechain[7].chain9.inv_chain[65] ;
 wire \thechain[7].chain9.inv_chain[66] ;
 wire \thechain[7].chain9.inv_chain[67] ;
 wire \thechain[7].chain9.inv_chain[68] ;
 wire \thechain[7].chain9.inv_chain[69] ;
 wire \thechain[7].chain9.inv_chain[6] ;
 wire \thechain[7].chain9.inv_chain[70] ;
 wire \thechain[7].chain9.inv_chain[71] ;
 wire \thechain[7].chain9.inv_chain[72] ;
 wire \thechain[7].chain9.inv_chain[73] ;
 wire \thechain[7].chain9.inv_chain[74] ;
 wire \thechain[7].chain9.inv_chain[75] ;
 wire \thechain[7].chain9.inv_chain[76] ;
 wire \thechain[7].chain9.inv_chain[77] ;
 wire \thechain[7].chain9.inv_chain[78] ;
 wire \thechain[7].chain9.inv_chain[79] ;
 wire \thechain[7].chain9.inv_chain[7] ;
 wire \thechain[7].chain9.inv_chain[80] ;
 wire \thechain[7].chain9.inv_chain[81] ;
 wire \thechain[7].chain9.inv_chain[82] ;
 wire \thechain[7].chain9.inv_chain[83] ;
 wire \thechain[7].chain9.inv_chain[84] ;
 wire \thechain[7].chain9.inv_chain[85] ;
 wire \thechain[7].chain9.inv_chain[86] ;
 wire \thechain[7].chain9.inv_chain[87] ;
 wire \thechain[7].chain9.inv_chain[88] ;
 wire \thechain[7].chain9.inv_chain[89] ;
 wire \thechain[7].chain9.inv_chain[8] ;
 wire \thechain[7].chain9.inv_chain[90] ;
 wire \thechain[7].chain9.inv_chain[91] ;
 wire \thechain[7].chain9.inv_chain[92] ;
 wire \thechain[7].chain9.inv_chain[93] ;
 wire \thechain[7].chain9.inv_chain[94] ;
 wire \thechain[7].chain9.inv_chain[95] ;
 wire \thechain[7].chain9.inv_chain[96] ;
 wire \thechain[7].chain9.inv_chain[97] ;
 wire \thechain[7].chain9.inv_chain[98] ;
 wire \thechain[7].chain9.inv_chain[99] ;
 wire \thechain[7].chain9.inv_chain[9] ;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;

 sky130_fd_sc_hd__mux2_1 _072_ (.A0(net137),
    .A1(\thechain[0].chain1.inv_chain[2] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _073_ (.A0(net146),
    .A1(\thechain[0].chain2.inv_chain[4] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _074_ (.A0(net155),
    .A1(\thechain[0].chain3.inv_chain[8] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _075_ (.A0(net164),
    .A1(\thechain[0].chain4.inv_chain[16] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _076_ (.A0(net162),
    .A1(\thechain[0].chain5.inv_chain[32] ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _077_ (.A0(net135),
    .A1(\thechain[0].chain6.inv_chain[64] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(net124),
    .A1(\thechain[0].chain7.inv_chain[128] ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _079_ (.A0(\thechain[0].chain8.inv_chain[0] ),
    .A1(\thechain[0].chain8.inv_chain[192] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _080_ (.A0(net169),
    .A1(\thechain[0].chain9.inv_chain[256] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _081_ (.A0(net150),
    .A1(\thechain[1].chain1.inv_chain[2] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _082_ (.A0(net153),
    .A1(\thechain[1].chain2.inv_chain[4] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _083_ (.A0(net133),
    .A1(\thechain[1].chain3.inv_chain[8] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _084_ (.A0(net182),
    .A1(\thechain[1].chain4.inv_chain[16] ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _085_ (.A0(net151),
    .A1(\thechain[1].chain5.inv_chain[32] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _086_ (.A0(net156),
    .A1(\thechain[1].chain6.inv_chain[64] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _087_ (.A0(net167),
    .A1(\thechain[1].chain7.inv_chain[128] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _088_ (.A0(net183),
    .A1(\thechain[1].chain8.inv_chain[192] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _089_ (.A0(net154),
    .A1(\thechain[1].chain9.inv_chain[256] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _090_ (.A0(net122),
    .A1(\thechain[2].chain1.inv_chain[2] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _091_ (.A0(net147),
    .A1(\thechain[2].chain2.inv_chain[4] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _092_ (.A0(net163),
    .A1(\thechain[2].chain3.inv_chain[8] ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _093_ (.A0(net142),
    .A1(\thechain[2].chain4.inv_chain[16] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _094_ (.A0(\thechain[2].chain5.inv_chain[0] ),
    .A1(\thechain[2].chain5.inv_chain[32] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _095_ (.A0(net134),
    .A1(\thechain[2].chain6.inv_chain[64] ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _096_ (.A0(net175),
    .A1(\thechain[2].chain7.inv_chain[128] ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _097_ (.A0(\thechain[2].chain8.inv_chain[0] ),
    .A1(\thechain[2].chain8.inv_chain[192] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _098_ (.A0(net139),
    .A1(\thechain[2].chain9.inv_chain[256] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _099_ (.A0(net132),
    .A1(\thechain[3].chain1.inv_chain[2] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _100_ (.A0(net149),
    .A1(\thechain[3].chain2.inv_chain[4] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _101_ (.A0(net173),
    .A1(\thechain[3].chain3.inv_chain[8] ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(net158),
    .A1(\thechain[3].chain4.inv_chain[16] ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _103_ (.A0(net172),
    .A1(\thechain[3].chain5.inv_chain[32] ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _104_ (.A0(net141),
    .A1(\thechain[3].chain6.inv_chain[64] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _105_ (.A0(net145),
    .A1(\thechain[3].chain7.inv_chain[128] ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _106_ (.A0(\thechain[3].chain8.inv_chain[0] ),
    .A1(\thechain[3].chain8.inv_chain[192] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _107_ (.A0(net166),
    .A1(\thechain[3].chain9.inv_chain[256] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _108_ (.A0(net143),
    .A1(\thechain[4].chain1.inv_chain[2] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _109_ (.A0(net125),
    .A1(\thechain[4].chain2.inv_chain[4] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _110_ (.A0(net157),
    .A1(\thechain[4].chain3.inv_chain[8] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _111_ (.A0(net174),
    .A1(\thechain[4].chain4.inv_chain[16] ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _112_ (.A0(net180),
    .A1(\thechain[4].chain5.inv_chain[32] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _113_ (.A0(net152),
    .A1(\thechain[4].chain6.inv_chain[64] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _114_ (.A0(net165),
    .A1(\thechain[4].chain7.inv_chain[128] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _115_ (.A0(\thechain[4].chain8.inv_chain[0] ),
    .A1(\thechain[4].chain8.inv_chain[192] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _116_ (.A0(net123),
    .A1(\thechain[4].chain9.inv_chain[256] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _117_ (.A0(net129),
    .A1(\thechain[5].chain1.inv_chain[2] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _118_ (.A0(net138),
    .A1(\thechain[5].chain2.inv_chain[4] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _119_ (.A0(net168),
    .A1(\thechain[5].chain3.inv_chain[8] ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _120_ (.A0(net120),
    .A1(\thechain[5].chain4.inv_chain[16] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _121_ (.A0(net176),
    .A1(\thechain[5].chain5.inv_chain[32] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _122_ (.A0(net130),
    .A1(\thechain[5].chain6.inv_chain[64] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _123_ (.A0(net177),
    .A1(\thechain[5].chain7.inv_chain[128] ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _124_ (.A0(\thechain[5].chain8.inv_chain[0] ),
    .A1(\thechain[5].chain8.inv_chain[192] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _125_ (.A0(net126),
    .A1(\thechain[5].chain9.inv_chain[256] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _126_ (.A0(net121),
    .A1(\thechain[6].chain1.inv_chain[2] ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _127_ (.A0(net128),
    .A1(\thechain[6].chain2.inv_chain[4] ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _128_ (.A0(net160),
    .A1(\thechain[6].chain3.inv_chain[8] ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _129_ (.A0(\thechain[6].chain4.inv_chain[0] ),
    .A1(\thechain[6].chain4.inv_chain[16] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _130_ (.A0(net148),
    .A1(\thechain[6].chain5.inv_chain[32] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _131_ (.A0(net136),
    .A1(\thechain[6].chain6.inv_chain[64] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _132_ (.A0(net161),
    .A1(\thechain[6].chain7.inv_chain[128] ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _133_ (.A0(\thechain[6].chain8.inv_chain[0] ),
    .A1(\thechain[6].chain8.inv_chain[192] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _134_ (.A0(net181),
    .A1(\thechain[6].chain9.inv_chain[256] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _135_ (.A0(net131),
    .A1(\thechain[7].chain1.inv_chain[2] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _136_ (.A0(net144),
    .A1(\thechain[7].chain2.inv_chain[4] ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _137_ (.A0(net140),
    .A1(\thechain[7].chain3.inv_chain[8] ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _138_ (.A0(net170),
    .A1(\thechain[7].chain4.inv_chain[16] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _139_ (.A0(net159),
    .A1(\thechain[7].chain5.inv_chain[32] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _140_ (.A0(net171),
    .A1(\thechain[7].chain6.inv_chain[64] ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _141_ (.A0(net127),
    .A1(\thechain[7].chain7.inv_chain[128] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _142_ (.A0(net179),
    .A1(\thechain[7].chain8.inv_chain[192] ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _143_ (.A0(net178),
    .A1(\thechain[7].chain9.inv_chain[256] ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_071_));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(clknet_4_2_0_clk),
    .D(net76),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _145_ (.CLK(clknet_4_10_0_clk),
    .D(_071_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _146_ (.CLK(clknet_4_15_0_clk),
    .D(_000_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _147_ (.CLK(clknet_4_15_0_clk),
    .D(net2),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _148_ (.CLK(clknet_4_15_0_clk),
    .D(_001_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _149_ (.CLK(clknet_4_15_0_clk),
    .D(net102),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _150_ (.CLK(clknet_4_15_0_clk),
    .D(_002_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _151_ (.CLK(clknet_4_15_0_clk),
    .D(net88),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _152_ (.CLK(clknet_4_13_0_clk),
    .D(_003_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _153_ (.CLK(clknet_4_15_0_clk),
    .D(net84),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _154_ (.CLK(clknet_4_13_0_clk),
    .D(_004_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _155_ (.CLK(clknet_4_13_0_clk),
    .D(net92),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _156_ (.CLK(clknet_4_7_0_clk),
    .D(_005_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _157_ (.CLK(clknet_4_7_0_clk),
    .D(net116),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _158_ (.CLK(clknet_4_13_0_clk),
    .D(_006_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _159_ (.CLK(clknet_4_7_0_clk),
    .D(net69),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _160_ (.CLK(clknet_4_8_0_clk),
    .D(_007_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_1 _161_ (.CLK(clknet_4_13_0_clk),
    .D(net86),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _162_ (.CLK(clknet_4_11_0_clk),
    .D(_008_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _163_ (.CLK(clknet_4_9_0_clk),
    .D(net103),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[0].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _164_ (.CLK(clknet_4_15_0_clk),
    .D(_009_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _165_ (.CLK(clknet_4_15_0_clk),
    .D(net3),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _166_ (.CLK(clknet_4_15_0_clk),
    .D(_010_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _167_ (.CLK(clknet_4_15_0_clk),
    .D(net105),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _168_ (.CLK(clknet_4_13_0_clk),
    .D(_011_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _169_ (.CLK(clknet_4_13_0_clk),
    .D(net112),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _170_ (.CLK(clknet_4_6_0_clk),
    .D(_012_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _171_ (.CLK(clknet_4_13_0_clk),
    .D(net109),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _172_ (.CLK(clknet_4_7_0_clk),
    .D(_013_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _173_ (.CLK(clknet_4_7_0_clk),
    .D(net70),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _174_ (.CLK(clknet_4_5_0_clk),
    .D(_014_),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _175_ (.CLK(clknet_4_7_0_clk),
    .D(net94),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _176_ (.CLK(clknet_4_5_0_clk),
    .D(_015_),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _177_ (.CLK(clknet_4_5_0_clk),
    .D(net64),
    .RESET_B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _178_ (.CLK(clknet_4_3_0_clk),
    .D(_016_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_1 _179_ (.CLK(clknet_4_5_0_clk),
    .D(net60),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _180_ (.CLK(clknet_4_6_0_clk),
    .D(_017_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _181_ (.CLK(clknet_4_3_0_clk),
    .D(net68),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[1].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _182_ (.CLK(clknet_4_14_0_clk),
    .D(_018_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _183_ (.CLK(clknet_4_14_0_clk),
    .D(net4),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _184_ (.CLK(clknet_4_14_0_clk),
    .D(_019_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _185_ (.CLK(clknet_4_15_0_clk),
    .D(net80),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _186_ (.CLK(clknet_4_15_0_clk),
    .D(_020_),
    .RESET_B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _187_ (.CLK(clknet_4_15_0_clk),
    .D(net56),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _188_ (.CLK(clknet_4_12_0_clk),
    .D(_021_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _189_ (.CLK(clknet_4_12_0_clk),
    .D(net115),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _190_ (.CLK(clknet_4_4_0_clk),
    .D(_022_),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _191_ (.CLK(clknet_4_13_0_clk),
    .D(net114),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _192_ (.CLK(clknet_4_5_0_clk),
    .D(_023_),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _193_ (.CLK(clknet_4_4_0_clk),
    .D(net77),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _194_ (.CLK(clknet_4_4_0_clk),
    .D(_024_),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _195_ (.CLK(clknet_4_5_0_clk),
    .D(net93),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _196_ (.CLK(clknet_4_8_0_clk),
    .D(_025_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_2 _197_ (.CLK(clknet_4_5_0_clk),
    .D(net95),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _198_ (.CLK(clknet_4_8_0_clk),
    .D(_026_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _199_ (.CLK(clknet_4_8_0_clk),
    .D(net62),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[2].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _200_ (.CLK(clknet_4_14_0_clk),
    .D(_027_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _201_ (.CLK(clknet_4_14_0_clk),
    .D(net5),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _202_ (.CLK(clknet_4_14_0_clk),
    .D(_028_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _203_ (.CLK(clknet_4_14_0_clk),
    .D(net61),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _204_ (.CLK(clknet_4_12_0_clk),
    .D(_029_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _205_ (.CLK(clknet_4_15_0_clk),
    .D(net58),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _206_ (.CLK(clknet_4_12_0_clk),
    .D(_030_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _207_ (.CLK(clknet_4_13_0_clk),
    .D(net57),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _208_ (.CLK(clknet_4_1_0_clk),
    .D(_031_),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _209_ (.CLK(clknet_4_7_0_clk),
    .D(net119),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _210_ (.CLK(clknet_4_1_0_clk),
    .D(_032_),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _211_ (.CLK(clknet_4_1_0_clk),
    .D(net113),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _212_ (.CLK(clknet_4_4_0_clk),
    .D(_033_),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _213_ (.CLK(clknet_4_4_0_clk),
    .D(net59),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _214_ (.CLK(clknet_4_8_0_clk),
    .D(_034_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_2 _215_ (.CLK(clknet_4_4_0_clk),
    .D(net65),
    .RESET_B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _216_ (.CLK(clknet_4_8_0_clk),
    .D(_035_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _217_ (.CLK(clknet_4_8_0_clk),
    .D(net63),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[3].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _218_ (.CLK(clknet_4_11_0_clk),
    .D(_036_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _219_ (.CLK(clknet_4_11_0_clk),
    .D(net6),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _220_ (.CLK(clknet_4_14_0_clk),
    .D(_037_),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _221_ (.CLK(clknet_4_14_0_clk),
    .D(net87),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _222_ (.CLK(clknet_4_12_0_clk),
    .D(_038_),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _223_ (.CLK(clknet_4_14_0_clk),
    .D(net83),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _224_ (.CLK(clknet_4_6_0_clk),
    .D(_039_),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _225_ (.CLK(clknet_4_12_0_clk),
    .D(net97),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _226_ (.CLK(clknet_4_1_0_clk),
    .D(_040_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _227_ (.CLK(clknet_4_3_0_clk),
    .D(net117),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _228_ (.CLK(clknet_4_0_0_clk),
    .D(_041_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _229_ (.CLK(clknet_4_0_0_clk),
    .D(net104),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _230_ (.CLK(clknet_4_0_0_clk),
    .D(_042_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _231_ (.CLK(clknet_4_1_0_clk),
    .D(net100),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _232_ (.CLK(clknet_4_10_0_clk),
    .D(_043_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_2 _233_ (.CLK(clknet_4_0_0_clk),
    .D(net99),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _234_ (.CLK(clknet_4_10_0_clk),
    .D(_044_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _235_ (.CLK(clknet_4_10_0_clk),
    .D(net73),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[4].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _236_ (.CLK(clknet_4_11_0_clk),
    .D(_045_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _237_ (.CLK(clknet_4_11_0_clk),
    .D(net7),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _238_ (.CLK(clknet_4_11_0_clk),
    .D(_046_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _239_ (.CLK(clknet_4_11_0_clk),
    .D(net81),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _240_ (.CLK(clknet_4_9_0_clk),
    .D(_047_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _241_ (.CLK(clknet_4_11_0_clk),
    .D(net108),
    .RESET_B(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _242_ (.CLK(clknet_4_9_0_clk),
    .D(_048_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _243_ (.CLK(clknet_4_9_0_clk),
    .D(net72),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _244_ (.CLK(clknet_4_3_0_clk),
    .D(_049_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _245_ (.CLK(clknet_4_12_0_clk),
    .D(net91),
    .RESET_B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _246_ (.CLK(clknet_4_6_0_clk),
    .D(_050_),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _247_ (.CLK(clknet_4_3_0_clk),
    .D(net98),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _248_ (.CLK(clknet_4_2_0_clk),
    .D(_051_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _249_ (.CLK(clknet_4_6_0_clk),
    .D(net96),
    .RESET_B(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _250_ (.CLK(clknet_4_10_0_clk),
    .D(_052_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_1 _251_ (.CLK(clknet_4_2_0_clk),
    .D(net85),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _252_ (.CLK(clknet_4_10_0_clk),
    .D(_053_),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _253_ (.CLK(clknet_4_10_0_clk),
    .D(net74),
    .RESET_B(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[5].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _254_ (.CLK(clknet_4_10_0_clk),
    .D(_054_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _255_ (.CLK(clknet_4_11_0_clk),
    .D(net8),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _256_ (.CLK(clknet_4_11_0_clk),
    .D(_055_),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _257_ (.CLK(clknet_4_11_0_clk),
    .D(net110),
    .RESET_B(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _258_ (.CLK(clknet_4_9_0_clk),
    .D(_056_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _259_ (.CLK(clknet_4_11_0_clk),
    .D(net66),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _260_ (.CLK(clknet_4_3_0_clk),
    .D(_057_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _261_ (.CLK(clknet_4_12_0_clk),
    .D(net71),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _262_ (.CLK(clknet_4_0_0_clk),
    .D(_058_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _263_ (.CLK(clknet_4_0_0_clk),
    .D(net118),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _264_ (.CLK(clknet_4_0_0_clk),
    .D(_059_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _265_ (.CLK(clknet_4_0_0_clk),
    .D(net90),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _266_ (.CLK(clknet_4_1_0_clk),
    .D(_060_),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _267_ (.CLK(clknet_4_0_0_clk),
    .D(net78),
    .RESET_B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _268_ (.CLK(clknet_4_2_0_clk),
    .D(_061_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_1 _269_ (.CLK(clknet_4_1_0_clk),
    .D(net67),
    .RESET_B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _270_ (.CLK(clknet_4_10_0_clk),
    .D(_062_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain9.dout ));
 sky130_fd_sc_hd__dfrtp_1 _271_ (.CLK(clknet_4_2_0_clk),
    .D(net79),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[6].chain9.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _272_ (.CLK(clknet_4_10_0_clk),
    .D(_063_),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.dout ));
 sky130_fd_sc_hd__dfrtp_1 _273_ (.CLK(clknet_4_10_0_clk),
    .D(net9),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain1.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _274_ (.CLK(clknet_4_8_0_clk),
    .D(_064_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain2.dout ));
 sky130_fd_sc_hd__dfrtp_1 _275_ (.CLK(clknet_4_10_0_clk),
    .D(net101),
    .RESET_B(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain2.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _276_ (.CLK(clknet_4_9_0_clk),
    .D(_065_),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain3.dout ));
 sky130_fd_sc_hd__dfrtp_1 _277_ (.CLK(clknet_4_9_0_clk),
    .D(net107),
    .RESET_B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain3.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _278_ (.CLK(clknet_4_2_0_clk),
    .D(_066_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain4.dout ));
 sky130_fd_sc_hd__dfrtp_1 _279_ (.CLK(clknet_4_8_0_clk),
    .D(net111),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain4.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _280_ (.CLK(clknet_4_2_0_clk),
    .D(_067_),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain5.dout ));
 sky130_fd_sc_hd__dfrtp_1 _281_ (.CLK(clknet_4_2_0_clk),
    .D(net106),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain5.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _282_ (.CLK(clknet_4_3_0_clk),
    .D(_068_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain6.dout ));
 sky130_fd_sc_hd__dfrtp_1 _283_ (.CLK(clknet_4_2_0_clk),
    .D(net89),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain6.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _284_ (.CLK(clknet_4_3_0_clk),
    .D(_069_),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain7.dout ));
 sky130_fd_sc_hd__dfrtp_1 _285_ (.CLK(clknet_4_3_0_clk),
    .D(net82),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain7.inv_chain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _286_ (.CLK(clknet_4_2_0_clk),
    .D(_070_),
    .RESET_B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain8.dout ));
 sky130_fd_sc_hd__dfrtp_1 _287_ (.CLK(clknet_4_3_0_clk),
    .D(net75),
    .RESET_B(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\thechain[7].chain8.inv_chain[0] ));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net41));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net42));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net43));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net44));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net45));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net46));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net47));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net48));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net49));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net50));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net51));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net52));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net53));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net54));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net55));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_2 _304_ (.A(\thechain[0].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _305_ (.A(\thechain[1].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__clkbuf_4 _306_ (.A(\thechain[2].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__clkbuf_4 _307_ (.A(\thechain[3].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _308_ (.A(\thechain[4].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _309_ (.A(\thechain[5].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _310_ (.A(\thechain[6].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _311_ (.A(\thechain[7].chain9.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[0].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[0].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[0].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[0].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[0].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[0].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[0].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[0].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[1].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[1].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[1].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[1].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[1].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[1].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[1].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[1].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[2].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[2].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[2].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[2].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[2].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[2].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[2].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[2].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[3].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[3].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[3].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[3].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[3].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[3].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[3].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[3].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[4].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[4].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[4].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[4].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[4].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[4].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[4].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[4].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[5].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[5].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[5].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[5].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[5].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[5].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[5].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[5].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[6].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[6].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[6].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[6].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[6].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[6].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[6].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[6].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain1.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain1.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain1.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain2.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain2.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain2.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain2.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain2.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain2.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain2.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain2.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain2.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain2.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain2.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain3.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain3.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain3.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[10].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[11].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[12].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[13].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[14].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[15].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[8].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain4.inv_pair[9].inv_gate/_0_  (.A(\thechain[7].chain4.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain4.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[10].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[11].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[12].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[13].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[14].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[15].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[16].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[17].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[18].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[19].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[20].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[21].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[22].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[23].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[24].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[25].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[26].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[27].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[28].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[29].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[30].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[31].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[8].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain5.inv_pair[9].inv_gate/_0_  (.A(\thechain[7].chain5.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain5.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[10].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[11].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[12].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[13].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[14].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[15].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[16].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[17].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[18].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[19].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[20].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[21].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[22].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[23].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[24].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[25].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[26].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[27].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[28].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[29].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[30].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[31].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[32].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[33].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[34].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[35].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[36].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[37].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[38].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[39].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[40].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[41].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[42].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[43].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[44].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[45].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[46].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[47].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[48].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[49].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[50].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[51].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[52].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[53].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[54].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[55].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[56].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[57].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[58].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[59].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[60].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[61].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[62].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[63].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[8].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain6.inv_pair[9].inv_gate/_0_  (.A(\thechain[7].chain6.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain6.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[100].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[101].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[102].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[103].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[104].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[105].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[106].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[107].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[108].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[109].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[10].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[110].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[111].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[112].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[113].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[114].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[115].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[116].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[117].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[118].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[119].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[11].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[120].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[121].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[122].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[123].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[124].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[125].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[126].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[127].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[12].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[13].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[14].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[15].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[16].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[17].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[18].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[19].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[20].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[21].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[22].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[23].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[24].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[25].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[26].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[27].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[28].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[29].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[30].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[31].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[32].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[33].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[34].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[35].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[36].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[37].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[38].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[39].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[40].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[41].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[42].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[43].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[44].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[45].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[46].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[47].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[48].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[49].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[50].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[51].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[52].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[53].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[54].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[55].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[56].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[57].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[58].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[59].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[60].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[61].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[62].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[63].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[64].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[65].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[66].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[67].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[68].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[69].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[70].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[71].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[72].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[73].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[74].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[75].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[76].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[77].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[78].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[79].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[80].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[81].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[82].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[83].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[84].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[85].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[86].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[87].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[88].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[89].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[8].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[90].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[91].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[92].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[93].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[94].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[95].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[96].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[97].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[98].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[99].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain7.inv_pair[9].inv_gate/_0_  (.A(\thechain[7].chain7.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain7.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[100].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[101].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[102].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[103].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[104].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[105].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[106].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[107].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[108].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[109].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[10].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[110].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[111].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[112].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[113].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[114].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[115].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[116].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[117].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[118].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[119].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[11].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[120].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[121].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[122].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[123].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[124].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[125].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[126].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[127].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[128].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[129].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[12].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[130].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[131].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[132].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[133].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[134].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[135].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[136].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[137].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[138].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[139].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[13].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[140].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[141].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[142].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[143].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[144].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[145].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[146].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[147].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[148].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[149].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[14].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[150].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[151].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[152].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[153].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[154].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[155].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[156].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[157].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[158].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[159].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[15].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[160].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[161].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[162].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[163].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[164].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[165].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[166].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[167].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[168].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[169].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[16].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[170].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[171].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[172].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[173].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[174].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[175].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[176].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[177].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[178].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[179].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[17].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[180].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[181].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[182].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[183].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[184].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[185].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[186].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[187].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[188].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[189].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[18].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[190].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[191].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[19].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[20].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[21].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[22].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[23].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[24].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[25].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[26].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[27].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[28].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[29].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[30].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[31].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[32].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[33].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[34].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[35].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[36].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[37].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[38].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[39].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[40].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[41].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[42].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[43].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[44].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[45].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[46].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[47].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[48].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[49].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[50].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[51].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[52].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[53].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[54].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[55].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[56].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[57].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[58].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[59].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[60].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[61].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[62].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[63].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[64].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[65].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[66].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[67].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[68].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[69].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[70].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[71].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[72].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[73].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[74].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[75].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[76].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[77].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[78].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[79].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[80].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[81].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[82].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[83].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[84].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[85].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[86].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[87].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[88].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[89].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[8].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[90].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[91].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[92].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[93].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[94].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[95].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[96].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[97].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[98].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[99].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain8.inv_pair[9].inv_gate/_0_  (.A(\thechain[7].chain8.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain8.inv_chain[10] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[0].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[1] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[100].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[101] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[101].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[102] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[102].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[103] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[103].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[104] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[104].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[105] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[105].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[106] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[106].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[107] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[107].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[108] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[108].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[109] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[109].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[110] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[10].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[11] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[110].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[111] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[111].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[112] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[112].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[113] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[113].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[114] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[114].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[115] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[115].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[116] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[116].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[117] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[117].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[118] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[118].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[119] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[119].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[120] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[11].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[12] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[120].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[121] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[121].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[122] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[122].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[123] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[123].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[124] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[124].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[125] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[125].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[126] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[126].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[127] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[127].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[128] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[128].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[129] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[129].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[130] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[12].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[13] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[130].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[131] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[131].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[132] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[132].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[133] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[133].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[134] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[134].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[135] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[135].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[136] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[136].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[137] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[137].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[138] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[138].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[139] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[139].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[140] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[13].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[14] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[140].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[141] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[141].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[142] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[142].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[143] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[143].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[144] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[144].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[145] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[145].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[146] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[146].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[147] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[147].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[148] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[148].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[149] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[149].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[150] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[14].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[15] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[150].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[151] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[151].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[152] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[152].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[153] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[153].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[154] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[154].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[155] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[155].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[156] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[156].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[157] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[157].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[158] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[158].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[159] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[159].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[160] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[15].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[16] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[160].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[161] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[161].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[162] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[162].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[163] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[163].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[164] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[164].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[165] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[165].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[166] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[166].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[167] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[167].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[168] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[168].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[169] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[169].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[170] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[16].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[17] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[170].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[171] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[171].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[172] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[172].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[173] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[173].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[174] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[174].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[175] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[175].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[176] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[176].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[177] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[177].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[178] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[178].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[179] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[179].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[180] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[17].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[18] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[180].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[181] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[181].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[182] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[182].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[183] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[183].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[184] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[184].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[185] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[185].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[186] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[186].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[187] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[187].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[188] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[188].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[189] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[189].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[190] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[18].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[19] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[190].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[191] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[191].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[192] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[192].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[193] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[193].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[193] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[194] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[194].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[195] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[195].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[196] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[196].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[196] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[197] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[197].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[198] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[198].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[199] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[199].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[199] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[200] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[19].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[20] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[1].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[2] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[200].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[201] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[201].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[202] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[202].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[202] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[203] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[203].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[204] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[204].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[204] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[205] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[205].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[206] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[206].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[206] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[207] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[207].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[208] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[208].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[208] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[209] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[209].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[210] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[20].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[21] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[210].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[210] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[211] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[211].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[212] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[212].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[212] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[213] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[213].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[214] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[214].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[214] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[215] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[215].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[216] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[216].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[216] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[217] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[217].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[218] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[218].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[218] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[219] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[219].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[220] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[21].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[22] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[220].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[220] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[221] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[221].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[222] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[222].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[222] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[223] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[223].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[224] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[224].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[224] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[225] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[225].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[226] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[226].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[226] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[227] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[227].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[228] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[228].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[229] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[229].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[229] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[230] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[22].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[23] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[230].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[231] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[231].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[232] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[232].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[232] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[233] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[233].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[234] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[234].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[235] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[235].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[235] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[236] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[236].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[237] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[237].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[238] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[238].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[238] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[239] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[239].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[240] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[23].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[24] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[240].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[240] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[241] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[241].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[242] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[242].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[242] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[243] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[243].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[244] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[244].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[244] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[245] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[245].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[246] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[246].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[246] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[247] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[247].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[248] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[248].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[249] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[249].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[249] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[250] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[24].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[25] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[250].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[251] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[251].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[252] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[252].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[252] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[253] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[253].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[254] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[254].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[255] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[255].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[255] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[256] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[25].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[26] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[26].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[27] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[27].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[28] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[28].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[29] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[29].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[30] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[2].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[3] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[30].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[31] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[31].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[32] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[32].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[33] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[33].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[34] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[34].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[35] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[35].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[36] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[36].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[37] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[37].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[38] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[38].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[39] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[39].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[40] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[3].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[4] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[40].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[41] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[41].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[42] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[42].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[43] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[43].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[44] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[44].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[45] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[45].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[46] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[46].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[47] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[47].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[48] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[48].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[49] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[49].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[50] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[4].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[5] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[50].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[51] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[51].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[52] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[52].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[53] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[53].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[54] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[54].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[55] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[55].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[56] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[56].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[57] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[57].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[58] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[58].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[59] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[59].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[60] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[5].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[6] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[60].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[61] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[61].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[62] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[62].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[63] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[63].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[64] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[64].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[65] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[65].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[66] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[66].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[67] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[67].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[68] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[68].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[69] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[69].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[70] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[6].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[7] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[70].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[71] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[71].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[72] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[72].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[73] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[73].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[74] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[74].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[75] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[75].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[76] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[76].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[77] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[77].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[78] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[78].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[79] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[79].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[80] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[7].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[8] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[80].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[81] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[81].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[82] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[82].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[83] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[83].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[84] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[84].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[85] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[85].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[86] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[86].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[87] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[87].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[88] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[88].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[89] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[89].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[90] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[8].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[9] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[90].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[91] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[91].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[92] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[92].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[93] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[93].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[94] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[94].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[95] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[95].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[96] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[96].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[97] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[97].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[98] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[98].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[99] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[99].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[100] ));
 sky130_fd_sc_hd__inv_2 \thechain[7].chain9.inv_pair[9].inv_gate/_0_  (.A(\thechain[7].chain9.inv_chain[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\thechain[7].chain9.inv_chain[10] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__buf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_4 fanout12 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 fanout33 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__conb_1 tt_um_delaychain_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net40));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload6 (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload8 (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload11 (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload13 (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload14 (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\thechain[2].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\thechain[3].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\thechain[3].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\thechain[3].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\thechain[1].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\thechain[3].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\thechain[2].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\thechain[3].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\thechain[1].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\thechain[3].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\thechain[6].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\thechain[6].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\thechain[1].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\thechain[0].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\thechain[1].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\thechain[6].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\thechain[5].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\thechain[4].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\thechain[5].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\thechain[7].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\thechain[7].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\thechain[2].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\thechain[6].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\thechain[6].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\thechain[2].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\thechain[5].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\thechain[7].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\thechain[4].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\thechain[0].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\thechain[5].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\thechain[0].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\thechain[4].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\thechain[0].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\thechain[7].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\thechain[6].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\thechain[5].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\thechain[0].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\thechain[2].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\thechain[1].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\thechain[2].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\thechain[5].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\thechain[4].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\thechain[5].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\thechain[4].chain7.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\thechain[4].chain6.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\thechain[7].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\thechain[0].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\thechain[0].chain8.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\thechain[4].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\thechain[1].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\thechain[7].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\thechain[7].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\thechain[5].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\thechain[1].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\thechain[6].chain1.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\thechain[7].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\thechain[1].chain2.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\thechain[3].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\thechain[2].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\thechain[2].chain3.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\thechain[0].chain5.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\thechain[4].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\thechain[6].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\thechain[3].chain4.dout ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\thechain[5].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\thechain[6].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\thechain[2].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\thechain[4].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\thechain[0].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\thechain[4].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\thechain[5].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\thechain[7].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\thechain[6].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\thechain[5].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\thechain[5].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\thechain[7].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\thechain[3].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\thechain[1].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\thechain[2].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\thechain[0].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\thechain[6].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\thechain[0].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\thechain[5].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\thechain[2].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\thechain[7].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\thechain[3].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\thechain[2].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\thechain[4].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\thechain[7].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\thechain[3].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\thechain[0].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\thechain[2].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\thechain[6].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\thechain[3].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\thechain[1].chain1.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\thechain[1].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\thechain[4].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\thechain[1].chain2.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\thechain[1].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\thechain[0].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\thechain[1].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\thechain[4].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\thechain[3].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\thechain[7].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\thechain[6].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\thechain[6].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\thechain[0].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\thechain[2].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\thechain[0].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\thechain[4].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\thechain[3].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\thechain[1].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\thechain[5].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\thechain[0].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\thechain[7].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\thechain[7].chain6.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\thechain[3].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\thechain[3].chain3.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\thechain[4].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\thechain[2].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\thechain[5].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\thechain[5].chain7.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\thechain[7].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\thechain[7].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\thechain[4].chain5.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\thechain[6].chain9.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\thechain[1].chain4.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\thechain[1].chain8.inv_chain[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_226 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_4_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_190 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_7_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_11_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_202 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_41_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_259 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_43_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_44_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_45_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_162 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_46_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_47_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_47_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_48_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_180 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_50_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_51_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_55_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_57_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_246 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_57_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_59_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_62_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_63_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_65_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_66_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_69_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_70_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_71_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_71_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_72_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_72_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_73_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_74_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_75_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_75_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_75_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_75_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_75_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_76_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_76_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_76_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_76_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_77_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_77_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_77_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_77_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_78_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_78_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_78_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_78_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_78_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_79_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_79_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_79_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_80_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_80_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_80_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_80_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_80_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_80_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net40;
 assign uio_oe[1] = net41;
 assign uio_oe[2] = net42;
 assign uio_oe[3] = net43;
 assign uio_oe[4] = net44;
 assign uio_oe[5] = net45;
 assign uio_oe[6] = net46;
 assign uio_oe[7] = net47;
 assign uio_out[0] = net48;
 assign uio_out[1] = net49;
 assign uio_out[2] = net50;
 assign uio_out[3] = net51;
 assign uio_out[4] = net52;
 assign uio_out[5] = net53;
 assign uio_out[6] = net54;
 assign uio_out[7] = net55;
endmodule
