module tt_um_FFT_engine (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire net31;
 wire net32;
 wire clknet_0_clk;
 wire \addr[0] ;
 wire \addr[1] ;
 wire \disp_inst.done ;
 wire \disp_inst.output_counter[0] ;
 wire \disp_inst.output_counter[1] ;
 wire \disp_inst.processing ;
 wire \fft0_imag[4] ;
 wire \fft0_imag[5] ;
 wire \fft0_imag[6] ;
 wire \fft0_imag[7] ;
 wire \fft0_real[4] ;
 wire \fft0_real[5] ;
 wire \fft0_real[6] ;
 wire \fft0_real[7] ;
 wire \fft1_imag[4] ;
 wire \fft1_imag[5] ;
 wire \fft1_imag[6] ;
 wire \fft1_imag[7] ;
 wire \fft1_real[4] ;
 wire \fft1_real[5] ;
 wire \fft1_real[6] ;
 wire \fft1_real[7] ;
 wire \fft2_imag[4] ;
 wire \fft2_imag[5] ;
 wire \fft2_imag[6] ;
 wire \fft2_imag[7] ;
 wire \fft2_real[4] ;
 wire \fft2_real[5] ;
 wire \fft2_real[6] ;
 wire \fft2_real[7] ;
 wire \fft3_imag[4] ;
 wire \fft3_imag[5] ;
 wire \fft3_imag[6] ;
 wire \fft3_imag[7] ;
 wire \fft3_real[4] ;
 wire \fft3_real[5] ;
 wire \fft3_real[6] ;
 wire \fft3_real[7] ;
 wire \fft_inst.bfly_neg_imag[4] ;
 wire \fft_inst.bfly_neg_imag[5] ;
 wire \fft_inst.bfly_neg_imag[6] ;
 wire \fft_inst.bfly_neg_imag[7] ;
 wire \fft_inst.bfly_neg_real[4] ;
 wire \fft_inst.bfly_neg_real[5] ;
 wire \fft_inst.bfly_neg_real[6] ;
 wire \fft_inst.bfly_neg_real[7] ;
 wire \fft_inst.bfly_pos_imag[4] ;
 wire \fft_inst.bfly_pos_imag[5] ;
 wire \fft_inst.bfly_pos_imag[6] ;
 wire \fft_inst.bfly_pos_imag[7] ;
 wire \fft_inst.bfly_pos_real[4] ;
 wire \fft_inst.bfly_pos_real[5] ;
 wire \fft_inst.bfly_pos_real[6] ;
 wire \fft_inst.bfly_pos_real[7] ;
 wire \fft_inst.bfly_stage1_0.A_imag[4] ;
 wire \fft_inst.bfly_stage1_0.A_imag[5] ;
 wire \fft_inst.bfly_stage1_0.A_imag[6] ;
 wire \fft_inst.bfly_stage1_0.A_imag[7] ;
 wire \fft_inst.bfly_stage1_0.A_real[4] ;
 wire \fft_inst.bfly_stage1_0.A_real[5] ;
 wire \fft_inst.bfly_stage1_0.A_real[6] ;
 wire \fft_inst.bfly_stage1_0.A_real[7] ;
 wire \fft_inst.bfly_stage1_0.B_imag[4] ;
 wire \fft_inst.bfly_stage1_0.B_imag[5] ;
 wire \fft_inst.bfly_stage1_0.B_imag[6] ;
 wire \fft_inst.bfly_stage1_0.B_imag[7] ;
 wire \fft_inst.bfly_stage1_0.B_real[4] ;
 wire \fft_inst.bfly_stage1_0.B_real[5] ;
 wire \fft_inst.bfly_stage1_0.B_real[6] ;
 wire \fft_inst.bfly_stage1_0.B_real[7] ;
 wire \fft_inst.bfly_stage1_1.A_imag[4] ;
 wire \fft_inst.bfly_stage1_1.A_imag[5] ;
 wire \fft_inst.bfly_stage1_1.A_imag[6] ;
 wire \fft_inst.bfly_stage1_1.A_imag[7] ;
 wire \fft_inst.bfly_stage1_1.A_real[4] ;
 wire \fft_inst.bfly_stage1_1.A_real[5] ;
 wire \fft_inst.bfly_stage1_1.A_real[6] ;
 wire \fft_inst.bfly_stage1_1.A_real[7] ;
 wire \fft_inst.bfly_stage1_1.B_imag[4] ;
 wire \fft_inst.bfly_stage1_1.B_imag[5] ;
 wire \fft_inst.bfly_stage1_1.B_imag[6] ;
 wire \fft_inst.bfly_stage1_1.B_imag[7] ;
 wire \fft_inst.bfly_stage1_1.B_real[4] ;
 wire \fft_inst.bfly_stage1_1.B_real[5] ;
 wire \fft_inst.bfly_stage1_1.B_real[6] ;
 wire \fft_inst.bfly_stage1_1.B_real[7] ;
 wire \fft_inst.rst ;
 wire \io_inst.prev_in0 ;
 wire \io_inst.prev_in1 ;
 wire \out_delay_gen[0].out_delay_inst.A ;
 wire \out_delay_gen[0].out_delay_inst.X ;
 wire \out_delay_gen[0].out_delay_inst.w1 ;
 wire \out_delay_gen[0].out_delay_inst.w10 ;
 wire \out_delay_gen[0].out_delay_inst.w11 ;
 wire \out_delay_gen[0].out_delay_inst.w12 ;
 wire \out_delay_gen[0].out_delay_inst.w13 ;
 wire \out_delay_gen[0].out_delay_inst.w14 ;
 wire \out_delay_gen[0].out_delay_inst.w15 ;
 wire \out_delay_gen[0].out_delay_inst.w16 ;
 wire \out_delay_gen[0].out_delay_inst.w17 ;
 wire \out_delay_gen[0].out_delay_inst.w18 ;
 wire \out_delay_gen[0].out_delay_inst.w19 ;
 wire \out_delay_gen[0].out_delay_inst.w2 ;
 wire \out_delay_gen[0].out_delay_inst.w20 ;
 wire \out_delay_gen[0].out_delay_inst.w21 ;
 wire \out_delay_gen[0].out_delay_inst.w22 ;
 wire \out_delay_gen[0].out_delay_inst.w23 ;
 wire \out_delay_gen[0].out_delay_inst.w24 ;
 wire \out_delay_gen[0].out_delay_inst.w25 ;
 wire \out_delay_gen[0].out_delay_inst.w26 ;
 wire \out_delay_gen[0].out_delay_inst.w27 ;
 wire \out_delay_gen[0].out_delay_inst.w28 ;
 wire \out_delay_gen[0].out_delay_inst.w29 ;
 wire \out_delay_gen[0].out_delay_inst.w3 ;
 wire \out_delay_gen[0].out_delay_inst.w30 ;
 wire \out_delay_gen[0].out_delay_inst.w31 ;
 wire \out_delay_gen[0].out_delay_inst.w32 ;
 wire \out_delay_gen[0].out_delay_inst.w33 ;
 wire \out_delay_gen[0].out_delay_inst.w34 ;
 wire \out_delay_gen[0].out_delay_inst.w35 ;
 wire \out_delay_gen[0].out_delay_inst.w36 ;
 wire \out_delay_gen[0].out_delay_inst.w37 ;
 wire \out_delay_gen[0].out_delay_inst.w38 ;
 wire \out_delay_gen[0].out_delay_inst.w39 ;
 wire \out_delay_gen[0].out_delay_inst.w4 ;
 wire \out_delay_gen[0].out_delay_inst.w5 ;
 wire \out_delay_gen[0].out_delay_inst.w6 ;
 wire \out_delay_gen[0].out_delay_inst.w7 ;
 wire \out_delay_gen[0].out_delay_inst.w8 ;
 wire \out_delay_gen[0].out_delay_inst.w9 ;
 wire \out_delay_gen[1].out_delay_inst.A ;
 wire \out_delay_gen[1].out_delay_inst.X ;
 wire \out_delay_gen[1].out_delay_inst.w1 ;
 wire \out_delay_gen[1].out_delay_inst.w10 ;
 wire \out_delay_gen[1].out_delay_inst.w11 ;
 wire \out_delay_gen[1].out_delay_inst.w12 ;
 wire \out_delay_gen[1].out_delay_inst.w13 ;
 wire \out_delay_gen[1].out_delay_inst.w14 ;
 wire \out_delay_gen[1].out_delay_inst.w15 ;
 wire \out_delay_gen[1].out_delay_inst.w16 ;
 wire \out_delay_gen[1].out_delay_inst.w17 ;
 wire \out_delay_gen[1].out_delay_inst.w18 ;
 wire \out_delay_gen[1].out_delay_inst.w19 ;
 wire \out_delay_gen[1].out_delay_inst.w2 ;
 wire \out_delay_gen[1].out_delay_inst.w20 ;
 wire \out_delay_gen[1].out_delay_inst.w21 ;
 wire \out_delay_gen[1].out_delay_inst.w22 ;
 wire \out_delay_gen[1].out_delay_inst.w23 ;
 wire \out_delay_gen[1].out_delay_inst.w24 ;
 wire \out_delay_gen[1].out_delay_inst.w25 ;
 wire \out_delay_gen[1].out_delay_inst.w26 ;
 wire \out_delay_gen[1].out_delay_inst.w27 ;
 wire \out_delay_gen[1].out_delay_inst.w28 ;
 wire \out_delay_gen[1].out_delay_inst.w29 ;
 wire \out_delay_gen[1].out_delay_inst.w3 ;
 wire \out_delay_gen[1].out_delay_inst.w30 ;
 wire \out_delay_gen[1].out_delay_inst.w31 ;
 wire \out_delay_gen[1].out_delay_inst.w32 ;
 wire \out_delay_gen[1].out_delay_inst.w33 ;
 wire \out_delay_gen[1].out_delay_inst.w34 ;
 wire \out_delay_gen[1].out_delay_inst.w35 ;
 wire \out_delay_gen[1].out_delay_inst.w36 ;
 wire \out_delay_gen[1].out_delay_inst.w37 ;
 wire \out_delay_gen[1].out_delay_inst.w38 ;
 wire \out_delay_gen[1].out_delay_inst.w39 ;
 wire \out_delay_gen[1].out_delay_inst.w4 ;
 wire \out_delay_gen[1].out_delay_inst.w5 ;
 wire \out_delay_gen[1].out_delay_inst.w6 ;
 wire \out_delay_gen[1].out_delay_inst.w7 ;
 wire \out_delay_gen[1].out_delay_inst.w8 ;
 wire \out_delay_gen[1].out_delay_inst.w9 ;
 wire \out_delay_gen[2].out_delay_inst.A ;
 wire \out_delay_gen[2].out_delay_inst.X ;
 wire \out_delay_gen[2].out_delay_inst.w1 ;
 wire \out_delay_gen[2].out_delay_inst.w10 ;
 wire \out_delay_gen[2].out_delay_inst.w11 ;
 wire \out_delay_gen[2].out_delay_inst.w12 ;
 wire \out_delay_gen[2].out_delay_inst.w13 ;
 wire \out_delay_gen[2].out_delay_inst.w14 ;
 wire \out_delay_gen[2].out_delay_inst.w15 ;
 wire \out_delay_gen[2].out_delay_inst.w16 ;
 wire \out_delay_gen[2].out_delay_inst.w17 ;
 wire \out_delay_gen[2].out_delay_inst.w18 ;
 wire \out_delay_gen[2].out_delay_inst.w19 ;
 wire \out_delay_gen[2].out_delay_inst.w2 ;
 wire \out_delay_gen[2].out_delay_inst.w20 ;
 wire \out_delay_gen[2].out_delay_inst.w21 ;
 wire \out_delay_gen[2].out_delay_inst.w22 ;
 wire \out_delay_gen[2].out_delay_inst.w23 ;
 wire \out_delay_gen[2].out_delay_inst.w24 ;
 wire \out_delay_gen[2].out_delay_inst.w25 ;
 wire \out_delay_gen[2].out_delay_inst.w26 ;
 wire \out_delay_gen[2].out_delay_inst.w27 ;
 wire \out_delay_gen[2].out_delay_inst.w28 ;
 wire \out_delay_gen[2].out_delay_inst.w29 ;
 wire \out_delay_gen[2].out_delay_inst.w3 ;
 wire \out_delay_gen[2].out_delay_inst.w30 ;
 wire \out_delay_gen[2].out_delay_inst.w31 ;
 wire \out_delay_gen[2].out_delay_inst.w32 ;
 wire \out_delay_gen[2].out_delay_inst.w33 ;
 wire \out_delay_gen[2].out_delay_inst.w34 ;
 wire \out_delay_gen[2].out_delay_inst.w35 ;
 wire \out_delay_gen[2].out_delay_inst.w36 ;
 wire \out_delay_gen[2].out_delay_inst.w37 ;
 wire \out_delay_gen[2].out_delay_inst.w38 ;
 wire \out_delay_gen[2].out_delay_inst.w39 ;
 wire \out_delay_gen[2].out_delay_inst.w4 ;
 wire \out_delay_gen[2].out_delay_inst.w5 ;
 wire \out_delay_gen[2].out_delay_inst.w6 ;
 wire \out_delay_gen[2].out_delay_inst.w7 ;
 wire \out_delay_gen[2].out_delay_inst.w8 ;
 wire \out_delay_gen[2].out_delay_inst.w9 ;
 wire \out_delay_gen[3].out_delay_inst.A ;
 wire \out_delay_gen[3].out_delay_inst.X ;
 wire \out_delay_gen[3].out_delay_inst.w1 ;
 wire \out_delay_gen[3].out_delay_inst.w10 ;
 wire \out_delay_gen[3].out_delay_inst.w11 ;
 wire \out_delay_gen[3].out_delay_inst.w12 ;
 wire \out_delay_gen[3].out_delay_inst.w13 ;
 wire \out_delay_gen[3].out_delay_inst.w14 ;
 wire \out_delay_gen[3].out_delay_inst.w15 ;
 wire \out_delay_gen[3].out_delay_inst.w16 ;
 wire \out_delay_gen[3].out_delay_inst.w17 ;
 wire \out_delay_gen[3].out_delay_inst.w18 ;
 wire \out_delay_gen[3].out_delay_inst.w19 ;
 wire \out_delay_gen[3].out_delay_inst.w2 ;
 wire \out_delay_gen[3].out_delay_inst.w20 ;
 wire \out_delay_gen[3].out_delay_inst.w21 ;
 wire \out_delay_gen[3].out_delay_inst.w22 ;
 wire \out_delay_gen[3].out_delay_inst.w23 ;
 wire \out_delay_gen[3].out_delay_inst.w24 ;
 wire \out_delay_gen[3].out_delay_inst.w25 ;
 wire \out_delay_gen[3].out_delay_inst.w26 ;
 wire \out_delay_gen[3].out_delay_inst.w27 ;
 wire \out_delay_gen[3].out_delay_inst.w28 ;
 wire \out_delay_gen[3].out_delay_inst.w29 ;
 wire \out_delay_gen[3].out_delay_inst.w3 ;
 wire \out_delay_gen[3].out_delay_inst.w30 ;
 wire \out_delay_gen[3].out_delay_inst.w31 ;
 wire \out_delay_gen[3].out_delay_inst.w32 ;
 wire \out_delay_gen[3].out_delay_inst.w33 ;
 wire \out_delay_gen[3].out_delay_inst.w34 ;
 wire \out_delay_gen[3].out_delay_inst.w35 ;
 wire \out_delay_gen[3].out_delay_inst.w36 ;
 wire \out_delay_gen[3].out_delay_inst.w37 ;
 wire \out_delay_gen[3].out_delay_inst.w38 ;
 wire \out_delay_gen[3].out_delay_inst.w39 ;
 wire \out_delay_gen[3].out_delay_inst.w4 ;
 wire \out_delay_gen[3].out_delay_inst.w5 ;
 wire \out_delay_gen[3].out_delay_inst.w6 ;
 wire \out_delay_gen[3].out_delay_inst.w7 ;
 wire \out_delay_gen[3].out_delay_inst.w8 ;
 wire \out_delay_gen[3].out_delay_inst.w9 ;
 wire \out_delay_gen[4].out_delay_inst.A ;
 wire \out_delay_gen[4].out_delay_inst.X ;
 wire \out_delay_gen[4].out_delay_inst.w1 ;
 wire \out_delay_gen[4].out_delay_inst.w10 ;
 wire \out_delay_gen[4].out_delay_inst.w11 ;
 wire \out_delay_gen[4].out_delay_inst.w12 ;
 wire \out_delay_gen[4].out_delay_inst.w13 ;
 wire \out_delay_gen[4].out_delay_inst.w14 ;
 wire \out_delay_gen[4].out_delay_inst.w15 ;
 wire \out_delay_gen[4].out_delay_inst.w16 ;
 wire \out_delay_gen[4].out_delay_inst.w17 ;
 wire \out_delay_gen[4].out_delay_inst.w18 ;
 wire \out_delay_gen[4].out_delay_inst.w19 ;
 wire \out_delay_gen[4].out_delay_inst.w2 ;
 wire \out_delay_gen[4].out_delay_inst.w20 ;
 wire \out_delay_gen[4].out_delay_inst.w21 ;
 wire \out_delay_gen[4].out_delay_inst.w22 ;
 wire \out_delay_gen[4].out_delay_inst.w23 ;
 wire \out_delay_gen[4].out_delay_inst.w24 ;
 wire \out_delay_gen[4].out_delay_inst.w25 ;
 wire \out_delay_gen[4].out_delay_inst.w26 ;
 wire \out_delay_gen[4].out_delay_inst.w27 ;
 wire \out_delay_gen[4].out_delay_inst.w28 ;
 wire \out_delay_gen[4].out_delay_inst.w29 ;
 wire \out_delay_gen[4].out_delay_inst.w3 ;
 wire \out_delay_gen[4].out_delay_inst.w30 ;
 wire \out_delay_gen[4].out_delay_inst.w31 ;
 wire \out_delay_gen[4].out_delay_inst.w32 ;
 wire \out_delay_gen[4].out_delay_inst.w33 ;
 wire \out_delay_gen[4].out_delay_inst.w34 ;
 wire \out_delay_gen[4].out_delay_inst.w35 ;
 wire \out_delay_gen[4].out_delay_inst.w36 ;
 wire \out_delay_gen[4].out_delay_inst.w37 ;
 wire \out_delay_gen[4].out_delay_inst.w38 ;
 wire \out_delay_gen[4].out_delay_inst.w39 ;
 wire \out_delay_gen[4].out_delay_inst.w4 ;
 wire \out_delay_gen[4].out_delay_inst.w5 ;
 wire \out_delay_gen[4].out_delay_inst.w6 ;
 wire \out_delay_gen[4].out_delay_inst.w7 ;
 wire \out_delay_gen[4].out_delay_inst.w8 ;
 wire \out_delay_gen[4].out_delay_inst.w9 ;
 wire \out_delay_gen[5].out_delay_inst.A ;
 wire \out_delay_gen[5].out_delay_inst.X ;
 wire \out_delay_gen[5].out_delay_inst.w1 ;
 wire \out_delay_gen[5].out_delay_inst.w10 ;
 wire \out_delay_gen[5].out_delay_inst.w11 ;
 wire \out_delay_gen[5].out_delay_inst.w12 ;
 wire \out_delay_gen[5].out_delay_inst.w13 ;
 wire \out_delay_gen[5].out_delay_inst.w14 ;
 wire \out_delay_gen[5].out_delay_inst.w15 ;
 wire \out_delay_gen[5].out_delay_inst.w16 ;
 wire \out_delay_gen[5].out_delay_inst.w17 ;
 wire \out_delay_gen[5].out_delay_inst.w18 ;
 wire \out_delay_gen[5].out_delay_inst.w19 ;
 wire \out_delay_gen[5].out_delay_inst.w2 ;
 wire \out_delay_gen[5].out_delay_inst.w20 ;
 wire \out_delay_gen[5].out_delay_inst.w21 ;
 wire \out_delay_gen[5].out_delay_inst.w22 ;
 wire \out_delay_gen[5].out_delay_inst.w23 ;
 wire \out_delay_gen[5].out_delay_inst.w24 ;
 wire \out_delay_gen[5].out_delay_inst.w25 ;
 wire \out_delay_gen[5].out_delay_inst.w26 ;
 wire \out_delay_gen[5].out_delay_inst.w27 ;
 wire \out_delay_gen[5].out_delay_inst.w28 ;
 wire \out_delay_gen[5].out_delay_inst.w29 ;
 wire \out_delay_gen[5].out_delay_inst.w3 ;
 wire \out_delay_gen[5].out_delay_inst.w30 ;
 wire \out_delay_gen[5].out_delay_inst.w31 ;
 wire \out_delay_gen[5].out_delay_inst.w32 ;
 wire \out_delay_gen[5].out_delay_inst.w33 ;
 wire \out_delay_gen[5].out_delay_inst.w34 ;
 wire \out_delay_gen[5].out_delay_inst.w35 ;
 wire \out_delay_gen[5].out_delay_inst.w36 ;
 wire \out_delay_gen[5].out_delay_inst.w37 ;
 wire \out_delay_gen[5].out_delay_inst.w38 ;
 wire \out_delay_gen[5].out_delay_inst.w39 ;
 wire \out_delay_gen[5].out_delay_inst.w4 ;
 wire \out_delay_gen[5].out_delay_inst.w5 ;
 wire \out_delay_gen[5].out_delay_inst.w6 ;
 wire \out_delay_gen[5].out_delay_inst.w7 ;
 wire \out_delay_gen[5].out_delay_inst.w8 ;
 wire \out_delay_gen[5].out_delay_inst.w9 ;
 wire \out_delay_gen[6].out_delay_inst.A ;
 wire \out_delay_gen[6].out_delay_inst.X ;
 wire \out_delay_gen[6].out_delay_inst.w1 ;
 wire \out_delay_gen[6].out_delay_inst.w10 ;
 wire \out_delay_gen[6].out_delay_inst.w11 ;
 wire \out_delay_gen[6].out_delay_inst.w12 ;
 wire \out_delay_gen[6].out_delay_inst.w13 ;
 wire \out_delay_gen[6].out_delay_inst.w14 ;
 wire \out_delay_gen[6].out_delay_inst.w15 ;
 wire \out_delay_gen[6].out_delay_inst.w16 ;
 wire \out_delay_gen[6].out_delay_inst.w17 ;
 wire \out_delay_gen[6].out_delay_inst.w18 ;
 wire \out_delay_gen[6].out_delay_inst.w19 ;
 wire \out_delay_gen[6].out_delay_inst.w2 ;
 wire \out_delay_gen[6].out_delay_inst.w20 ;
 wire \out_delay_gen[6].out_delay_inst.w21 ;
 wire \out_delay_gen[6].out_delay_inst.w22 ;
 wire \out_delay_gen[6].out_delay_inst.w23 ;
 wire \out_delay_gen[6].out_delay_inst.w24 ;
 wire \out_delay_gen[6].out_delay_inst.w25 ;
 wire \out_delay_gen[6].out_delay_inst.w26 ;
 wire \out_delay_gen[6].out_delay_inst.w27 ;
 wire \out_delay_gen[6].out_delay_inst.w28 ;
 wire \out_delay_gen[6].out_delay_inst.w29 ;
 wire \out_delay_gen[6].out_delay_inst.w3 ;
 wire \out_delay_gen[6].out_delay_inst.w30 ;
 wire \out_delay_gen[6].out_delay_inst.w31 ;
 wire \out_delay_gen[6].out_delay_inst.w32 ;
 wire \out_delay_gen[6].out_delay_inst.w33 ;
 wire \out_delay_gen[6].out_delay_inst.w34 ;
 wire \out_delay_gen[6].out_delay_inst.w35 ;
 wire \out_delay_gen[6].out_delay_inst.w36 ;
 wire \out_delay_gen[6].out_delay_inst.w37 ;
 wire \out_delay_gen[6].out_delay_inst.w38 ;
 wire \out_delay_gen[6].out_delay_inst.w39 ;
 wire \out_delay_gen[6].out_delay_inst.w4 ;
 wire \out_delay_gen[6].out_delay_inst.w5 ;
 wire \out_delay_gen[6].out_delay_inst.w6 ;
 wire \out_delay_gen[6].out_delay_inst.w7 ;
 wire \out_delay_gen[6].out_delay_inst.w8 ;
 wire \out_delay_gen[6].out_delay_inst.w9 ;
 wire \out_delay_gen[7].out_delay_inst.A ;
 wire \out_delay_gen[7].out_delay_inst.X ;
 wire \out_delay_gen[7].out_delay_inst.w1 ;
 wire \out_delay_gen[7].out_delay_inst.w10 ;
 wire \out_delay_gen[7].out_delay_inst.w11 ;
 wire \out_delay_gen[7].out_delay_inst.w12 ;
 wire \out_delay_gen[7].out_delay_inst.w13 ;
 wire \out_delay_gen[7].out_delay_inst.w14 ;
 wire \out_delay_gen[7].out_delay_inst.w15 ;
 wire \out_delay_gen[7].out_delay_inst.w16 ;
 wire \out_delay_gen[7].out_delay_inst.w17 ;
 wire \out_delay_gen[7].out_delay_inst.w18 ;
 wire \out_delay_gen[7].out_delay_inst.w19 ;
 wire \out_delay_gen[7].out_delay_inst.w2 ;
 wire \out_delay_gen[7].out_delay_inst.w20 ;
 wire \out_delay_gen[7].out_delay_inst.w21 ;
 wire \out_delay_gen[7].out_delay_inst.w22 ;
 wire \out_delay_gen[7].out_delay_inst.w23 ;
 wire \out_delay_gen[7].out_delay_inst.w24 ;
 wire \out_delay_gen[7].out_delay_inst.w25 ;
 wire \out_delay_gen[7].out_delay_inst.w26 ;
 wire \out_delay_gen[7].out_delay_inst.w27 ;
 wire \out_delay_gen[7].out_delay_inst.w28 ;
 wire \out_delay_gen[7].out_delay_inst.w29 ;
 wire \out_delay_gen[7].out_delay_inst.w3 ;
 wire \out_delay_gen[7].out_delay_inst.w30 ;
 wire \out_delay_gen[7].out_delay_inst.w31 ;
 wire \out_delay_gen[7].out_delay_inst.w32 ;
 wire \out_delay_gen[7].out_delay_inst.w33 ;
 wire \out_delay_gen[7].out_delay_inst.w34 ;
 wire \out_delay_gen[7].out_delay_inst.w35 ;
 wire \out_delay_gen[7].out_delay_inst.w36 ;
 wire \out_delay_gen[7].out_delay_inst.w37 ;
 wire \out_delay_gen[7].out_delay_inst.w38 ;
 wire \out_delay_gen[7].out_delay_inst.w39 ;
 wire \out_delay_gen[7].out_delay_inst.w4 ;
 wire \out_delay_gen[7].out_delay_inst.w5 ;
 wire \out_delay_gen[7].out_delay_inst.w6 ;
 wire \out_delay_gen[7].out_delay_inst.w7 ;
 wire \out_delay_gen[7].out_delay_inst.w8 ;
 wire \out_delay_gen[7].out_delay_inst.w9 ;
 wire processing_dly;
 wire \rst_delay.X ;
 wire \rst_delay.w1 ;
 wire \rst_delay.w10 ;
 wire \rst_delay.w11 ;
 wire \rst_delay.w12 ;
 wire \rst_delay.w13 ;
 wire \rst_delay.w14 ;
 wire \rst_delay.w15 ;
 wire \rst_delay.w16 ;
 wire \rst_delay.w17 ;
 wire \rst_delay.w18 ;
 wire \rst_delay.w19 ;
 wire \rst_delay.w2 ;
 wire \rst_delay.w20 ;
 wire \rst_delay.w21 ;
 wire \rst_delay.w22 ;
 wire \rst_delay.w23 ;
 wire \rst_delay.w24 ;
 wire \rst_delay.w25 ;
 wire \rst_delay.w26 ;
 wire \rst_delay.w27 ;
 wire \rst_delay.w28 ;
 wire \rst_delay.w29 ;
 wire \rst_delay.w3 ;
 wire \rst_delay.w30 ;
 wire \rst_delay.w31 ;
 wire \rst_delay.w32 ;
 wire \rst_delay.w33 ;
 wire \rst_delay.w34 ;
 wire \rst_delay.w35 ;
 wire \rst_delay.w36 ;
 wire \rst_delay.w37 ;
 wire \rst_delay.w38 ;
 wire \rst_delay.w39 ;
 wire \rst_delay.w4 ;
 wire \rst_delay.w5 ;
 wire \rst_delay.w6 ;
 wire \rst_delay.w7 ;
 wire \rst_delay.w8 ;
 wire \rst_delay.w9 ;
 wire rst_sync1;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.A ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[0].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[1].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[2].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[3].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[4].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[5].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[6].uio_oe_delay_inst.w9 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.X ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w1 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w10 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w11 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w12 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w13 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w14 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w15 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w16 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w17 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w18 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w19 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w2 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w20 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w21 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w22 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w23 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w24 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w25 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w26 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w27 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w28 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w29 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w3 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w30 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w31 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w32 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w33 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w34 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w35 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w36 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w37 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w38 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w39 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w4 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w5 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w6 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w7 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w8 ;
 wire \uio_oe_delay_gen[7].uio_oe_delay_inst.w9 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.X ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[0].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.A ;
 wire \uo_out_delay_gen[1].uo_delay_inst.X ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[1].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.A ;
 wire \uo_out_delay_gen[2].uo_delay_inst.X ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[2].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.A ;
 wire \uo_out_delay_gen[3].uo_delay_inst.X ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[3].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.A ;
 wire \uo_out_delay_gen[4].uo_delay_inst.X ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[4].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.A ;
 wire \uo_out_delay_gen[5].uo_delay_inst.X ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[5].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.A ;
 wire \uo_out_delay_gen[6].uo_delay_inst.X ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[6].uo_delay_inst.w9 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.X ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w1 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w10 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w11 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w12 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w13 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w14 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w15 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w16 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w17 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w18 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w19 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w2 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w20 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w21 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w22 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w23 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w24 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w25 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w26 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w27 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w28 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w29 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w3 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w30 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w31 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w32 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w33 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w34 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w35 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w36 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w37 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w38 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w39 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w4 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w5 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w6 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w7 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w8 ;
 wire \uo_out_delay_gen[7].uo_delay_inst.w9 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;

 sky130_fd_sc_hd__inv_2 _377_ (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_160_));
 sky130_fd_sc_hd__inv_2 _378_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_161_));
 sky130_fd_sc_hd__inv_2 _379_ (.A(\fft_inst.bfly_stage1_1.A_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_162_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_163_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(\fft3_imag[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_164_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_016_));
 sky130_fd_sc_hd__and3b_2 _383_ (.A_N(\io_inst.prev_in0 ),
    .B(net2),
    .C(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_165_));
 sky130_fd_sc_hd__or2_1 _384_ (.A(\addr[1] ),
    .B(\addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_166_));
 sky130_fd_sc_hd__or3b_4 _385_ (.A(\addr[1] ),
    .B(\addr[0] ),
    .C_N(_165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(net7),
    .A1(net59),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_159_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(net6),
    .A1(\fft_inst.bfly_stage1_0.A_imag[6] ),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _388_ (.A0(net5),
    .A1(\fft_inst.bfly_stage1_0.A_imag[5] ),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(net4),
    .A1(net69),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_156_));
 sky130_fd_sc_hd__nand2_1 _390_ (.A(\addr[0] ),
    .B(_165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _391_ (.A(\addr[1] ),
    .B(\addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_169_));
 sky130_fd_sc_hd__nand3_4 _392_ (.A(\addr[1] ),
    .B(\addr[0] ),
    .C(_165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_170_));
 sky130_fd_sc_hd__mux2_1 _393_ (.A0(net7),
    .A1(net57),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_155_));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(net6),
    .A1(net56),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(net5),
    .A1(\fft_inst.bfly_stage1_1.B_imag[5] ),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(net4),
    .A1(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(net47),
    .A1(net3),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_151_));
 sky130_fd_sc_hd__nor2_4 _398_ (.A(\addr[1] ),
    .B(_168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_171_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(net52),
    .A1(net11),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_150_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(net66),
    .A1(net10),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(\fft_inst.bfly_stage1_1.A_real[5] ),
    .A1(net9),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\fft_inst.bfly_stage1_1.A_real[4] ),
    .A1(net8),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(net51),
    .A1(net7),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _404_ (.A0(net68),
    .A1(net6),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(\fft_inst.bfly_stage1_1.A_imag[5] ),
    .A1(net5),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(\fft_inst.bfly_stage1_1.A_imag[4] ),
    .A1(net4),
    .S(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_143_));
 sky130_fd_sc_hd__and3b_4 _407_ (.A_N(\addr[0] ),
    .B(_165_),
    .C(\addr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(net50),
    .A1(net11),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _409_ (.A0(net48),
    .A1(net10),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(\fft_inst.bfly_stage1_0.B_real[5] ),
    .A1(net9),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_140_));
 sky130_fd_sc_hd__mux2_1 _411_ (.A0(\fft_inst.bfly_stage1_0.B_real[4] ),
    .A1(net8),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _412_ (.A0(net11),
    .A1(net53),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _413_ (.A0(net10),
    .A1(net61),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(net9),
    .A1(\fft_inst.bfly_stage1_1.B_real[5] ),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(net8),
    .A1(\fft_inst.bfly_stage1_1.B_real[4] ),
    .S(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _416_ (.A0(net49),
    .A1(net7),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(net58),
    .A1(net6),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _418_ (.A0(\fft_inst.bfly_stage1_0.B_imag[5] ),
    .A1(net5),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .A1(net4),
    .S(_172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _420_ (.A0(net36),
    .A1(net2),
    .S(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(net11),
    .A1(net60),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _422_ (.A0(net10),
    .A1(\fft_inst.bfly_stage1_0.A_real[6] ),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(net9),
    .A1(\fft_inst.bfly_stage1_0.A_real[5] ),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(net8),
    .A1(net70),
    .S(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_126_));
 sky130_fd_sc_hd__and2_1 _425_ (.A(\addr[1] ),
    .B(_168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_173_));
 sky130_fd_sc_hd__or2_1 _426_ (.A(_171_),
    .B(_173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_125_));
 sky130_fd_sc_hd__or2_1 _427_ (.A(\addr[0] ),
    .B(_165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_174_));
 sky130_fd_sc_hd__and2_1 _428_ (.A(_168_),
    .B(_174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_124_));
 sky130_fd_sc_hd__nor2_2 _429_ (.A(net27),
    .B(\disp_inst.processing ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_175_));
 sky130_fd_sc_hd__o21ba_1 _430_ (.A1(net29),
    .A2(net40),
    .B1_N(_175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_123_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(net24),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_176_));
 sky130_fd_sc_hd__or4_1 _432_ (.A(\io_inst.prev_in1 ),
    .B(_160_),
    .C(net27),
    .D(_176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_177_));
 sky130_fd_sc_hd__a22o_1 _433_ (.A1(net40),
    .A2(_175_),
    .B1(_177_),
    .B2(\disp_inst.done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_122_));
 sky130_fd_sc_hd__a21bo_1 _434_ (.A1(_161_),
    .A2(net45),
    .B1_N(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_121_));
 sky130_fd_sc_hd__and3_1 _435_ (.A(net24),
    .B(net25),
    .C(\fft3_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_178_));
 sky130_fd_sc_hd__and2_1 _436_ (.A(_163_),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_179_));
 sky130_fd_sc_hd__nor2_2 _437_ (.A(_163_),
    .B(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_180_));
 sky130_fd_sc_hd__a221o_1 _438_ (.A1(\fft1_real[7] ),
    .A2(_179_),
    .B1(_180_),
    .B2(\fft2_real[7] ),
    .C1(_178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_181_));
 sky130_fd_sc_hd__nor2_2 _439_ (.A(net24),
    .B(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_182_));
 sky130_fd_sc_hd__a21o_1 _440_ (.A1(net64),
    .A2(_182_),
    .B1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_183_));
 sky130_fd_sc_hd__o22a_1 _441_ (.A1(net28),
    .A2(\out_delay_gen[7].out_delay_inst.A ),
    .B1(_181_),
    .B2(_183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_120_));
 sky130_fd_sc_hd__a221o_1 _442_ (.A1(_163_),
    .A2(\fft1_real[6] ),
    .B1(_180_),
    .B2(\fft2_real[6] ),
    .C1(_182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_184_));
 sky130_fd_sc_hd__a31o_1 _443_ (.A1(net24),
    .A2(net25),
    .A3(\fft3_real[6] ),
    .B1(_184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_185_));
 sky130_fd_sc_hd__o31a_1 _444_ (.A1(net24),
    .A2(net25),
    .A3(\fft0_real[6] ),
    .B1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_186_));
 sky130_fd_sc_hd__a22o_1 _445_ (.A1(net27),
    .A2(net67),
    .B1(_185_),
    .B2(_186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_119_));
 sky130_fd_sc_hd__a21o_1 _446_ (.A1(\fft0_real[5] ),
    .A2(_182_),
    .B1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_187_));
 sky130_fd_sc_hd__and3_1 _447_ (.A(net24),
    .B(net25),
    .C(\fft3_real[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_188_));
 sky130_fd_sc_hd__a221o_1 _448_ (.A1(\fft1_real[5] ),
    .A2(_179_),
    .B1(_180_),
    .B2(\fft2_real[5] ),
    .C1(_188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_189_));
 sky130_fd_sc_hd__o22a_1 _449_ (.A1(net28),
    .A2(net63),
    .B1(_187_),
    .B2(_189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_118_));
 sky130_fd_sc_hd__mux4_1 _450_ (.A0(\fft0_real[4] ),
    .A1(\fft1_real[4] ),
    .A2(\fft2_real[4] ),
    .A3(\fft3_real[4] ),
    .S0(net25),
    .S1(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_190_));
 sky130_fd_sc_hd__mux2_1 _451_ (.A0(net54),
    .A1(_190_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_117_));
 sky130_fd_sc_hd__mux4_1 _452_ (.A0(\fft0_imag[7] ),
    .A1(\fft1_imag[7] ),
    .A2(\fft2_imag[7] ),
    .A3(\fft3_imag[7] ),
    .S0(net26),
    .S1(\disp_inst.output_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_191_));
 sky130_fd_sc_hd__mux2_1 _453_ (.A0(net37),
    .A1(_191_),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_116_));
 sky130_fd_sc_hd__and3_1 _454_ (.A(\disp_inst.output_counter[1] ),
    .B(net26),
    .C(\fft3_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_192_));
 sky130_fd_sc_hd__a221o_1 _455_ (.A1(\fft1_imag[6] ),
    .A2(_179_),
    .B1(_180_),
    .B2(\fft2_imag[6] ),
    .C1(_192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_193_));
 sky130_fd_sc_hd__a21o_1 _456_ (.A1(\fft0_imag[6] ),
    .A2(_182_),
    .B1(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_194_));
 sky130_fd_sc_hd__o22a_1 _457_ (.A1(net29),
    .A2(net42),
    .B1(_193_),
    .B2(_194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_115_));
 sky130_fd_sc_hd__a2bb2o_1 _458_ (.A1_N(_164_),
    .A2_N(_176_),
    .B1(\fft1_imag[5] ),
    .B2(_163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_195_));
 sky130_fd_sc_hd__a211o_1 _459_ (.A1(\fft2_imag[5] ),
    .A2(_180_),
    .B1(_182_),
    .C1(_195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_196_));
 sky130_fd_sc_hd__o31a_1 _460_ (.A1(net24),
    .A2(net26),
    .A3(\fft0_imag[5] ),
    .B1(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_197_));
 sky130_fd_sc_hd__a22o_1 _461_ (.A1(_161_),
    .A2(net55),
    .B1(_196_),
    .B2(_197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_114_));
 sky130_fd_sc_hd__mux4_1 _462_ (.A0(\fft0_imag[4] ),
    .A1(\fft1_imag[4] ),
    .A2(\fft2_imag[4] ),
    .A3(\fft3_imag[4] ),
    .S0(net25),
    .S1(\disp_inst.output_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_198_));
 sky130_fd_sc_hd__mux2_1 _463_ (.A0(net62),
    .A1(_198_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_113_));
 sky130_fd_sc_hd__and4b_1 _464_ (.A_N(\io_inst.prev_in1 ),
    .B(net3),
    .C(net29),
    .D(\disp_inst.done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_199_));
 sky130_fd_sc_hd__a21o_1 _465_ (.A1(net27),
    .A2(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .B1(_199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_112_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(net25),
    .B(_199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_200_));
 sky130_fd_sc_hd__xnor2_1 _467_ (.A(net24),
    .B(_200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_111_));
 sky130_fd_sc_hd__or2_1 _468_ (.A(net25),
    .B(_199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_201_));
 sky130_fd_sc_hd__and2_1 _469_ (.A(_200_),
    .B(_201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_110_));
 sky130_fd_sc_hd__nand2_1 _470_ (.A(\disp_inst.done ),
    .B(_180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_202_));
 sky130_fd_sc_hd__a21o_1 _471_ (.A1(_166_),
    .A2(_169_),
    .B1(\disp_inst.done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_203_));
 sky130_fd_sc_hd__a32o_1 _472_ (.A1(_175_),
    .A2(_202_),
    .A3(_203_),
    .B1(net39),
    .B2(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_109_));
 sky130_fd_sc_hd__o21ai_1 _473_ (.A1(_163_),
    .A2(net25),
    .B1(\disp_inst.done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_204_));
 sky130_fd_sc_hd__o2bb2a_1 _474_ (.A1_N(_175_),
    .A2_N(_204_),
    .B1(net28),
    .B2(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_108_));
 sky130_fd_sc_hd__nand2_1 _475_ (.A(\addr[1] ),
    .B(_175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_205_));
 sky130_fd_sc_hd__nand2b_1 _476_ (.A_N(\disp_inst.done ),
    .B(\addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_206_));
 sky130_fd_sc_hd__nand2_1 _477_ (.A(_175_),
    .B(_206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_207_));
 sky130_fd_sc_hd__a22o_1 _478_ (.A1(\disp_inst.done ),
    .A2(_179_),
    .B1(_205_),
    .B2(_207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_208_));
 sky130_fd_sc_hd__o21a_1 _479_ (.A1(net28),
    .A2(net35),
    .B1(_208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_107_));
 sky130_fd_sc_hd__o22a_1 _480_ (.A1(net28),
    .A2(net41),
    .B1(_205_),
    .B2(_206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_106_));
 sky130_fd_sc_hd__a22o_1 _481_ (.A1(net27),
    .A2(net44),
    .B1(_175_),
    .B2(_206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_105_));
 sky130_fd_sc_hd__a32o_1 _482_ (.A1(_175_),
    .A2(_203_),
    .A3(_204_),
    .B1(net38),
    .B2(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_104_));
 sky130_fd_sc_hd__nand2b_2 _483_ (.A_N(\fft_inst.bfly_stage1_0.A_imag[4] ),
    .B(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_209_));
 sky130_fd_sc_hd__nand2b_1 _484_ (.A_N(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .B(\fft_inst.bfly_stage1_0.A_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_210_));
 sky130_fd_sc_hd__nand2_2 _485_ (.A(_209_),
    .B(_210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_211_));
 sky130_fd_sc_hd__nand2_2 _486_ (.A(\fft_inst.bfly_stage1_1.A_real[4] ),
    .B(\fft_inst.bfly_stage1_1.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_212_));
 sky130_fd_sc_hd__or2_1 _487_ (.A(\fft_inst.bfly_stage1_1.A_real[4] ),
    .B(\fft_inst.bfly_stage1_1.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_213_));
 sky130_fd_sc_hd__nand2_4 _488_ (.A(_212_),
    .B(_213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_214_));
 sky130_fd_sc_hd__nand2b_1 _489_ (.A_N(_214_),
    .B(_211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_215_));
 sky130_fd_sc_hd__xnor2_1 _490_ (.A(_211_),
    .B(_214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_neg_imag[4] ));
 sky130_fd_sc_hd__nand2b_1 _491_ (.A_N(\fft_inst.bfly_stage1_1.A_imag[4] ),
    .B(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_216_));
 sky130_fd_sc_hd__xnor2_4 _492_ (.A(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .B(\fft_inst.bfly_stage1_1.A_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_217_));
 sky130_fd_sc_hd__nand2_2 _493_ (.A(\fft_inst.bfly_stage1_0.B_real[4] ),
    .B(\fft_inst.bfly_stage1_0.A_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_218_));
 sky130_fd_sc_hd__or2_1 _494_ (.A(\fft_inst.bfly_stage1_0.B_real[4] ),
    .B(\fft_inst.bfly_stage1_0.A_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_219_));
 sky130_fd_sc_hd__and2_1 _495_ (.A(_218_),
    .B(_219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_220_));
 sky130_fd_sc_hd__nand2_2 _496_ (.A(_218_),
    .B(_219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_221_));
 sky130_fd_sc_hd__nor2_1 _497_ (.A(_217_),
    .B(_221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_222_));
 sky130_fd_sc_hd__and2_1 _498_ (.A(_217_),
    .B(_221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_223_));
 sky130_fd_sc_hd__nor2_1 _499_ (.A(_222_),
    .B(_223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_neg_real[4] ));
 sky130_fd_sc_hd__or2_2 _500_ (.A(_211_),
    .B(_217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_224_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(_211_),
    .B(_217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_225_));
 sky130_fd_sc_hd__a21oi_1 _502_ (.A1(_209_),
    .A2(_210_),
    .B1(_217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_226_));
 sky130_fd_sc_hd__inv_2 _503_ (.A(_226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_227_));
 sky130_fd_sc_hd__nand2_1 _504_ (.A(_224_),
    .B(_225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_012_));
 sky130_fd_sc_hd__or2_1 _505_ (.A(_214_),
    .B(_220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_228_));
 sky130_fd_sc_hd__nand2_1 _506_ (.A(_214_),
    .B(_220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_229_));
 sky130_fd_sc_hd__nand2_1 _507_ (.A(_228_),
    .B(_229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_004_));
 sky130_fd_sc_hd__nand2b_1 _508_ (.A_N(\fft_inst.bfly_stage1_0.A_real[4] ),
    .B(\fft_inst.bfly_stage1_0.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_230_));
 sky130_fd_sc_hd__xor2_4 _509_ (.A(\fft_inst.bfly_stage1_0.B_real[5] ),
    .B(\fft_inst.bfly_stage1_0.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_231_));
 sky130_fd_sc_hd__nand2_1 _510_ (.A(\fft_inst.bfly_stage1_0.A_real[5] ),
    .B(_231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_232_));
 sky130_fd_sc_hd__xnor2_4 _511_ (.A(\fft_inst.bfly_stage1_0.A_real[5] ),
    .B(_231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_233_));
 sky130_fd_sc_hd__xnor2_2 _512_ (.A(_230_),
    .B(_233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_234_));
 sky130_fd_sc_hd__xor2_4 _513_ (.A(\fft_inst.bfly_stage1_1.B_imag[5] ),
    .B(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_235_));
 sky130_fd_sc_hd__nand2_1 _514_ (.A(\fft_inst.bfly_stage1_1.A_imag[5] ),
    .B(_235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_236_));
 sky130_fd_sc_hd__xnor2_4 _515_ (.A(\fft_inst.bfly_stage1_1.A_imag[5] ),
    .B(_235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_237_));
 sky130_fd_sc_hd__xnor2_2 _516_ (.A(_216_),
    .B(_237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_238_));
 sky130_fd_sc_hd__and2b_1 _517_ (.A_N(_234_),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_239_));
 sky130_fd_sc_hd__xnor2_2 _518_ (.A(_234_),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_240_));
 sky130_fd_sc_hd__xnor2_1 _519_ (.A(_222_),
    .B(_240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_pos_real[5] ));
 sky130_fd_sc_hd__or2_1 _520_ (.A(_234_),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_241_));
 sky130_fd_sc_hd__o31a_1 _521_ (.A1(_217_),
    .A2(_221_),
    .A3(_240_),
    .B1(_241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_242_));
 sky130_fd_sc_hd__and2b_1 _522_ (.A_N(_231_),
    .B(\fft_inst.bfly_stage1_0.A_real[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_243_));
 sky130_fd_sc_hd__a21o_1 _523_ (.A1(_230_),
    .A2(_233_),
    .B1(_243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_244_));
 sky130_fd_sc_hd__or3_1 _524_ (.A(\fft_inst.bfly_stage1_0.B_real[6] ),
    .B(\fft_inst.bfly_stage1_0.B_real[5] ),
    .C(\fft_inst.bfly_stage1_0.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_245_));
 sky130_fd_sc_hd__o21ai_1 _525_ (.A1(\fft_inst.bfly_stage1_0.B_real[5] ),
    .A2(\fft_inst.bfly_stage1_0.B_real[4] ),
    .B1(\fft_inst.bfly_stage1_0.B_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_246_));
 sky130_fd_sc_hd__and2_2 _526_ (.A(_245_),
    .B(_246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_247_));
 sky130_fd_sc_hd__and3_1 _527_ (.A(\fft_inst.bfly_stage1_0.A_real[6] ),
    .B(_245_),
    .C(_246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_248_));
 sky130_fd_sc_hd__or2_1 _528_ (.A(\fft_inst.bfly_stage1_0.A_real[6] ),
    .B(_247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_249_));
 sky130_fd_sc_hd__and2b_1 _529_ (.A_N(_247_),
    .B(\fft_inst.bfly_stage1_0.A_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_250_));
 sky130_fd_sc_hd__xnor2_4 _530_ (.A(\fft_inst.bfly_stage1_0.A_real[6] ),
    .B(_247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_251_));
 sky130_fd_sc_hd__xnor2_2 _531_ (.A(_244_),
    .B(_251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_252_));
 sky130_fd_sc_hd__or3_2 _532_ (.A(\fft_inst.bfly_stage1_1.B_imag[6] ),
    .B(\fft_inst.bfly_stage1_1.B_imag[5] ),
    .C(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_253_));
 sky130_fd_sc_hd__o21ai_1 _533_ (.A1(\fft_inst.bfly_stage1_1.B_imag[5] ),
    .A2(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .B1(\fft_inst.bfly_stage1_1.B_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_254_));
 sky130_fd_sc_hd__and3_1 _534_ (.A(_162_),
    .B(_253_),
    .C(_254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_255_));
 sky130_fd_sc_hd__a21oi_1 _535_ (.A1(_253_),
    .A2(_254_),
    .B1(_162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_256_));
 sky130_fd_sc_hd__or2_2 _536_ (.A(_255_),
    .B(_256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_257_));
 sky130_fd_sc_hd__o21ba_1 _537_ (.A1(\fft_inst.bfly_stage1_1.A_imag[5] ),
    .A2(_216_),
    .B1_N(_235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_258_));
 sky130_fd_sc_hd__a21o_1 _538_ (.A1(\fft_inst.bfly_stage1_1.A_imag[5] ),
    .A2(_216_),
    .B1(_258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_259_));
 sky130_fd_sc_hd__xnor2_2 _539_ (.A(_257_),
    .B(_259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_260_));
 sky130_fd_sc_hd__nor2_1 _540_ (.A(_252_),
    .B(_260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_261_));
 sky130_fd_sc_hd__nand2b_1 _541_ (.A_N(_252_),
    .B(_260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_262_));
 sky130_fd_sc_hd__xor2_2 _542_ (.A(_252_),
    .B(_260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_263_));
 sky130_fd_sc_hd__xor2_1 _543_ (.A(_242_),
    .B(_263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\fft_inst.bfly_pos_real[6] ));
 sky130_fd_sc_hd__o21ai_1 _544_ (.A1(_242_),
    .A2(_263_),
    .B1(_262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_264_));
 sky130_fd_sc_hd__a21oi_1 _545_ (.A1(_244_),
    .A2(_251_),
    .B1(_250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_265_));
 sky130_fd_sc_hd__o21ba_1 _546_ (.A1(_256_),
    .A2(_259_),
    .B1_N(_255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_266_));
 sky130_fd_sc_hd__xnor2_1 _547_ (.A(\fft_inst.bfly_stage1_1.B_imag[7] ),
    .B(\fft_inst.bfly_stage1_1.A_imag[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_267_));
 sky130_fd_sc_hd__xnor2_2 _548_ (.A(_253_),
    .B(_267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_268_));
 sky130_fd_sc_hd__xnor2_1 _549_ (.A(\fft_inst.bfly_stage1_0.B_real[7] ),
    .B(\fft_inst.bfly_stage1_0.A_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_269_));
 sky130_fd_sc_hd__xnor2_1 _550_ (.A(_245_),
    .B(_269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_270_));
 sky130_fd_sc_hd__xor2_1 _551_ (.A(_268_),
    .B(_270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_271_));
 sky130_fd_sc_hd__xnor2_1 _552_ (.A(_265_),
    .B(_271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_272_));
 sky130_fd_sc_hd__xnor2_1 _553_ (.A(_266_),
    .B(_272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_273_));
 sky130_fd_sc_hd__xnor2_1 _554_ (.A(_264_),
    .B(_273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_pos_real[7] ));
 sky130_fd_sc_hd__xor2_4 _555_ (.A(\fft_inst.bfly_stage1_1.B_real[5] ),
    .B(\fft_inst.bfly_stage1_1.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_274_));
 sky130_fd_sc_hd__nand2_1 _556_ (.A(\fft_inst.bfly_stage1_1.A_real[5] ),
    .B(_274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_275_));
 sky130_fd_sc_hd__xnor2_4 _557_ (.A(\fft_inst.bfly_stage1_1.A_real[5] ),
    .B(_274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_276_));
 sky130_fd_sc_hd__nand2b_2 _558_ (.A_N(\fft_inst.bfly_stage1_1.B_real[4] ),
    .B(\fft_inst.bfly_stage1_1.A_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_277_));
 sky130_fd_sc_hd__and2_1 _559_ (.A(_276_),
    .B(_277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_278_));
 sky130_fd_sc_hd__nor2_1 _560_ (.A(_276_),
    .B(_277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_279_));
 sky130_fd_sc_hd__xor2_2 _561_ (.A(_276_),
    .B(_277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_280_));
 sky130_fd_sc_hd__xor2_4 _562_ (.A(\fft_inst.bfly_stage1_0.B_imag[5] ),
    .B(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_281_));
 sky130_fd_sc_hd__nand2_1 _563_ (.A(\fft_inst.bfly_stage1_0.A_imag[5] ),
    .B(_281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_282_));
 sky130_fd_sc_hd__xnor2_4 _564_ (.A(\fft_inst.bfly_stage1_0.A_imag[5] ),
    .B(_281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_283_));
 sky130_fd_sc_hd__xnor2_2 _565_ (.A(_209_),
    .B(_283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_284_));
 sky130_fd_sc_hd__nor2_1 _566_ (.A(_280_),
    .B(_284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_285_));
 sky130_fd_sc_hd__xor2_2 _567_ (.A(_280_),
    .B(_284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_286_));
 sky130_fd_sc_hd__or2_1 _568_ (.A(_211_),
    .B(_214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_287_));
 sky130_fd_sc_hd__xor2_1 _569_ (.A(_286_),
    .B(_287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\fft_inst.bfly_neg_imag[5] ));
 sky130_fd_sc_hd__a21o_1 _570_ (.A1(_286_),
    .A2(_287_),
    .B1(_285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_288_));
 sky130_fd_sc_hd__and2b_1 _571_ (.A_N(\fft_inst.bfly_stage1_1.A_real[5] ),
    .B(_274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_289_));
 sky130_fd_sc_hd__a21o_1 _572_ (.A1(_276_),
    .A2(_277_),
    .B1(_289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_290_));
 sky130_fd_sc_hd__or3_1 _573_ (.A(\fft_inst.bfly_stage1_1.B_real[6] ),
    .B(\fft_inst.bfly_stage1_1.B_real[5] ),
    .C(\fft_inst.bfly_stage1_1.B_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_291_));
 sky130_fd_sc_hd__o21ai_1 _574_ (.A1(\fft_inst.bfly_stage1_1.B_real[5] ),
    .A2(\fft_inst.bfly_stage1_1.B_real[4] ),
    .B1(\fft_inst.bfly_stage1_1.B_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_292_));
 sky130_fd_sc_hd__and3_1 _575_ (.A(\fft_inst.bfly_stage1_1.A_real[6] ),
    .B(_291_),
    .C(_292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_293_));
 sky130_fd_sc_hd__a21oi_1 _576_ (.A1(_291_),
    .A2(_292_),
    .B1(\fft_inst.bfly_stage1_1.A_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_294_));
 sky130_fd_sc_hd__and3b_1 _577_ (.A_N(\fft_inst.bfly_stage1_1.A_real[6] ),
    .B(_291_),
    .C(_292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_295_));
 sky130_fd_sc_hd__or2_2 _578_ (.A(_293_),
    .B(_294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_296_));
 sky130_fd_sc_hd__xor2_1 _579_ (.A(_290_),
    .B(_296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_297_));
 sky130_fd_sc_hd__xnor2_1 _580_ (.A(_290_),
    .B(_296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_298_));
 sky130_fd_sc_hd__and2b_1 _581_ (.A_N(_281_),
    .B(\fft_inst.bfly_stage1_0.A_imag[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_299_));
 sky130_fd_sc_hd__a21o_1 _582_ (.A1(_209_),
    .A2(_283_),
    .B1(_299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_300_));
 sky130_fd_sc_hd__or3_1 _583_ (.A(\fft_inst.bfly_stage1_0.B_imag[6] ),
    .B(\fft_inst.bfly_stage1_0.B_imag[5] ),
    .C(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_301_));
 sky130_fd_sc_hd__o21ai_1 _584_ (.A1(\fft_inst.bfly_stage1_0.B_imag[5] ),
    .A2(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .B1(\fft_inst.bfly_stage1_0.B_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_302_));
 sky130_fd_sc_hd__and2_2 _585_ (.A(_301_),
    .B(_302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_303_));
 sky130_fd_sc_hd__nand2_1 _586_ (.A(\fft_inst.bfly_stage1_0.A_imag[6] ),
    .B(_303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_304_));
 sky130_fd_sc_hd__and2b_1 _587_ (.A_N(_303_),
    .B(\fft_inst.bfly_stage1_0.A_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_305_));
 sky130_fd_sc_hd__xnor2_4 _588_ (.A(\fft_inst.bfly_stage1_0.A_imag[6] ),
    .B(_303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_306_));
 sky130_fd_sc_hd__xor2_1 _589_ (.A(_300_),
    .B(_306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_307_));
 sky130_fd_sc_hd__xnor2_1 _590_ (.A(_300_),
    .B(_306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_308_));
 sky130_fd_sc_hd__nor2_1 _591_ (.A(_297_),
    .B(_308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_309_));
 sky130_fd_sc_hd__nor2_1 _592_ (.A(_298_),
    .B(_308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_310_));
 sky130_fd_sc_hd__xnor2_1 _593_ (.A(_297_),
    .B(_307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_311_));
 sky130_fd_sc_hd__xnor2_1 _594_ (.A(_298_),
    .B(_307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_312_));
 sky130_fd_sc_hd__xnor2_1 _595_ (.A(_288_),
    .B(_312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_neg_imag[6] ));
 sky130_fd_sc_hd__a21oi_1 _596_ (.A1(_288_),
    .A2(_311_),
    .B1(_309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_313_));
 sky130_fd_sc_hd__a21oi_1 _597_ (.A1(_290_),
    .A2(_296_),
    .B1(_295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_314_));
 sky130_fd_sc_hd__a21oi_1 _598_ (.A1(_300_),
    .A2(_306_),
    .B1(_305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_315_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(_314_),
    .B(_315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_316_));
 sky130_fd_sc_hd__xnor2_1 _600_ (.A(\fft_inst.bfly_stage1_1.A_real[7] ),
    .B(\fft_inst.bfly_stage1_1.B_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_317_));
 sky130_fd_sc_hd__xnor2_1 _601_ (.A(_291_),
    .B(_317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_318_));
 sky130_fd_sc_hd__xnor2_1 _602_ (.A(\fft_inst.bfly_stage1_0.A_imag[7] ),
    .B(\fft_inst.bfly_stage1_0.B_imag[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_319_));
 sky130_fd_sc_hd__xnor2_1 _603_ (.A(_301_),
    .B(_319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_320_));
 sky130_fd_sc_hd__xnor2_1 _604_ (.A(_318_),
    .B(_320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_321_));
 sky130_fd_sc_hd__xnor2_1 _605_ (.A(_316_),
    .B(_321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_322_));
 sky130_fd_sc_hd__xnor2_1 _606_ (.A(_313_),
    .B(_322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_neg_imag[7] ));
 sky130_fd_sc_hd__xor2_1 _607_ (.A(_215_),
    .B(_286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\fft_inst.bfly_pos_imag[5] ));
 sky130_fd_sc_hd__or3_1 _608_ (.A(_278_),
    .B(_279_),
    .C(_284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_323_));
 sky130_fd_sc_hd__o21ai_1 _609_ (.A1(_215_),
    .A2(_286_),
    .B1(_323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_324_));
 sky130_fd_sc_hd__xnor2_1 _610_ (.A(_311_),
    .B(_324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_pos_imag[6] ));
 sky130_fd_sc_hd__a21o_1 _611_ (.A1(_312_),
    .A2(_324_),
    .B1(_310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_325_));
 sky130_fd_sc_hd__xnor2_1 _612_ (.A(_322_),
    .B(_325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_pos_imag[7] ));
 sky130_fd_sc_hd__or2_1 _613_ (.A(_217_),
    .B(_220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_326_));
 sky130_fd_sc_hd__xor2_1 _614_ (.A(_240_),
    .B(_326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\fft_inst.bfly_neg_real[5] ));
 sky130_fd_sc_hd__a21o_1 _615_ (.A1(_240_),
    .A2(_326_),
    .B1(_239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_327_));
 sky130_fd_sc_hd__xor2_1 _616_ (.A(_263_),
    .B(_327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\fft_inst.bfly_neg_real[6] ));
 sky130_fd_sc_hd__a21oi_1 _617_ (.A1(_263_),
    .A2(_327_),
    .B1(_261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_328_));
 sky130_fd_sc_hd__xnor2_1 _618_ (.A(_273_),
    .B(_328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_neg_real[7] ));
 sky130_fd_sc_hd__nand2_1 _619_ (.A(\fft_inst.bfly_stage1_1.B_imag[4] ),
    .B(\fft_inst.bfly_stage1_1.A_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_329_));
 sky130_fd_sc_hd__xor2_2 _620_ (.A(_237_),
    .B(_329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_330_));
 sky130_fd_sc_hd__nand2_1 _621_ (.A(\fft_inst.bfly_stage1_0.A_imag[4] ),
    .B(\fft_inst.bfly_stage1_0.B_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_331_));
 sky130_fd_sc_hd__xor2_2 _622_ (.A(_283_),
    .B(_331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_332_));
 sky130_fd_sc_hd__and2b_1 _623_ (.A_N(_330_),
    .B(_332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_333_));
 sky130_fd_sc_hd__xnor2_2 _624_ (.A(_330_),
    .B(_332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_334_));
 sky130_fd_sc_hd__xnor2_1 _625_ (.A(_226_),
    .B(_334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _626_ (.A(_330_),
    .B(_332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_335_));
 sky130_fd_sc_hd__o21ai_1 _627_ (.A1(_227_),
    .A2(_334_),
    .B1(_335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_336_));
 sky130_fd_sc_hd__o21ai_2 _628_ (.A1(_237_),
    .A2(_329_),
    .B1(_236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_337_));
 sky130_fd_sc_hd__xnor2_2 _629_ (.A(_257_),
    .B(_337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_338_));
 sky130_fd_sc_hd__o21a_1 _630_ (.A1(_283_),
    .A2(_331_),
    .B1(_282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_339_));
 sky130_fd_sc_hd__xnor2_2 _631_ (.A(_306_),
    .B(_339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_340_));
 sky130_fd_sc_hd__nor2_1 _632_ (.A(_338_),
    .B(_340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_341_));
 sky130_fd_sc_hd__nand2b_1 _633_ (.A_N(_340_),
    .B(_338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_342_));
 sky130_fd_sc_hd__xor2_2 _634_ (.A(_338_),
    .B(_340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_343_));
 sky130_fd_sc_hd__xor2_1 _635_ (.A(_336_),
    .B(_343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__a21o_1 _636_ (.A1(_336_),
    .A2(_343_),
    .B1(_341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_344_));
 sky130_fd_sc_hd__xor2_1 _637_ (.A(_268_),
    .B(_320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_345_));
 sky130_fd_sc_hd__o21a_1 _638_ (.A1(_306_),
    .A2(_339_),
    .B1(_304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_346_));
 sky130_fd_sc_hd__a32o_1 _639_ (.A1(\fft_inst.bfly_stage1_1.A_imag[6] ),
    .A2(_253_),
    .A3(_254_),
    .B1(_257_),
    .B2(_337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_347_));
 sky130_fd_sc_hd__xnor2_1 _640_ (.A(_345_),
    .B(_347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_348_));
 sky130_fd_sc_hd__xnor2_1 _641_ (.A(_346_),
    .B(_348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_349_));
 sky130_fd_sc_hd__xnor2_1 _642_ (.A(_344_),
    .B(_349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_011_));
 sky130_fd_sc_hd__xor2_1 _643_ (.A(_224_),
    .B(_334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__a21oi_1 _644_ (.A1(_224_),
    .A2(_334_),
    .B1(_333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_350_));
 sky130_fd_sc_hd__xor2_1 _645_ (.A(_343_),
    .B(_350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__o21a_1 _646_ (.A1(_343_),
    .A2(_350_),
    .B1(_342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_351_));
 sky130_fd_sc_hd__xnor2_1 _647_ (.A(_349_),
    .B(_351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_015_));
 sky130_fd_sc_hd__xor2_2 _648_ (.A(_212_),
    .B(_276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_352_));
 sky130_fd_sc_hd__xor2_2 _649_ (.A(_218_),
    .B(_233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_353_));
 sky130_fd_sc_hd__and2b_1 _650_ (.A_N(_352_),
    .B(_353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_354_));
 sky130_fd_sc_hd__xnor2_2 _651_ (.A(_352_),
    .B(_353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_355_));
 sky130_fd_sc_hd__xor2_1 _652_ (.A(_228_),
    .B(_355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__a21oi_1 _653_ (.A1(_228_),
    .A2(_355_),
    .B1(_354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_356_));
 sky130_fd_sc_hd__o21a_1 _654_ (.A1(_212_),
    .A2(_276_),
    .B1(_275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_357_));
 sky130_fd_sc_hd__xnor2_2 _655_ (.A(_296_),
    .B(_357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_358_));
 sky130_fd_sc_hd__o21ai_2 _656_ (.A1(_218_),
    .A2(_233_),
    .B1(_232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_359_));
 sky130_fd_sc_hd__xor2_2 _657_ (.A(_251_),
    .B(_359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_360_));
 sky130_fd_sc_hd__nor2_1 _658_ (.A(_358_),
    .B(_360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_361_));
 sky130_fd_sc_hd__nand2b_1 _659_ (.A_N(_360_),
    .B(_358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_362_));
 sky130_fd_sc_hd__xor2_2 _660_ (.A(_358_),
    .B(_360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_363_));
 sky130_fd_sc_hd__xor2_1 _661_ (.A(_356_),
    .B(_363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__o21ai_1 _662_ (.A1(_356_),
    .A2(_363_),
    .B1(_362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_364_));
 sky130_fd_sc_hd__o21ba_1 _663_ (.A1(_296_),
    .A2(_357_),
    .B1_N(_293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_365_));
 sky130_fd_sc_hd__xor2_1 _664_ (.A(_270_),
    .B(_318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_366_));
 sky130_fd_sc_hd__a21oi_1 _665_ (.A1(_249_),
    .A2(_359_),
    .B1(_248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_367_));
 sky130_fd_sc_hd__xnor2_1 _666_ (.A(_366_),
    .B(_367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_368_));
 sky130_fd_sc_hd__xnor2_1 _667_ (.A(_365_),
    .B(_368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_369_));
 sky130_fd_sc_hd__xnor2_1 _668_ (.A(_364_),
    .B(_369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_1 _669_ (.A(_214_),
    .B(_221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_370_));
 sky130_fd_sc_hd__xnor2_1 _670_ (.A(_355_),
    .B(_370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _671_ (.A(_352_),
    .B(_353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_371_));
 sky130_fd_sc_hd__o31ai_2 _672_ (.A1(_214_),
    .A2(_221_),
    .A3(_355_),
    .B1(_371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_372_));
 sky130_fd_sc_hd__xor2_1 _673_ (.A(_363_),
    .B(_372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__a21oi_1 _674_ (.A1(_363_),
    .A2(_372_),
    .B1(_361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_373_));
 sky130_fd_sc_hd__xnor2_1 _675_ (.A(_369_),
    .B(_373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_003_));
 sky130_fd_sc_hd__xnor2_1 _676_ (.A(_211_),
    .B(_214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_pos_imag[4] ));
 sky130_fd_sc_hd__nor2_1 _677_ (.A(_222_),
    .B(_223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\fft_inst.bfly_pos_real[4] ));
 sky130_fd_sc_hd__nand2_1 _678_ (.A(_224_),
    .B(_225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_1 _679_ (.A(_228_),
    .B(_229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _680_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _681_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _682_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _683_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _684_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _685_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _686_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _687_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _688_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _689_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _690_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _691_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _692_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _693_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _694_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _695_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _696_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _697_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _698_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _699_ (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _700_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _701_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _702_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _703_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _704_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _705_ (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _706_ (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _707_ (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _708_ (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _709_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _710_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _711_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _712_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _713_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _714_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _715_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _716_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _717_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _718_ (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _719_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _720_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _721_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _722_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _723_ (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _724_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _725_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _726_ (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _727_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _728_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _729_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _730_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _731_ (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _732_ (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _733_ (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _734_ (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _735_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _736_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _737_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _738_ (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _739_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _740_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _741_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _742_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _743_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _744_ (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _745_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _746_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _747_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _748_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _749_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _750_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _751_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _752_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _753_ (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _754_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _755_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _756_ (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _757_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _758_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _759_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _760_ (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _761_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _762_ (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _763_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _764_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _765_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _766_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_103_));
 sky130_fd_sc_hd__dfrtp_1 _767_ (.CLK(clknet_3_0__leaf_clk),
    .D(_104_),
    .RESET_B(_016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uo_out_delay_gen[1].uo_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _768_ (.CLK(clknet_3_2__leaf_clk),
    .D(_105_),
    .RESET_B(_017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uo_out_delay_gen[2].uo_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _769_ (.CLK(clknet_3_0__leaf_clk),
    .D(_106_),
    .RESET_B(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uo_out_delay_gen[3].uo_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _770_ (.CLK(clknet_3_0__leaf_clk),
    .D(_107_),
    .RESET_B(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uo_out_delay_gen[4].uo_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _771_ (.CLK(clknet_3_0__leaf_clk),
    .D(_108_),
    .RESET_B(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uo_out_delay_gen[5].uo_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _772_ (.CLK(clknet_3_0__leaf_clk),
    .D(_109_),
    .RESET_B(_021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uo_out_delay_gen[6].uo_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _773_ (.CLK(clknet_3_0__leaf_clk),
    .D(_110_),
    .RESET_B(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\disp_inst.output_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _774_ (.CLK(clknet_3_0__leaf_clk),
    .D(_111_),
    .RESET_B(_023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\disp_inst.output_counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _775_ (.CLK(clknet_3_0__leaf_clk),
    .D(_112_),
    .RESET_B(_024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _776_ (.CLK(clknet_3_0__leaf_clk),
    .D(_113_),
    .RESET_B(_025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[0].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _777_ (.CLK(clknet_3_2__leaf_clk),
    .D(_114_),
    .RESET_B(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[1].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _778_ (.CLK(clknet_3_3__leaf_clk),
    .D(net43),
    .RESET_B(_027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[2].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _779_ (.CLK(clknet_3_2__leaf_clk),
    .D(_116_),
    .RESET_B(_028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[3].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _780_ (.CLK(clknet_3_0__leaf_clk),
    .D(_117_),
    .RESET_B(_029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[4].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _781_ (.CLK(clknet_3_1__leaf_clk),
    .D(_118_),
    .RESET_B(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[5].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _782_ (.CLK(clknet_3_1__leaf_clk),
    .D(_119_),
    .RESET_B(_031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[6].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _783_ (.CLK(clknet_3_3__leaf_clk),
    .D(net65),
    .RESET_B(_032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\out_delay_gen[7].out_delay_inst.A ));
 sky130_fd_sc_hd__dfrtp_1 _784_ (.CLK(clknet_3_0__leaf_clk),
    .D(_121_),
    .RESET_B(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\disp_inst.processing ));
 sky130_fd_sc_hd__dfrtp_2 _785_ (.CLK(clknet_3_2__leaf_clk),
    .D(_122_),
    .RESET_B(_034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\disp_inst.done ));
 sky130_fd_sc_hd__dfrtp_1 _786_ (.CLK(clknet_3_2__leaf_clk),
    .D(_123_),
    .RESET_B(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(processing_dly));
 sky130_fd_sc_hd__dfstp_1 _787_ (.CLK(clknet_3_2__leaf_clk),
    .D(net30),
    .SET_B(\rst_delay.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(rst_sync1));
 sky130_fd_sc_hd__dfstp_1 _788_ (.CLK(clknet_3_2__leaf_clk),
    .D(net34),
    .SET_B(\rst_delay.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.rst ));
 sky130_fd_sc_hd__dfrtp_4 _789_ (.CLK(clknet_3_6__leaf_clk),
    .D(_124_),
    .RESET_B(_036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _790_ (.CLK(clknet_3_7__leaf_clk),
    .D(_125_),
    .RESET_B(_037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _791_ (.CLK(clknet_3_4__leaf_clk),
    .D(_126_),
    .RESET_B(_038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_real[4] ));
 sky130_fd_sc_hd__dfrtp_4 _792_ (.CLK(clknet_3_4__leaf_clk),
    .D(_127_),
    .RESET_B(_039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_real[5] ));
 sky130_fd_sc_hd__dfrtp_4 _793_ (.CLK(clknet_3_5__leaf_clk),
    .D(_128_),
    .RESET_B(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _794_ (.CLK(clknet_3_5__leaf_clk),
    .D(_129_),
    .RESET_B(_041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_real[7] ));
 sky130_fd_sc_hd__dfrtp_1 _795_ (.CLK(clknet_3_6__leaf_clk),
    .D(_130_),
    .RESET_B(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\io_inst.prev_in0 ));
 sky130_fd_sc_hd__dfrtp_4 _796_ (.CLK(clknet_3_6__leaf_clk),
    .D(_131_),
    .RESET_B(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_imag[4] ));
 sky130_fd_sc_hd__dfrtp_4 _797_ (.CLK(clknet_3_7__leaf_clk),
    .D(_132_),
    .RESET_B(_044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _798_ (.CLK(clknet_3_7__leaf_clk),
    .D(_133_),
    .RESET_B(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _799_ (.CLK(clknet_3_7__leaf_clk),
    .D(_134_),
    .RESET_B(_046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_imag[7] ));
 sky130_fd_sc_hd__dfrtp_4 _800_ (.CLK(clknet_3_4__leaf_clk),
    .D(_135_),
    .RESET_B(_047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_real[4] ));
 sky130_fd_sc_hd__dfrtp_4 _801_ (.CLK(clknet_3_5__leaf_clk),
    .D(_136_),
    .RESET_B(_048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _802_ (.CLK(clknet_3_5__leaf_clk),
    .D(_137_),
    .RESET_B(_049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _803_ (.CLK(clknet_3_5__leaf_clk),
    .D(_138_),
    .RESET_B(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_real[7] ));
 sky130_fd_sc_hd__dfrtp_4 _804_ (.CLK(clknet_3_4__leaf_clk),
    .D(_139_),
    .RESET_B(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_real[4] ));
 sky130_fd_sc_hd__dfrtp_4 _805_ (.CLK(clknet_3_5__leaf_clk),
    .D(_140_),
    .RESET_B(_052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _806_ (.CLK(clknet_3_4__leaf_clk),
    .D(_141_),
    .RESET_B(_053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _807_ (.CLK(clknet_3_5__leaf_clk),
    .D(_142_),
    .RESET_B(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.B_real[7] ));
 sky130_fd_sc_hd__dfrtp_4 _808_ (.CLK(clknet_3_7__leaf_clk),
    .D(_143_),
    .RESET_B(_055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_imag[4] ));
 sky130_fd_sc_hd__dfrtp_4 _809_ (.CLK(clknet_3_6__leaf_clk),
    .D(_144_),
    .RESET_B(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _810_ (.CLK(clknet_3_7__leaf_clk),
    .D(_145_),
    .RESET_B(_057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _811_ (.CLK(clknet_3_5__leaf_clk),
    .D(_146_),
    .RESET_B(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_imag[7] ));
 sky130_fd_sc_hd__dfrtp_1 _812_ (.CLK(clknet_3_4__leaf_clk),
    .D(_147_),
    .RESET_B(_059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_real[4] ));
 sky130_fd_sc_hd__dfrtp_4 _813_ (.CLK(clknet_3_4__leaf_clk),
    .D(_148_),
    .RESET_B(_060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _814_ (.CLK(clknet_3_5__leaf_clk),
    .D(_149_),
    .RESET_B(_061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _815_ (.CLK(clknet_3_5__leaf_clk),
    .D(_150_),
    .RESET_B(_062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.A_real[7] ));
 sky130_fd_sc_hd__dfrtp_1 _816_ (.CLK(clknet_3_2__leaf_clk),
    .D(_151_),
    .RESET_B(_063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\io_inst.prev_in1 ));
 sky130_fd_sc_hd__dfrtp_4 _817_ (.CLK(clknet_3_7__leaf_clk),
    .D(_152_),
    .RESET_B(_064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_imag[4] ));
 sky130_fd_sc_hd__dfrtp_4 _818_ (.CLK(clknet_3_7__leaf_clk),
    .D(_153_),
    .RESET_B(_065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _819_ (.CLK(clknet_3_6__leaf_clk),
    .D(_154_),
    .RESET_B(_066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _820_ (.CLK(clknet_3_5__leaf_clk),
    .D(_155_),
    .RESET_B(_067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_1.B_imag[7] ));
 sky130_fd_sc_hd__dfrtp_1 _821_ (.CLK(clknet_3_6__leaf_clk),
    .D(_156_),
    .RESET_B(_068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_imag[4] ));
 sky130_fd_sc_hd__dfrtp_4 _822_ (.CLK(clknet_3_6__leaf_clk),
    .D(_157_),
    .RESET_B(_069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_imag[5] ));
 sky130_fd_sc_hd__dfrtp_4 _823_ (.CLK(clknet_3_7__leaf_clk),
    .D(_158_),
    .RESET_B(_070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _824_ (.CLK(clknet_3_5__leaf_clk),
    .D(_159_),
    .RESET_B(_071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft_inst.bfly_stage1_0.A_imag[7] ));
 sky130_fd_sc_hd__dfrtp_1 _825_ (.CLK(clknet_3_2__leaf_clk),
    .D(\fft_inst.bfly_pos_imag[4] ),
    .RESET_B(_072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_imag[4] ));
 sky130_fd_sc_hd__dfrtp_1 _826_ (.CLK(clknet_3_2__leaf_clk),
    .D(\fft_inst.bfly_pos_imag[5] ),
    .RESET_B(_073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _827_ (.CLK(clknet_3_3__leaf_clk),
    .D(\fft_inst.bfly_pos_imag[6] ),
    .RESET_B(_074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _828_ (.CLK(clknet_3_3__leaf_clk),
    .D(\fft_inst.bfly_pos_imag[7] ),
    .RESET_B(_075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_imag[7] ));
 sky130_fd_sc_hd__dfrtp_1 _829_ (.CLK(clknet_3_0__leaf_clk),
    .D(_004_),
    .RESET_B(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_real[4] ));
 sky130_fd_sc_hd__dfrtp_1 _830_ (.CLK(clknet_3_1__leaf_clk),
    .D(_005_),
    .RESET_B(_077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _831_ (.CLK(clknet_3_1__leaf_clk),
    .D(_006_),
    .RESET_B(_078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _832_ (.CLK(clknet_3_1__leaf_clk),
    .D(_007_),
    .RESET_B(_079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_real[7] ));
 sky130_fd_sc_hd__dfrtp_1 _833_ (.CLK(clknet_3_0__leaf_clk),
    .D(\fft_inst.bfly_pos_real[4] ),
    .RESET_B(_080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_real[4] ));
 sky130_fd_sc_hd__dfrtp_1 _834_ (.CLK(clknet_3_1__leaf_clk),
    .D(\fft_inst.bfly_pos_real[5] ),
    .RESET_B(_081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _835_ (.CLK(clknet_3_1__leaf_clk),
    .D(\fft_inst.bfly_pos_real[6] ),
    .RESET_B(_082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _836_ (.CLK(clknet_3_1__leaf_clk),
    .D(\fft_inst.bfly_pos_real[7] ),
    .RESET_B(_083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft1_real[7] ));
 sky130_fd_sc_hd__dfrtp_1 _837_ (.CLK(clknet_3_0__leaf_clk),
    .D(\fft_inst.bfly_neg_real[4] ),
    .RESET_B(_084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_real[4] ));
 sky130_fd_sc_hd__dfrtp_1 _838_ (.CLK(clknet_3_1__leaf_clk),
    .D(\fft_inst.bfly_neg_real[5] ),
    .RESET_B(_085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _839_ (.CLK(clknet_3_1__leaf_clk),
    .D(\fft_inst.bfly_neg_real[6] ),
    .RESET_B(_086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _840_ (.CLK(clknet_3_4__leaf_clk),
    .D(\fft_inst.bfly_neg_real[7] ),
    .RESET_B(_087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_real[7] ));
 sky130_fd_sc_hd__dfrtp_1 _841_ (.CLK(clknet_3_2__leaf_clk),
    .D(_008_),
    .RESET_B(_088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_imag[4] ));
 sky130_fd_sc_hd__dfrtp_1 _842_ (.CLK(clknet_3_2__leaf_clk),
    .D(_009_),
    .RESET_B(_089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _843_ (.CLK(clknet_3_3__leaf_clk),
    .D(_010_),
    .RESET_B(_090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _844_ (.CLK(clknet_3_3__leaf_clk),
    .D(_011_),
    .RESET_B(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_imag[7] ));
 sky130_fd_sc_hd__dfrtp_1 _845_ (.CLK(clknet_3_2__leaf_clk),
    .D(_012_),
    .RESET_B(_092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_imag[4] ));
 sky130_fd_sc_hd__dfrtp_1 _846_ (.CLK(clknet_3_2__leaf_clk),
    .D(_013_),
    .RESET_B(_093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _847_ (.CLK(clknet_3_3__leaf_clk),
    .D(_014_),
    .RESET_B(_094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _848_ (.CLK(clknet_3_3__leaf_clk),
    .D(_015_),
    .RESET_B(_095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft2_imag[7] ));
 sky130_fd_sc_hd__dfrtp_1 _849_ (.CLK(clknet_3_0__leaf_clk),
    .D(_000_),
    .RESET_B(_096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_real[4] ));
 sky130_fd_sc_hd__dfrtp_1 _850_ (.CLK(clknet_3_0__leaf_clk),
    .D(_001_),
    .RESET_B(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_real[5] ));
 sky130_fd_sc_hd__dfrtp_1 _851_ (.CLK(clknet_3_1__leaf_clk),
    .D(_002_),
    .RESET_B(_098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_real[6] ));
 sky130_fd_sc_hd__dfrtp_1 _852_ (.CLK(clknet_3_1__leaf_clk),
    .D(_003_),
    .RESET_B(_099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft0_real[7] ));
 sky130_fd_sc_hd__dfrtp_1 _853_ (.CLK(clknet_3_2__leaf_clk),
    .D(\fft_inst.bfly_neg_imag[4] ),
    .RESET_B(_100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_imag[4] ));
 sky130_fd_sc_hd__dfrtp_1 _854_ (.CLK(clknet_3_3__leaf_clk),
    .D(\fft_inst.bfly_neg_imag[5] ),
    .RESET_B(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_imag[5] ));
 sky130_fd_sc_hd__dfrtp_1 _855_ (.CLK(clknet_3_3__leaf_clk),
    .D(\fft_inst.bfly_neg_imag[6] ),
    .RESET_B(_102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_imag[6] ));
 sky130_fd_sc_hd__dfrtp_1 _856_ (.CLK(clknet_3_3__leaf_clk),
    .D(\fft_inst.bfly_neg_imag[7] ),
    .RESET_B(_103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\fft3_imag[7] ));
 sky130_fd_sc_hd__conb_1 \uo_out_delay_gen[0].uo_delay_inst.buf1_31  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__conb_1 \uo_out_delay_gen[7].uo_delay_inst.buf1_32  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_2 _860_ (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__buf_2 _861_ (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__buf_2 _862_ (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__buf_2 _863_ (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[3]));
 sky130_fd_sc_hd__buf_2 _864_ (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[4]));
 sky130_fd_sc_hd__buf_2 _865_ (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[5]));
 sky130_fd_sc_hd__buf_2 _866_ (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__buf_2 _867_ (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__buf_2 _868_ (.A(\out_delay_gen[0].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__buf_2 _869_ (.A(\out_delay_gen[1].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _870_ (.A(\out_delay_gen[2].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__buf_2 _871_ (.A(\out_delay_gen[3].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__buf_2 _872_ (.A(\out_delay_gen[4].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__buf_2 _873_ (.A(\out_delay_gen[5].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__buf_2 _874_ (.A(\out_delay_gen[6].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__buf_2 _875_ (.A(\out_delay_gen[7].out_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__buf_2 _876_ (.A(\uo_out_delay_gen[0].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _877_ (.A(\uo_out_delay_gen[1].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _878_ (.A(\uo_out_delay_gen[2].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__buf_2 _879_ (.A(\uo_out_delay_gen[3].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _880_ (.A(\uo_out_delay_gen[4].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__buf_2 _881_ (.A(\uo_out_delay_gen[5].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _882_ (.A(\uo_out_delay_gen[6].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _883_ (.A(\uo_out_delay_gen[7].uo_delay_inst.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf1  (.A(\out_delay_gen[0].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf10  (.A(\out_delay_gen[0].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf11  (.A(\out_delay_gen[0].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf12  (.A(\out_delay_gen[0].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf13  (.A(\out_delay_gen[0].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf14  (.A(\out_delay_gen[0].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf15  (.A(\out_delay_gen[0].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf16  (.A(\out_delay_gen[0].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf17  (.A(\out_delay_gen[0].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf18  (.A(\out_delay_gen[0].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf19  (.A(\out_delay_gen[0].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf2  (.A(\out_delay_gen[0].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf20  (.A(\out_delay_gen[0].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf21  (.A(\out_delay_gen[0].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf22  (.A(\out_delay_gen[0].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf23  (.A(\out_delay_gen[0].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf24  (.A(\out_delay_gen[0].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf25  (.A(\out_delay_gen[0].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf26  (.A(\out_delay_gen[0].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf27  (.A(\out_delay_gen[0].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf28  (.A(\out_delay_gen[0].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf29  (.A(\out_delay_gen[0].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf3  (.A(\out_delay_gen[0].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf30  (.A(\out_delay_gen[0].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf31  (.A(\out_delay_gen[0].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf32  (.A(\out_delay_gen[0].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf33  (.A(\out_delay_gen[0].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf34  (.A(\out_delay_gen[0].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf35  (.A(\out_delay_gen[0].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf36  (.A(\out_delay_gen[0].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf37  (.A(\out_delay_gen[0].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf38  (.A(\out_delay_gen[0].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf39  (.A(\out_delay_gen[0].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf4  (.A(\out_delay_gen[0].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf40  (.A(\out_delay_gen[0].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf5  (.A(\out_delay_gen[0].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf6  (.A(\out_delay_gen[0].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf7  (.A(\out_delay_gen[0].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf8  (.A(\out_delay_gen[0].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[0].out_delay_inst.buf9  (.A(\out_delay_gen[0].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[0].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf1  (.A(\out_delay_gen[1].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf10  (.A(\out_delay_gen[1].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf11  (.A(\out_delay_gen[1].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf12  (.A(\out_delay_gen[1].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf13  (.A(\out_delay_gen[1].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf14  (.A(\out_delay_gen[1].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf15  (.A(\out_delay_gen[1].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf16  (.A(\out_delay_gen[1].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf17  (.A(\out_delay_gen[1].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf18  (.A(\out_delay_gen[1].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf19  (.A(\out_delay_gen[1].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf2  (.A(\out_delay_gen[1].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf20  (.A(\out_delay_gen[1].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf21  (.A(\out_delay_gen[1].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf22  (.A(\out_delay_gen[1].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf23  (.A(\out_delay_gen[1].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf24  (.A(\out_delay_gen[1].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf25  (.A(\out_delay_gen[1].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf26  (.A(\out_delay_gen[1].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf27  (.A(\out_delay_gen[1].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf28  (.A(\out_delay_gen[1].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf29  (.A(\out_delay_gen[1].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf3  (.A(\out_delay_gen[1].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf30  (.A(\out_delay_gen[1].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf31  (.A(\out_delay_gen[1].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf32  (.A(\out_delay_gen[1].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf33  (.A(\out_delay_gen[1].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf34  (.A(\out_delay_gen[1].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf35  (.A(\out_delay_gen[1].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf36  (.A(\out_delay_gen[1].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf37  (.A(\out_delay_gen[1].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf38  (.A(\out_delay_gen[1].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf39  (.A(\out_delay_gen[1].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf4  (.A(\out_delay_gen[1].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf40  (.A(\out_delay_gen[1].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf5  (.A(\out_delay_gen[1].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf6  (.A(\out_delay_gen[1].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf7  (.A(\out_delay_gen[1].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf8  (.A(\out_delay_gen[1].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[1].out_delay_inst.buf9  (.A(\out_delay_gen[1].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[1].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf1  (.A(\out_delay_gen[2].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf10  (.A(\out_delay_gen[2].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf11  (.A(\out_delay_gen[2].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf12  (.A(\out_delay_gen[2].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf13  (.A(\out_delay_gen[2].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf14  (.A(\out_delay_gen[2].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf15  (.A(\out_delay_gen[2].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf16  (.A(\out_delay_gen[2].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf17  (.A(\out_delay_gen[2].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf18  (.A(\out_delay_gen[2].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf19  (.A(\out_delay_gen[2].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf2  (.A(\out_delay_gen[2].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf20  (.A(\out_delay_gen[2].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf21  (.A(\out_delay_gen[2].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf22  (.A(\out_delay_gen[2].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf23  (.A(\out_delay_gen[2].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf24  (.A(\out_delay_gen[2].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf25  (.A(\out_delay_gen[2].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf26  (.A(\out_delay_gen[2].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf27  (.A(\out_delay_gen[2].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf28  (.A(\out_delay_gen[2].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf29  (.A(\out_delay_gen[2].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf3  (.A(\out_delay_gen[2].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf30  (.A(\out_delay_gen[2].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf31  (.A(\out_delay_gen[2].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf32  (.A(\out_delay_gen[2].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf33  (.A(\out_delay_gen[2].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf34  (.A(\out_delay_gen[2].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf35  (.A(\out_delay_gen[2].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf36  (.A(\out_delay_gen[2].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf37  (.A(\out_delay_gen[2].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf38  (.A(\out_delay_gen[2].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf39  (.A(\out_delay_gen[2].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf4  (.A(\out_delay_gen[2].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf40  (.A(\out_delay_gen[2].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.X ));
 sky130_fd_sc_hd__buf_1 \out_delay_gen[2].out_delay_inst.buf5  (.A(\out_delay_gen[2].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf6  (.A(\out_delay_gen[2].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf7  (.A(\out_delay_gen[2].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf8  (.A(\out_delay_gen[2].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[2].out_delay_inst.buf9  (.A(\out_delay_gen[2].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[2].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf1  (.A(\out_delay_gen[3].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf10  (.A(\out_delay_gen[3].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf11  (.A(\out_delay_gen[3].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf12  (.A(\out_delay_gen[3].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf13  (.A(\out_delay_gen[3].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf14  (.A(\out_delay_gen[3].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf15  (.A(\out_delay_gen[3].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf16  (.A(\out_delay_gen[3].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf17  (.A(\out_delay_gen[3].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf18  (.A(\out_delay_gen[3].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf19  (.A(\out_delay_gen[3].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf2  (.A(\out_delay_gen[3].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf20  (.A(\out_delay_gen[3].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf21  (.A(\out_delay_gen[3].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf22  (.A(\out_delay_gen[3].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf23  (.A(\out_delay_gen[3].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf24  (.A(\out_delay_gen[3].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf25  (.A(\out_delay_gen[3].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf26  (.A(\out_delay_gen[3].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf27  (.A(\out_delay_gen[3].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf28  (.A(\out_delay_gen[3].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf29  (.A(\out_delay_gen[3].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf3  (.A(\out_delay_gen[3].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf30  (.A(\out_delay_gen[3].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf31  (.A(\out_delay_gen[3].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf32  (.A(\out_delay_gen[3].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf33  (.A(\out_delay_gen[3].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf34  (.A(\out_delay_gen[3].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf35  (.A(\out_delay_gen[3].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf36  (.A(\out_delay_gen[3].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf37  (.A(\out_delay_gen[3].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf38  (.A(\out_delay_gen[3].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf39  (.A(\out_delay_gen[3].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf4  (.A(\out_delay_gen[3].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf40  (.A(\out_delay_gen[3].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf5  (.A(\out_delay_gen[3].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf6  (.A(\out_delay_gen[3].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w6 ));
 sky130_fd_sc_hd__buf_1 \out_delay_gen[3].out_delay_inst.buf7  (.A(\out_delay_gen[3].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf8  (.A(\out_delay_gen[3].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[3].out_delay_inst.buf9  (.A(\out_delay_gen[3].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[3].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf1  (.A(\out_delay_gen[4].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf10  (.A(\out_delay_gen[4].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf11  (.A(\out_delay_gen[4].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf12  (.A(\out_delay_gen[4].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf13  (.A(\out_delay_gen[4].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf14  (.A(\out_delay_gen[4].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf15  (.A(\out_delay_gen[4].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf16  (.A(\out_delay_gen[4].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf17  (.A(\out_delay_gen[4].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf18  (.A(\out_delay_gen[4].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf19  (.A(\out_delay_gen[4].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf2  (.A(\out_delay_gen[4].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf20  (.A(\out_delay_gen[4].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf21  (.A(\out_delay_gen[4].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf22  (.A(\out_delay_gen[4].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf23  (.A(\out_delay_gen[4].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf24  (.A(\out_delay_gen[4].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf25  (.A(\out_delay_gen[4].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf26  (.A(\out_delay_gen[4].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf27  (.A(\out_delay_gen[4].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf28  (.A(\out_delay_gen[4].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf29  (.A(\out_delay_gen[4].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf3  (.A(\out_delay_gen[4].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf30  (.A(\out_delay_gen[4].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf31  (.A(\out_delay_gen[4].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf32  (.A(\out_delay_gen[4].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf33  (.A(\out_delay_gen[4].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf34  (.A(\out_delay_gen[4].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf35  (.A(\out_delay_gen[4].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf36  (.A(\out_delay_gen[4].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf37  (.A(\out_delay_gen[4].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf38  (.A(\out_delay_gen[4].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf39  (.A(\out_delay_gen[4].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf4  (.A(\out_delay_gen[4].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf40  (.A(\out_delay_gen[4].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf5  (.A(\out_delay_gen[4].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf6  (.A(\out_delay_gen[4].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf7  (.A(\out_delay_gen[4].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf8  (.A(\out_delay_gen[4].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[4].out_delay_inst.buf9  (.A(\out_delay_gen[4].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[4].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf1  (.A(\out_delay_gen[5].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf10  (.A(\out_delay_gen[5].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf11  (.A(\out_delay_gen[5].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf12  (.A(\out_delay_gen[5].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf13  (.A(\out_delay_gen[5].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf14  (.A(\out_delay_gen[5].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf15  (.A(\out_delay_gen[5].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf16  (.A(\out_delay_gen[5].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf17  (.A(\out_delay_gen[5].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf18  (.A(\out_delay_gen[5].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf19  (.A(\out_delay_gen[5].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf2  (.A(\out_delay_gen[5].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf20  (.A(\out_delay_gen[5].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf21  (.A(\out_delay_gen[5].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf22  (.A(\out_delay_gen[5].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf23  (.A(\out_delay_gen[5].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf24  (.A(\out_delay_gen[5].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf25  (.A(\out_delay_gen[5].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf26  (.A(\out_delay_gen[5].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf27  (.A(\out_delay_gen[5].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf28  (.A(\out_delay_gen[5].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf29  (.A(\out_delay_gen[5].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf3  (.A(\out_delay_gen[5].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf30  (.A(\out_delay_gen[5].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf31  (.A(\out_delay_gen[5].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf32  (.A(\out_delay_gen[5].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf33  (.A(\out_delay_gen[5].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf34  (.A(\out_delay_gen[5].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf35  (.A(\out_delay_gen[5].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf36  (.A(\out_delay_gen[5].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf37  (.A(\out_delay_gen[5].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf38  (.A(\out_delay_gen[5].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf39  (.A(\out_delay_gen[5].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf4  (.A(\out_delay_gen[5].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf40  (.A(\out_delay_gen[5].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf5  (.A(\out_delay_gen[5].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf6  (.A(\out_delay_gen[5].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf7  (.A(\out_delay_gen[5].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf8  (.A(\out_delay_gen[5].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[5].out_delay_inst.buf9  (.A(\out_delay_gen[5].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[5].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf1  (.A(\out_delay_gen[6].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf10  (.A(\out_delay_gen[6].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf11  (.A(\out_delay_gen[6].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf12  (.A(\out_delay_gen[6].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf13  (.A(\out_delay_gen[6].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf14  (.A(\out_delay_gen[6].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf15  (.A(\out_delay_gen[6].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf16  (.A(\out_delay_gen[6].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf17  (.A(\out_delay_gen[6].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf18  (.A(\out_delay_gen[6].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf19  (.A(\out_delay_gen[6].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf2  (.A(\out_delay_gen[6].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf20  (.A(\out_delay_gen[6].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf21  (.A(\out_delay_gen[6].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf22  (.A(\out_delay_gen[6].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf23  (.A(\out_delay_gen[6].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf24  (.A(\out_delay_gen[6].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf25  (.A(\out_delay_gen[6].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf26  (.A(\out_delay_gen[6].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf27  (.A(\out_delay_gen[6].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf28  (.A(\out_delay_gen[6].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf29  (.A(\out_delay_gen[6].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf3  (.A(\out_delay_gen[6].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf30  (.A(\out_delay_gen[6].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf31  (.A(\out_delay_gen[6].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf32  (.A(\out_delay_gen[6].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf33  (.A(\out_delay_gen[6].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf34  (.A(\out_delay_gen[6].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf35  (.A(\out_delay_gen[6].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf36  (.A(\out_delay_gen[6].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf37  (.A(\out_delay_gen[6].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf38  (.A(\out_delay_gen[6].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf39  (.A(\out_delay_gen[6].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf4  (.A(\out_delay_gen[6].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf40  (.A(\out_delay_gen[6].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf5  (.A(\out_delay_gen[6].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf6  (.A(\out_delay_gen[6].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf7  (.A(\out_delay_gen[6].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf8  (.A(\out_delay_gen[6].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[6].out_delay_inst.buf9  (.A(\out_delay_gen[6].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[6].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf1  (.A(\out_delay_gen[7].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf10  (.A(\out_delay_gen[7].out_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf11  (.A(\out_delay_gen[7].out_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf12  (.A(\out_delay_gen[7].out_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf13  (.A(\out_delay_gen[7].out_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf14  (.A(\out_delay_gen[7].out_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf15  (.A(\out_delay_gen[7].out_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf16  (.A(\out_delay_gen[7].out_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf17  (.A(\out_delay_gen[7].out_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf18  (.A(\out_delay_gen[7].out_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf19  (.A(\out_delay_gen[7].out_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf2  (.A(\out_delay_gen[7].out_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf20  (.A(\out_delay_gen[7].out_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf21  (.A(\out_delay_gen[7].out_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf22  (.A(\out_delay_gen[7].out_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf23  (.A(\out_delay_gen[7].out_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf24  (.A(\out_delay_gen[7].out_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf25  (.A(\out_delay_gen[7].out_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf26  (.A(\out_delay_gen[7].out_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf27  (.A(\out_delay_gen[7].out_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf28  (.A(\out_delay_gen[7].out_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf29  (.A(\out_delay_gen[7].out_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf3  (.A(\out_delay_gen[7].out_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf30  (.A(\out_delay_gen[7].out_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf31  (.A(\out_delay_gen[7].out_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf32  (.A(\out_delay_gen[7].out_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf33  (.A(\out_delay_gen[7].out_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf34  (.A(\out_delay_gen[7].out_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf35  (.A(\out_delay_gen[7].out_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf36  (.A(\out_delay_gen[7].out_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf37  (.A(\out_delay_gen[7].out_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf38  (.A(\out_delay_gen[7].out_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf39  (.A(\out_delay_gen[7].out_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf4  (.A(\out_delay_gen[7].out_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf40  (.A(\out_delay_gen[7].out_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf5  (.A(\out_delay_gen[7].out_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf6  (.A(\out_delay_gen[7].out_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf7  (.A(\out_delay_gen[7].out_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf8  (.A(\out_delay_gen[7].out_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \out_delay_gen[7].out_delay_inst.buf9  (.A(\out_delay_gen[7].out_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\out_delay_gen[7].out_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf1  (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf10  (.A(\rst_delay.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf11  (.A(\rst_delay.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf12  (.A(\rst_delay.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf13  (.A(\rst_delay.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf14  (.A(\rst_delay.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf15  (.A(\rst_delay.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf16  (.A(\rst_delay.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf17  (.A(\rst_delay.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf18  (.A(\rst_delay.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf19  (.A(\rst_delay.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf2  (.A(\rst_delay.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf20  (.A(\rst_delay.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf21  (.A(\rst_delay.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf22  (.A(\rst_delay.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf23  (.A(\rst_delay.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf24  (.A(\rst_delay.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf25  (.A(\rst_delay.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf26  (.A(\rst_delay.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf27  (.A(\rst_delay.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf28  (.A(\rst_delay.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf29  (.A(\rst_delay.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf3  (.A(\rst_delay.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf30  (.A(\rst_delay.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf31  (.A(\rst_delay.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf32  (.A(\rst_delay.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf33  (.A(\rst_delay.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf34  (.A(\rst_delay.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf35  (.A(\rst_delay.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf36  (.A(\rst_delay.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf37  (.A(\rst_delay.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf38  (.A(\rst_delay.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf39  (.A(\rst_delay.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf4  (.A(\rst_delay.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w4 ));
 sky130_fd_sc_hd__buf_1 \rst_delay.buf40  (.A(\rst_delay.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.X ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf5  (.A(\rst_delay.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf6  (.A(\rst_delay.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w6 ));
 sky130_fd_sc_hd__buf_1 \rst_delay.buf7  (.A(\rst_delay.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf8  (.A(\rst_delay.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \rst_delay.buf9  (.A(\rst_delay.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\rst_delay.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[0].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[0].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[1].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[1].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[1].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[2].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[2].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[2].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[3].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[3].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[3].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[4].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[4].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[4].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[5].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[5].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[5].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[6].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[6].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[6].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf1  (.A(\uio_oe_delay_gen[0].uio_oe_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf10  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf11  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf12  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf13  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf14  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf15  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf16  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf17  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf18  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf19  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf2  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf20  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf21  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf22  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf23  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf24  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf25  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf26  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf27  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf28  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf29  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf3  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf30  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf31  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf32  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf33  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf34  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf35  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf36  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf37  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf38  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf39  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf4  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf40  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf5  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf6  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf7  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf8  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uio_oe_delay_gen[7].uio_oe_delay_inst.buf9  (.A(\uio_oe_delay_gen[7].uio_oe_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uio_oe_delay_gen[7].uio_oe_delay_inst.w9 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf1  (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[0].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[0].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[0].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[0].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[0].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[0].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[0].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[0].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[0].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[0].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[0].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[0].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[0].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[0].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[0].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[0].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[0].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[0].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[0].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[0].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[0].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[0].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[0].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[0].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[0].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[0].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[0].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[0].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[0].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[0].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[0].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[0].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[0].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[0].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.X ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[0].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[0].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[0].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[0].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[0].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[0].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[0].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf1  (.A(\uo_out_delay_gen[1].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[1].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[1].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[1].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[1].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[1].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[1].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[1].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[1].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[1].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[1].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[1].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[1].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[1].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[1].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[1].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[1].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[1].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[1].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[1].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[1].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[1].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[1].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[1].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[1].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[1].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[1].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[1].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[1].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[1].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[1].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[1].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[1].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[1].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[1].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[1].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[1].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[1].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[1].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[1].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[1].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[1].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf1  (.A(\uo_out_delay_gen[2].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[2].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[2].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[2].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[2].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[2].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[2].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[2].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[2].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[2].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[2].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[2].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[2].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[2].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[2].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[2].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[2].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[2].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[2].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[2].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[2].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[2].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[2].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[2].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[2].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[2].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[2].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[2].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[2].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[2].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[2].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[2].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[2].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[2].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[2].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[2].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[2].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[2].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[2].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[2].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[2].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[2].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf1  (.A(\uo_out_delay_gen[3].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[3].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[3].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[3].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[3].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[3].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[3].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[3].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[3].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[3].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[3].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[3].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[3].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[3].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[3].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[3].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[3].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[3].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[3].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[3].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[3].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[3].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[3].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[3].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[3].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[3].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[3].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[3].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[3].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[3].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[3].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[3].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[3].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[3].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[3].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[3].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[3].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[3].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[3].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[3].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[3].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[3].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf1  (.A(\uo_out_delay_gen[4].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[4].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[4].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[4].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[4].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[4].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[4].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[4].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[4].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[4].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[4].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[4].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[4].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[4].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[4].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[4].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[4].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[4].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[4].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[4].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[4].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[4].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[4].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[4].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[4].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[4].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[4].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[4].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[4].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[4].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[4].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[4].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[4].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[4].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[4].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[4].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[4].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[4].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[4].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[4].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[4].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[4].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf1  (.A(\uo_out_delay_gen[5].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[5].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[5].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[5].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[5].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[5].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[5].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[5].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[5].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[5].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[5].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[5].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[5].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[5].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[5].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[5].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[5].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[5].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[5].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[5].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[5].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[5].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[5].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[5].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[5].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[5].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[5].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[5].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[5].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[5].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[5].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[5].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[5].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[5].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[5].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[5].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[5].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[5].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[5].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[5].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[5].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[5].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf1  (.A(\uo_out_delay_gen[6].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[6].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[6].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[6].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[6].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[6].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[6].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[6].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[6].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[6].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[6].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[6].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[6].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[6].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[6].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[6].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[6].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[6].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[6].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[6].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[6].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[6].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[6].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[6].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[6].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[6].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[6].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[6].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[6].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[6].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[6].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[6].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[6].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[6].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[6].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.X ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[6].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[6].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[6].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[6].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__clkbuf_1 \uo_out_delay_gen[6].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[6].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[6].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf1  (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w1 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf10  (.A(\uo_out_delay_gen[7].uo_delay_inst.w9 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w10 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf11  (.A(\uo_out_delay_gen[7].uo_delay_inst.w10 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w11 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf12  (.A(\uo_out_delay_gen[7].uo_delay_inst.w11 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w12 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf13  (.A(\uo_out_delay_gen[7].uo_delay_inst.w12 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w13 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf14  (.A(\uo_out_delay_gen[7].uo_delay_inst.w13 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w14 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf15  (.A(\uo_out_delay_gen[7].uo_delay_inst.w14 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w15 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf16  (.A(\uo_out_delay_gen[7].uo_delay_inst.w15 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w16 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf17  (.A(\uo_out_delay_gen[7].uo_delay_inst.w16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w17 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf18  (.A(\uo_out_delay_gen[7].uo_delay_inst.w17 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w18 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf19  (.A(\uo_out_delay_gen[7].uo_delay_inst.w18 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w19 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf2  (.A(\uo_out_delay_gen[7].uo_delay_inst.w1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w2 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf20  (.A(\uo_out_delay_gen[7].uo_delay_inst.w19 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w20 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf21  (.A(\uo_out_delay_gen[7].uo_delay_inst.w20 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w21 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf22  (.A(\uo_out_delay_gen[7].uo_delay_inst.w21 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w22 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf23  (.A(\uo_out_delay_gen[7].uo_delay_inst.w22 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w23 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf24  (.A(\uo_out_delay_gen[7].uo_delay_inst.w23 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w24 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf25  (.A(\uo_out_delay_gen[7].uo_delay_inst.w24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w25 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf26  (.A(\uo_out_delay_gen[7].uo_delay_inst.w25 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w26 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf27  (.A(\uo_out_delay_gen[7].uo_delay_inst.w26 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w27 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf28  (.A(\uo_out_delay_gen[7].uo_delay_inst.w27 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w28 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf29  (.A(\uo_out_delay_gen[7].uo_delay_inst.w28 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w29 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf3  (.A(\uo_out_delay_gen[7].uo_delay_inst.w2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w3 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf30  (.A(\uo_out_delay_gen[7].uo_delay_inst.w29 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w30 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf31  (.A(\uo_out_delay_gen[7].uo_delay_inst.w30 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w31 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf32  (.A(\uo_out_delay_gen[7].uo_delay_inst.w31 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w32 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf33  (.A(\uo_out_delay_gen[7].uo_delay_inst.w32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w33 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf34  (.A(\uo_out_delay_gen[7].uo_delay_inst.w33 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w34 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf35  (.A(\uo_out_delay_gen[7].uo_delay_inst.w34 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w35 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf36  (.A(\uo_out_delay_gen[7].uo_delay_inst.w35 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w36 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf37  (.A(\uo_out_delay_gen[7].uo_delay_inst.w36 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w37 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf38  (.A(\uo_out_delay_gen[7].uo_delay_inst.w37 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w38 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf39  (.A(\uo_out_delay_gen[7].uo_delay_inst.w38 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w39 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf4  (.A(\uo_out_delay_gen[7].uo_delay_inst.w3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w4 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf40  (.A(\uo_out_delay_gen[7].uo_delay_inst.w39 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.X ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf5  (.A(\uo_out_delay_gen[7].uo_delay_inst.w4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w5 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf6  (.A(\uo_out_delay_gen[7].uo_delay_inst.w5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w6 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf7  (.A(\uo_out_delay_gen[7].uo_delay_inst.w6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w7 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf8  (.A(\uo_out_delay_gen[7].uo_delay_inst.w7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w8 ));
 sky130_fd_sc_hd__buf_4 \uo_out_delay_gen[7].uo_delay_inst.buf9  (.A(\uo_out_delay_gen[7].uo_delay_inst.w8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\uo_out_delay_gen[7].uo_delay_inst.w9 ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(uio_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(uio_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(uio_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(uio_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(uio_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(uio_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(uio_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_4 fanout12 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_4 fanout14 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_4 fanout16 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout21 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 fanout23 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(\disp_inst.output_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(\disp_inst.output_counter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(\disp_inst.output_counter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(_161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout29 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__conb_1 _787__30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_8 clkload5 (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\fft_inst.rst ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_sync1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\uo_out_delay_gen[4].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\io_inst.prev_in0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\out_delay_gen[3].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\uo_out_delay_gen[1].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\uo_out_delay_gen[6].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(processing_dly),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\uo_out_delay_gen[3].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\out_delay_gen[2].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\uo_out_delay_gen[2].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\disp_inst.processing ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\uo_out_delay_gen[5].uo_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\io_inst.prev_in1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\fft_inst.bfly_stage1_0.B_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\fft_inst.bfly_stage1_0.B_imag[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\fft_inst.bfly_stage1_0.B_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\fft_inst.bfly_stage1_1.A_imag[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\fft_inst.bfly_stage1_1.A_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\fft_inst.bfly_stage1_1.B_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\out_delay_gen[4].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\out_delay_gen[1].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\fft_inst.bfly_stage1_1.B_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\fft_inst.bfly_stage1_1.B_imag[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\fft_inst.bfly_stage1_0.B_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\fft_inst.bfly_stage1_0.A_imag[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\fft_inst.bfly_stage1_0.A_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\fft_inst.bfly_stage1_1.B_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\out_delay_gen[0].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\out_delay_gen[5].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\fft0_real[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\fft_inst.bfly_stage1_1.A_real[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\out_delay_gen[6].out_delay_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\fft_inst.bfly_stage1_1.A_imag[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\fft_inst.bfly_stage1_0.A_imag[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\fft_inst.bfly_stage1_0.A_real[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_207 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_100 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_304 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_70 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_103 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_2_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_226 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_5_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_82 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_8 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_157 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_9_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_11_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_46 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_12_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_13_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_13_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_13_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_16 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_14_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_15_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_50 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_16_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_163 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_16_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_73 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_17_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_17_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_19_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_230 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_19_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_279 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_17 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_23_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_23_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_142 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_23_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_23_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_25_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_25_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_58 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_26_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_108 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_28_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_77 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_29_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_56 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_30_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_40 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_61 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_32_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_45 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_32 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_35_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_35_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_13 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_92 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_36_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_16 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_37_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_100 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
