VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_emmersonv_tiq_adc
  CLASS BLOCK ;
  FOREIGN tt_um_emmersonv_tiq_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 36.968998 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 195.889191 ;
    ANTENNADIFFAREA 109.297394 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    USE POWER ;
    ANTENNAGATEAREA 123.837997 ;
    ANTENNADIFFAREA 144.727646 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 92.190 35.065 124.310 36.670 ;
        RECT 128.520 35.780 132.230 38.540 ;
      LAYER pwell ;
        RECT 128.570 34.890 129.560 35.570 ;
        RECT 129.880 34.890 130.870 35.570 ;
        RECT 131.190 34.890 132.180 35.570 ;
        RECT 92.385 33.865 93.755 34.675 ;
        RECT 93.765 33.865 99.275 34.675 ;
        RECT 99.285 33.865 104.795 34.675 ;
        RECT 105.275 33.950 105.705 34.735 ;
        RECT 105.725 33.865 111.235 34.675 ;
        RECT 111.245 33.865 116.755 34.675 ;
        RECT 116.765 33.865 118.135 34.675 ;
        RECT 118.155 33.950 118.585 34.735 ;
        RECT 118.605 33.865 119.975 34.675 ;
        RECT 119.985 33.865 121.355 34.645 ;
        RECT 121.365 33.865 122.735 34.645 ;
        RECT 122.745 33.865 124.115 34.675 ;
        RECT 92.525 33.655 92.695 33.865 ;
        RECT 93.905 33.655 94.075 33.865 ;
        RECT 99.425 33.655 99.595 33.865 ;
        RECT 104.945 33.815 105.115 33.845 ;
        RECT 104.940 33.705 105.115 33.815 ;
        RECT 104.945 33.655 105.115 33.705 ;
        RECT 105.865 33.675 106.035 33.865 ;
        RECT 110.465 33.655 110.635 33.845 ;
        RECT 111.385 33.675 111.555 33.865 ;
        RECT 115.985 33.655 116.155 33.845 ;
        RECT 116.905 33.675 117.075 33.865 ;
        RECT 117.820 33.705 117.940 33.815 ;
        RECT 118.745 33.655 118.915 33.865 ;
        RECT 121.035 33.675 121.205 33.865 ;
        RECT 122.415 33.675 122.585 33.865 ;
        RECT 123.805 33.655 123.975 33.865 ;
        RECT 92.385 32.845 93.755 33.655 ;
        RECT 93.765 32.845 99.275 33.655 ;
        RECT 99.285 32.845 104.795 33.655 ;
        RECT 104.805 32.845 110.315 33.655 ;
        RECT 110.325 32.845 115.835 33.655 ;
        RECT 115.845 32.845 117.675 33.655 ;
        RECT 118.155 32.785 118.585 33.570 ;
        RECT 118.605 32.845 122.275 33.655 ;
        RECT 122.745 32.845 124.115 33.655 ;
        RECT 128.390 33.620 132.580 34.880 ;
      LAYER nwell ;
        RECT 92.190 29.625 124.310 32.455 ;
        RECT 128.520 30.860 132.230 33.620 ;
      LAYER pwell ;
        RECT 128.570 29.970 129.560 30.650 ;
        RECT 129.880 29.970 130.870 30.650 ;
        RECT 131.190 29.970 132.180 30.650 ;
        RECT 92.385 28.425 93.755 29.235 ;
        RECT 93.765 28.425 99.275 29.235 ;
        RECT 99.285 28.425 104.795 29.235 ;
        RECT 105.275 28.510 105.705 29.295 ;
        RECT 105.725 28.425 111.235 29.235 ;
        RECT 111.245 28.425 116.755 29.235 ;
        RECT 116.765 28.425 120.435 29.235 ;
        RECT 121.365 28.425 122.735 29.205 ;
        RECT 122.745 28.425 124.115 29.235 ;
        RECT 128.390 28.700 132.580 29.960 ;
        RECT 92.525 28.215 92.695 28.425 ;
        RECT 93.905 28.215 94.075 28.425 ;
        RECT 99.425 28.215 99.595 28.425 ;
        RECT 104.945 28.375 105.115 28.405 ;
        RECT 104.940 28.265 105.115 28.375 ;
        RECT 104.945 28.215 105.115 28.265 ;
        RECT 105.865 28.235 106.035 28.425 ;
        RECT 110.465 28.215 110.635 28.405 ;
        RECT 111.385 28.235 111.555 28.425 ;
        RECT 115.985 28.215 116.155 28.405 ;
        RECT 116.905 28.235 117.075 28.425 ;
        RECT 118.745 28.215 118.915 28.405 ;
        RECT 120.595 28.270 120.755 28.380 ;
        RECT 121.510 28.215 121.680 28.405 ;
        RECT 122.425 28.235 122.595 28.425 ;
        RECT 123.805 28.215 123.975 28.425 ;
        RECT 92.385 27.405 93.755 28.215 ;
        RECT 93.765 27.405 99.275 28.215 ;
        RECT 99.285 27.405 104.795 28.215 ;
        RECT 104.805 27.405 110.315 28.215 ;
        RECT 110.325 27.405 115.835 28.215 ;
        RECT 115.845 27.535 118.135 28.215 ;
        RECT 117.215 27.305 118.135 27.535 ;
        RECT 118.155 27.345 118.585 28.130 ;
        RECT 118.615 27.305 121.345 28.215 ;
        RECT 121.365 27.305 122.715 28.215 ;
        RECT 122.745 27.405 124.115 28.215 ;
      LAYER nwell ;
        RECT 92.190 24.185 124.310 27.015 ;
        RECT 128.520 25.930 132.230 28.690 ;
      LAYER pwell ;
        RECT 128.570 25.040 129.560 25.720 ;
        RECT 129.880 25.040 130.870 25.720 ;
        RECT 131.190 25.040 132.180 25.720 ;
        RECT 128.390 24.960 132.580 25.030 ;
        RECT 92.385 22.985 93.755 23.795 ;
        RECT 93.765 22.985 99.275 23.795 ;
        RECT 99.285 22.985 104.795 23.795 ;
        RECT 105.275 23.070 105.705 23.855 ;
        RECT 105.725 22.985 111.235 23.795 ;
        RECT 111.245 22.985 113.995 23.795 ;
        RECT 114.705 22.985 120.895 23.895 ;
        RECT 128.380 23.850 132.590 24.960 ;
        RECT 121.365 22.985 122.735 23.765 ;
        RECT 122.745 22.985 124.115 23.795 ;
        RECT 128.390 23.770 132.580 23.850 ;
        RECT 92.525 22.775 92.695 22.985 ;
        RECT 93.905 22.775 94.075 22.985 ;
        RECT 99.425 22.775 99.595 22.985 ;
        RECT 104.945 22.935 105.115 22.965 ;
        RECT 104.940 22.825 105.115 22.935 ;
        RECT 104.945 22.775 105.115 22.825 ;
        RECT 105.865 22.795 106.035 22.985 ;
        RECT 110.465 22.775 110.635 22.965 ;
        RECT 111.385 22.795 111.555 22.985 ;
        RECT 113.220 22.825 113.340 22.935 ;
        RECT 113.690 22.795 113.860 22.965 ;
        RECT 114.140 22.825 114.260 22.935 ;
        RECT 113.715 22.775 113.860 22.795 ;
        RECT 116.905 22.775 117.075 22.965 ;
        RECT 118.740 22.825 118.860 22.935 ;
        RECT 120.580 22.795 120.750 22.985 ;
        RECT 121.040 22.825 121.160 22.935 ;
        RECT 121.965 22.775 122.135 22.965 ;
        RECT 122.425 22.935 122.595 22.985 ;
        RECT 122.420 22.825 122.595 22.935 ;
        RECT 122.425 22.795 122.595 22.825 ;
        RECT 123.805 22.775 123.975 22.985 ;
        RECT 92.385 21.965 93.755 22.775 ;
        RECT 93.765 21.965 99.275 22.775 ;
        RECT 99.285 21.965 104.795 22.775 ;
        RECT 104.805 21.965 110.315 22.775 ;
        RECT 110.325 21.965 113.075 22.775 ;
        RECT 113.715 21.865 116.755 22.775 ;
        RECT 116.765 21.965 118.135 22.775 ;
        RECT 118.155 21.905 118.585 22.690 ;
        RECT 119.065 22.095 122.275 22.775 ;
        RECT 119.065 21.865 120.200 22.095 ;
        RECT 122.745 21.965 124.115 22.775 ;
      LAYER nwell ;
        RECT 92.190 18.745 124.310 21.575 ;
        RECT 128.520 21.010 132.230 23.770 ;
      LAYER pwell ;
        RECT 128.570 20.120 129.560 20.800 ;
        RECT 129.880 20.120 130.870 20.800 ;
        RECT 131.190 20.120 132.180 20.800 ;
        RECT 128.390 18.850 132.580 20.110 ;
        RECT 92.385 17.545 93.755 18.355 ;
        RECT 93.765 17.545 99.275 18.355 ;
        RECT 99.285 17.545 104.795 18.355 ;
        RECT 105.275 17.630 105.705 18.415 ;
        RECT 105.725 17.545 111.235 18.355 ;
        RECT 111.245 17.545 113.075 18.355 ;
        RECT 113.545 17.545 121.355 18.455 ;
        RECT 121.365 17.545 122.735 18.325 ;
        RECT 122.745 17.545 124.115 18.355 ;
        RECT 92.525 17.335 92.695 17.545 ;
        RECT 93.905 17.335 94.075 17.545 ;
        RECT 99.425 17.335 99.595 17.545 ;
        RECT 104.945 17.495 105.115 17.525 ;
        RECT 104.940 17.385 105.115 17.495 ;
        RECT 104.945 17.335 105.115 17.385 ;
        RECT 105.865 17.355 106.035 17.545 ;
        RECT 110.465 17.335 110.635 17.525 ;
        RECT 111.385 17.355 111.555 17.545 ;
        RECT 113.220 17.385 113.340 17.495 ;
        RECT 113.690 17.355 113.860 17.545 ;
        RECT 122.425 17.525 122.595 17.545 ;
        RECT 117.825 17.335 117.995 17.525 ;
        RECT 118.740 17.385 118.860 17.495 ;
        RECT 121.045 17.335 121.215 17.525 ;
        RECT 122.415 17.355 122.595 17.525 ;
        RECT 122.415 17.335 122.585 17.355 ;
        RECT 123.805 17.335 123.975 17.545 ;
        RECT 92.385 16.525 93.755 17.335 ;
        RECT 93.765 16.525 99.275 17.335 ;
        RECT 99.285 16.525 104.795 17.335 ;
        RECT 104.805 16.525 110.315 17.335 ;
        RECT 110.325 16.525 115.835 17.335 ;
        RECT 115.845 16.655 118.135 17.335 ;
        RECT 115.845 16.425 116.765 16.655 ;
        RECT 118.155 16.465 118.585 17.250 ;
        RECT 119.065 16.425 121.355 17.335 ;
        RECT 121.365 16.555 122.735 17.335 ;
        RECT 122.745 16.525 124.115 17.335 ;
      LAYER nwell ;
        RECT 92.190 13.305 124.310 16.135 ;
        RECT 128.520 16.090 132.230 18.850 ;
      LAYER pwell ;
        RECT 128.570 15.200 129.560 15.880 ;
        RECT 129.880 15.200 130.870 15.880 ;
        RECT 131.190 15.200 132.180 15.880 ;
        RECT 128.390 13.930 132.580 15.190 ;
        RECT 92.385 12.105 93.755 12.915 ;
        RECT 93.765 12.105 99.275 12.915 ;
        RECT 99.285 12.105 104.795 12.915 ;
        RECT 105.275 12.190 105.705 12.975 ;
        RECT 105.725 12.105 111.235 12.915 ;
        RECT 111.245 12.105 114.915 12.915 ;
        RECT 114.945 12.105 116.295 13.015 ;
        RECT 116.615 12.785 117.545 13.015 ;
        RECT 118.805 12.925 119.755 13.015 ;
        RECT 116.615 12.105 118.450 12.785 ;
        RECT 118.805 12.105 120.735 12.925 ;
        RECT 121.365 12.105 122.735 12.885 ;
        RECT 122.745 12.105 124.115 12.915 ;
        RECT 92.525 11.895 92.695 12.105 ;
        RECT 93.905 11.895 94.075 12.105 ;
        RECT 99.425 11.895 99.595 12.105 ;
        RECT 104.945 12.055 105.115 12.085 ;
        RECT 104.940 11.945 105.115 12.055 ;
        RECT 104.945 11.895 105.115 11.945 ;
        RECT 105.865 11.915 106.035 12.105 ;
        RECT 110.465 11.895 110.635 12.085 ;
        RECT 111.385 11.915 111.555 12.105 ;
        RECT 115.980 12.085 116.150 12.105 ;
        RECT 118.285 12.085 118.450 12.105 ;
        RECT 120.585 12.085 120.735 12.105 ;
        RECT 115.980 11.915 116.155 12.085 ;
        RECT 117.820 11.945 117.940 12.055 ;
        RECT 118.285 11.915 118.455 12.085 ;
        RECT 115.985 11.895 116.155 11.915 ;
        RECT 118.745 11.895 118.915 12.085 ;
        RECT 120.585 11.915 120.755 12.085 ;
        RECT 121.040 11.945 121.160 12.055 ;
        RECT 122.415 11.915 122.585 12.105 ;
        RECT 123.805 11.895 123.975 12.105 ;
        RECT 92.385 11.085 93.755 11.895 ;
        RECT 93.765 11.085 99.275 11.895 ;
        RECT 99.285 11.085 104.795 11.895 ;
        RECT 104.805 11.085 110.315 11.895 ;
        RECT 110.325 11.085 115.835 11.895 ;
        RECT 115.845 11.085 117.675 11.895 ;
        RECT 118.155 11.025 118.585 11.810 ;
        RECT 118.605 11.085 122.275 11.895 ;
        RECT 122.745 11.085 124.115 11.895 ;
      LAYER nwell ;
        RECT 128.520 11.170 132.230 13.930 ;
        RECT 92.190 7.865 124.310 10.695 ;
      LAYER pwell ;
        RECT 128.570 10.280 129.560 10.960 ;
        RECT 129.880 10.280 130.870 10.960 ;
        RECT 131.190 10.280 132.180 10.960 ;
        RECT 128.390 9.010 132.580 10.270 ;
        RECT 92.385 6.665 93.755 7.475 ;
        RECT 93.765 6.665 99.275 7.475 ;
        RECT 99.285 6.665 104.795 7.475 ;
        RECT 105.275 6.750 105.705 7.535 ;
        RECT 105.725 6.665 111.235 7.475 ;
        RECT 111.245 6.665 116.755 7.475 ;
        RECT 116.765 6.665 118.135 7.475 ;
        RECT 118.155 6.750 118.585 7.535 ;
        RECT 118.605 6.665 121.355 7.475 ;
        RECT 121.365 6.665 122.735 7.445 ;
        RECT 122.745 6.665 124.115 7.475 ;
        RECT 92.525 6.475 92.695 6.665 ;
        RECT 93.905 6.475 94.075 6.665 ;
        RECT 99.425 6.475 99.595 6.665 ;
        RECT 104.940 6.505 105.060 6.615 ;
        RECT 105.865 6.475 106.035 6.665 ;
        RECT 111.385 6.475 111.555 6.665 ;
        RECT 116.905 6.475 117.075 6.665 ;
        RECT 118.745 6.475 118.915 6.665 ;
        RECT 122.415 6.475 122.585 6.665 ;
        RECT 123.805 6.475 123.975 6.665 ;
      LAYER nwell ;
        RECT 128.520 6.250 132.230 9.010 ;
      LAYER pwell ;
        RECT 132.770 7.890 134.030 33.760 ;
        RECT 134.040 32.070 140.970 33.580 ;
        RECT 134.040 30.550 140.970 32.060 ;
        RECT 134.040 29.030 140.970 30.540 ;
        RECT 136.210 27.510 140.970 29.020 ;
      LAYER nwell ;
        RECT 141.180 28.980 152.880 33.630 ;
      LAYER pwell ;
        RECT 136.210 25.990 140.970 27.500 ;
      LAYER nwell ;
        RECT 141.550 26.030 152.880 28.980 ;
      LAYER pwell ;
        RECT 138.210 24.470 140.970 25.980 ;
        RECT 138.210 22.950 140.970 24.460 ;
        RECT 138.210 21.130 140.970 22.640 ;
        RECT 139.210 19.370 140.970 20.360 ;
      LAYER nwell ;
        RECT 141.180 18.840 152.880 26.030 ;
      LAYER pwell ;
        RECT 139.650 16.350 140.910 17.340 ;
        RECT 140.180 10.810 140.910 11.800 ;
      LAYER nwell ;
        RECT 141.120 8.280 152.880 18.840 ;
      LAYER pwell ;
        RECT 128.570 5.360 129.560 6.040 ;
        RECT 129.880 5.360 130.870 6.040 ;
        RECT 131.190 5.360 132.180 6.040 ;
        RECT 128.390 4.090 132.580 5.350 ;
      LAYER li1 ;
        RECT 128.520 37.430 132.450 38.290 ;
        RECT 92.380 36.395 124.120 36.565 ;
        RECT 92.465 35.305 93.675 36.395 ;
        RECT 93.845 35.960 99.190 36.395 ;
        RECT 99.365 35.960 104.710 36.395 ;
        RECT 92.465 34.595 92.985 35.135 ;
        RECT 93.155 34.765 93.675 35.305 ;
        RECT 92.465 33.845 93.675 34.595 ;
        RECT 95.430 34.390 95.770 35.220 ;
        RECT 97.250 34.710 97.600 35.960 ;
        RECT 100.950 34.390 101.290 35.220 ;
        RECT 102.770 34.710 103.120 35.960 ;
        RECT 105.345 35.230 105.635 36.395 ;
        RECT 105.805 35.960 111.150 36.395 ;
        RECT 111.325 35.960 116.670 36.395 ;
        RECT 93.845 33.845 99.190 34.390 ;
        RECT 99.365 33.845 104.710 34.390 ;
        RECT 105.345 33.845 105.635 34.570 ;
        RECT 107.390 34.390 107.730 35.220 ;
        RECT 109.210 34.710 109.560 35.960 ;
        RECT 112.910 34.390 113.250 35.220 ;
        RECT 114.730 34.710 115.080 35.960 ;
        RECT 116.845 35.305 118.055 36.395 ;
        RECT 116.845 34.595 117.365 35.135 ;
        RECT 117.535 34.765 118.055 35.305 ;
        RECT 118.225 35.230 118.515 36.395 ;
        RECT 118.685 35.305 119.895 36.395 ;
        RECT 118.685 34.595 119.205 35.135 ;
        RECT 119.375 34.765 119.895 35.305 ;
        RECT 120.065 35.320 120.335 36.225 ;
        RECT 120.505 35.635 120.835 36.395 ;
        RECT 121.015 35.465 121.195 36.225 ;
        RECT 105.805 33.845 111.150 34.390 ;
        RECT 111.325 33.845 116.670 34.390 ;
        RECT 116.845 33.845 118.055 34.595 ;
        RECT 118.225 33.845 118.515 34.570 ;
        RECT 118.685 33.845 119.895 34.595 ;
        RECT 120.065 34.520 120.245 35.320 ;
        RECT 120.520 35.295 121.195 35.465 ;
        RECT 121.445 35.320 121.715 36.225 ;
        RECT 121.885 35.635 122.215 36.395 ;
        RECT 122.395 35.465 122.575 36.225 ;
        RECT 120.520 35.150 120.690 35.295 ;
        RECT 120.415 34.820 120.690 35.150 ;
        RECT 120.520 34.565 120.690 34.820 ;
        RECT 120.915 34.745 121.255 35.115 ;
        RECT 120.065 34.015 120.325 34.520 ;
        RECT 120.520 34.395 121.185 34.565 ;
        RECT 120.505 33.845 120.835 34.225 ;
        RECT 121.015 34.015 121.185 34.395 ;
        RECT 121.445 34.520 121.625 35.320 ;
        RECT 121.900 35.295 122.575 35.465 ;
        RECT 122.825 35.305 124.035 36.395 ;
        RECT 128.240 35.830 128.570 35.900 ;
        RECT 128.760 35.830 128.930 37.110 ;
        RECT 129.200 36.070 129.370 37.430 ;
        RECT 128.240 35.630 128.930 35.830 ;
        RECT 128.240 35.560 128.570 35.630 ;
        RECT 121.900 35.150 122.070 35.295 ;
        RECT 121.795 34.820 122.070 35.150 ;
        RECT 121.900 34.565 122.070 34.820 ;
        RECT 122.295 34.745 122.635 35.115 ;
        RECT 122.825 34.765 123.345 35.305 ;
        RECT 123.515 34.595 124.035 35.135 ;
        RECT 128.760 35.000 128.930 35.630 ;
        RECT 129.500 35.830 129.830 35.910 ;
        RECT 130.070 35.830 130.240 37.110 ;
        RECT 130.510 36.070 130.680 37.430 ;
        RECT 129.500 35.630 130.240 35.830 ;
        RECT 129.500 35.570 129.830 35.630 ;
        RECT 129.200 34.670 129.370 35.460 ;
        RECT 130.070 35.000 130.240 35.630 ;
        RECT 130.810 35.830 131.140 35.910 ;
        RECT 131.380 35.830 131.550 37.110 ;
        RECT 131.820 36.070 131.990 37.430 ;
        RECT 130.810 35.630 131.550 35.830 ;
        RECT 130.810 35.570 131.140 35.630 ;
        RECT 130.510 34.670 130.680 35.460 ;
        RECT 131.380 35.000 131.550 35.630 ;
        RECT 132.120 35.570 132.450 35.910 ;
        RECT 131.820 34.670 131.990 35.460 ;
        RECT 121.445 34.015 121.705 34.520 ;
        RECT 121.900 34.395 122.565 34.565 ;
        RECT 121.885 33.845 122.215 34.225 ;
        RECT 122.395 34.015 122.565 34.395 ;
        RECT 122.825 33.845 124.035 34.595 ;
        RECT 92.380 33.675 124.120 33.845 ;
        RECT 128.520 33.830 132.450 34.670 ;
        RECT 92.465 32.925 93.675 33.675 ;
        RECT 93.845 33.130 99.190 33.675 ;
        RECT 99.365 33.130 104.710 33.675 ;
        RECT 104.885 33.130 110.230 33.675 ;
        RECT 110.405 33.130 115.750 33.675 ;
        RECT 92.465 32.385 92.985 32.925 ;
        RECT 93.155 32.215 93.675 32.755 ;
        RECT 95.430 32.300 95.770 33.130 ;
        RECT 92.465 31.125 93.675 32.215 ;
        RECT 97.250 31.560 97.600 32.810 ;
        RECT 100.950 32.300 101.290 33.130 ;
        RECT 102.770 31.560 103.120 32.810 ;
        RECT 106.470 32.300 106.810 33.130 ;
        RECT 108.290 31.560 108.640 32.810 ;
        RECT 111.990 32.300 112.330 33.130 ;
        RECT 115.925 32.905 117.595 33.675 ;
        RECT 118.225 32.950 118.515 33.675 ;
        RECT 118.685 32.905 122.195 33.675 ;
        RECT 122.825 32.925 124.035 33.675 ;
        RECT 132.980 33.390 133.820 33.630 ;
        RECT 113.810 31.560 114.160 32.810 ;
        RECT 115.925 32.385 116.675 32.905 ;
        RECT 116.845 32.215 117.595 32.735 ;
        RECT 118.685 32.385 120.335 32.905 ;
        RECT 93.845 31.125 99.190 31.560 ;
        RECT 99.365 31.125 104.710 31.560 ;
        RECT 104.885 31.125 110.230 31.560 ;
        RECT 110.405 31.125 115.750 31.560 ;
        RECT 115.925 31.125 117.595 32.215 ;
        RECT 118.225 31.125 118.515 32.290 ;
        RECT 120.505 32.215 122.195 32.735 ;
        RECT 118.685 31.125 122.195 32.215 ;
        RECT 122.825 32.215 123.345 32.755 ;
        RECT 123.515 32.385 124.035 32.925 ;
        RECT 128.520 32.510 132.450 33.370 ;
        RECT 132.980 33.220 140.860 33.390 ;
        RECT 122.825 31.125 124.035 32.215 ;
        RECT 92.380 30.955 124.120 31.125 ;
        RECT 92.465 29.865 93.675 30.955 ;
        RECT 93.845 30.520 99.190 30.955 ;
        RECT 99.365 30.520 104.710 30.955 ;
        RECT 92.465 29.155 92.985 29.695 ;
        RECT 93.155 29.325 93.675 29.865 ;
        RECT 92.465 28.405 93.675 29.155 ;
        RECT 95.430 28.950 95.770 29.780 ;
        RECT 97.250 29.270 97.600 30.520 ;
        RECT 100.950 28.950 101.290 29.780 ;
        RECT 102.770 29.270 103.120 30.520 ;
        RECT 105.345 29.790 105.635 30.955 ;
        RECT 105.805 30.520 111.150 30.955 ;
        RECT 111.325 30.520 116.670 30.955 ;
        RECT 93.845 28.405 99.190 28.950 ;
        RECT 99.365 28.405 104.710 28.950 ;
        RECT 105.345 28.405 105.635 29.130 ;
        RECT 107.390 28.950 107.730 29.780 ;
        RECT 109.210 29.270 109.560 30.520 ;
        RECT 112.910 28.950 113.250 29.780 ;
        RECT 114.730 29.270 115.080 30.520 ;
        RECT 116.845 29.865 120.355 30.955 ;
        RECT 116.845 29.175 118.495 29.695 ;
        RECT 118.665 29.345 120.355 29.865 ;
        RECT 121.445 29.880 121.715 30.785 ;
        RECT 121.885 30.195 122.215 30.955 ;
        RECT 122.395 30.025 122.565 30.785 ;
        RECT 105.805 28.405 111.150 28.950 ;
        RECT 111.325 28.405 116.670 28.950 ;
        RECT 116.845 28.405 120.355 29.175 ;
        RECT 121.445 29.080 121.615 29.880 ;
        RECT 121.900 29.855 122.565 30.025 ;
        RECT 122.825 29.865 124.035 30.955 ;
        RECT 128.240 30.910 128.570 30.960 ;
        RECT 128.760 30.910 128.930 32.190 ;
        RECT 129.200 31.150 129.370 32.510 ;
        RECT 128.240 30.710 128.930 30.910 ;
        RECT 128.240 30.620 128.570 30.710 ;
        RECT 128.760 30.080 128.930 30.710 ;
        RECT 129.500 30.910 129.830 30.990 ;
        RECT 130.070 30.910 130.240 32.190 ;
        RECT 130.510 31.150 130.680 32.510 ;
        RECT 129.500 30.710 130.240 30.910 ;
        RECT 129.500 30.650 129.830 30.710 ;
        RECT 121.900 29.710 122.070 29.855 ;
        RECT 121.785 29.380 122.070 29.710 ;
        RECT 121.900 29.125 122.070 29.380 ;
        RECT 122.305 29.305 122.635 29.675 ;
        RECT 122.825 29.325 123.345 29.865 ;
        RECT 129.200 29.750 129.370 30.540 ;
        RECT 130.070 30.080 130.240 30.710 ;
        RECT 130.810 30.910 131.140 30.990 ;
        RECT 131.380 30.910 131.550 32.190 ;
        RECT 131.820 31.150 131.990 32.510 ;
        RECT 132.980 32.430 133.820 33.220 ;
        RECT 141.030 33.120 141.360 33.450 ;
        RECT 134.150 32.740 141.230 32.910 ;
        RECT 132.980 32.260 140.860 32.430 ;
        RECT 132.980 31.870 133.820 32.260 ;
        RECT 132.980 31.700 140.860 31.870 ;
        RECT 130.810 30.710 131.550 30.910 ;
        RECT 130.810 30.650 131.140 30.710 ;
        RECT 130.510 29.750 130.680 30.540 ;
        RECT 131.380 30.080 131.550 30.710 ;
        RECT 132.120 30.650 132.450 30.990 ;
        RECT 132.980 30.910 133.820 31.700 ;
        RECT 141.030 31.390 141.230 32.740 ;
        RECT 151.770 31.830 152.630 33.630 ;
        RECT 141.470 31.660 152.630 31.830 ;
        RECT 134.150 31.220 141.980 31.390 ;
        RECT 132.980 30.740 140.860 30.910 ;
        RECT 131.820 29.750 131.990 30.540 ;
        RECT 132.980 30.350 133.820 30.740 ;
        RECT 132.980 30.180 140.860 30.350 ;
        RECT 123.515 29.155 124.035 29.695 ;
        RECT 121.445 28.575 121.705 29.080 ;
        RECT 121.900 28.955 122.565 29.125 ;
        RECT 121.885 28.405 122.215 28.785 ;
        RECT 122.395 28.575 122.565 28.955 ;
        RECT 122.825 28.405 124.035 29.155 ;
        RECT 128.520 28.910 132.450 29.750 ;
        RECT 132.980 29.390 133.820 30.180 ;
        RECT 141.030 29.870 141.230 31.220 ;
        RECT 134.150 29.700 141.230 29.870 ;
        RECT 141.030 29.490 141.230 29.700 ;
        RECT 132.980 29.220 140.860 29.390 ;
        RECT 132.980 28.830 133.820 29.220 ;
        RECT 141.030 29.160 141.360 29.490 ;
        RECT 132.980 28.660 140.860 28.830 ;
        RECT 92.380 28.235 124.120 28.405 ;
        RECT 92.465 27.485 93.675 28.235 ;
        RECT 93.845 27.690 99.190 28.235 ;
        RECT 99.365 27.690 104.710 28.235 ;
        RECT 104.885 27.690 110.230 28.235 ;
        RECT 110.405 27.690 115.750 28.235 ;
        RECT 115.925 27.855 116.815 28.025 ;
        RECT 92.465 26.945 92.985 27.485 ;
        RECT 93.155 26.775 93.675 27.315 ;
        RECT 95.430 26.860 95.770 27.690 ;
        RECT 92.465 25.685 93.675 26.775 ;
        RECT 97.250 26.120 97.600 27.370 ;
        RECT 100.950 26.860 101.290 27.690 ;
        RECT 102.770 26.120 103.120 27.370 ;
        RECT 106.470 26.860 106.810 27.690 ;
        RECT 108.290 26.120 108.640 27.370 ;
        RECT 111.990 26.860 112.330 27.690 ;
        RECT 113.810 26.120 114.160 27.370 ;
        RECT 115.925 27.300 116.475 27.685 ;
        RECT 116.645 27.130 116.815 27.855 ;
        RECT 115.925 27.060 116.815 27.130 ;
        RECT 116.985 27.555 117.205 28.015 ;
        RECT 117.375 27.695 117.625 28.235 ;
        RECT 117.795 27.585 118.055 28.065 ;
        RECT 116.985 27.530 117.235 27.555 ;
        RECT 116.985 27.105 117.315 27.530 ;
        RECT 115.925 27.035 116.820 27.060 ;
        RECT 115.925 27.020 116.830 27.035 ;
        RECT 115.925 27.005 116.835 27.020 ;
        RECT 115.925 27.000 116.845 27.005 ;
        RECT 115.925 26.990 116.850 27.000 ;
        RECT 115.925 26.980 116.855 26.990 ;
        RECT 115.925 26.975 116.865 26.980 ;
        RECT 115.925 26.965 116.875 26.975 ;
        RECT 115.925 26.960 116.885 26.965 ;
        RECT 115.925 26.510 116.185 26.960 ;
        RECT 116.550 26.955 116.885 26.960 ;
        RECT 116.550 26.950 116.900 26.955 ;
        RECT 116.550 26.940 116.915 26.950 ;
        RECT 116.550 26.935 116.940 26.940 ;
        RECT 117.485 26.935 117.715 27.330 ;
        RECT 116.550 26.930 117.715 26.935 ;
        RECT 116.580 26.895 117.715 26.930 ;
        RECT 116.615 26.870 117.715 26.895 ;
        RECT 116.645 26.840 117.715 26.870 ;
        RECT 116.665 26.810 117.715 26.840 ;
        RECT 116.685 26.780 117.715 26.810 ;
        RECT 116.755 26.770 117.715 26.780 ;
        RECT 116.780 26.760 117.715 26.770 ;
        RECT 116.800 26.745 117.715 26.760 ;
        RECT 116.820 26.730 117.715 26.745 ;
        RECT 116.825 26.720 117.610 26.730 ;
        RECT 116.840 26.685 117.610 26.720 ;
        RECT 116.355 26.365 116.685 26.610 ;
        RECT 116.855 26.435 117.610 26.685 ;
        RECT 117.885 26.555 118.055 27.585 ;
        RECT 118.225 27.510 118.515 28.235 ;
        RECT 116.355 26.340 116.540 26.365 ;
        RECT 115.925 26.240 116.540 26.340 ;
        RECT 93.845 25.685 99.190 26.120 ;
        RECT 99.365 25.685 104.710 26.120 ;
        RECT 104.885 25.685 110.230 26.120 ;
        RECT 110.405 25.685 115.750 26.120 ;
        RECT 115.925 25.685 116.530 26.240 ;
        RECT 116.705 25.855 117.185 26.195 ;
        RECT 117.355 25.685 117.610 26.230 ;
        RECT 117.780 25.855 118.055 26.555 ;
        RECT 118.225 25.685 118.515 26.850 ;
        RECT 118.695 25.865 118.955 28.055 ;
        RECT 119.215 27.865 119.885 28.235 ;
        RECT 120.065 27.685 120.375 28.055 ;
        RECT 119.145 27.485 120.375 27.685 ;
        RECT 119.145 26.815 119.435 27.485 ;
        RECT 120.555 27.305 120.785 27.945 ;
        RECT 120.965 27.505 121.255 28.235 ;
        RECT 121.465 27.425 121.705 28.235 ;
        RECT 121.875 27.425 122.205 28.065 ;
        RECT 122.375 27.425 122.645 28.235 ;
        RECT 122.825 27.485 124.035 28.235 ;
        RECT 128.520 27.580 132.450 28.440 ;
        RECT 132.980 27.870 133.820 28.660 ;
        RECT 141.030 28.560 141.360 28.890 ;
        RECT 136.320 28.180 141.230 28.350 ;
        RECT 132.980 27.700 140.860 27.870 ;
        RECT 119.615 26.995 120.080 27.305 ;
        RECT 120.260 26.995 120.785 27.305 ;
        RECT 120.965 26.995 121.265 27.325 ;
        RECT 121.445 26.995 121.795 27.245 ;
        RECT 121.965 26.825 122.135 27.425 ;
        RECT 122.305 26.995 122.655 27.245 ;
        RECT 119.145 26.595 119.915 26.815 ;
        RECT 119.125 25.685 119.465 26.415 ;
        RECT 119.645 25.865 119.915 26.595 ;
        RECT 120.095 26.575 121.255 26.815 ;
        RECT 120.095 25.865 120.325 26.575 ;
        RECT 120.495 25.685 120.825 26.395 ;
        RECT 120.995 25.865 121.255 26.575 ;
        RECT 121.455 26.655 122.135 26.825 ;
        RECT 121.455 25.870 121.785 26.655 ;
        RECT 122.315 25.685 122.645 26.825 ;
        RECT 122.825 26.775 123.345 27.315 ;
        RECT 123.515 26.945 124.035 27.485 ;
        RECT 122.825 25.685 124.035 26.775 ;
        RECT 128.240 25.980 128.570 26.050 ;
        RECT 128.760 25.980 128.930 27.260 ;
        RECT 129.200 26.220 129.370 27.580 ;
        RECT 128.240 25.780 128.930 25.980 ;
        RECT 128.240 25.710 128.570 25.780 ;
        RECT 92.380 25.515 124.120 25.685 ;
        RECT 92.465 24.425 93.675 25.515 ;
        RECT 93.845 25.080 99.190 25.515 ;
        RECT 99.365 25.080 104.710 25.515 ;
        RECT 92.465 23.715 92.985 24.255 ;
        RECT 93.155 23.885 93.675 24.425 ;
        RECT 92.465 22.965 93.675 23.715 ;
        RECT 95.430 23.510 95.770 24.340 ;
        RECT 97.250 23.830 97.600 25.080 ;
        RECT 100.950 23.510 101.290 24.340 ;
        RECT 102.770 23.830 103.120 25.080 ;
        RECT 105.345 24.350 105.635 25.515 ;
        RECT 105.805 25.080 111.150 25.515 ;
        RECT 93.845 22.965 99.190 23.510 ;
        RECT 99.365 22.965 104.710 23.510 ;
        RECT 105.345 22.965 105.635 23.690 ;
        RECT 107.390 23.510 107.730 24.340 ;
        RECT 109.210 23.830 109.560 25.080 ;
        RECT 111.325 24.425 113.915 25.515 ;
        RECT 114.795 25.005 115.125 25.515 ;
        RECT 115.295 24.835 115.465 25.345 ;
        RECT 115.635 25.005 115.965 25.515 ;
        RECT 116.135 24.835 116.305 25.345 ;
        RECT 116.475 25.005 116.805 25.515 ;
        RECT 117.075 25.175 118.085 25.345 ;
        RECT 111.325 23.735 112.535 24.255 ;
        RECT 112.705 23.905 113.915 24.425 ;
        RECT 114.605 24.665 116.365 24.835 ;
        RECT 117.075 24.675 117.245 25.175 ;
        RECT 105.805 22.965 111.150 23.510 ;
        RECT 111.325 22.965 113.915 23.735 ;
        RECT 114.605 23.705 114.775 24.665 ;
        RECT 117.415 24.505 117.745 24.995 ;
        RECT 117.915 24.835 118.085 25.175 ;
        RECT 118.375 25.005 118.705 25.515 ;
        RECT 118.875 24.835 119.045 25.345 ;
        RECT 119.215 25.005 119.545 25.515 ;
        RECT 119.715 24.835 119.885 25.345 ;
        RECT 120.055 25.005 120.385 25.515 ;
        RECT 120.555 24.835 120.725 25.345 ;
        RECT 117.915 24.665 120.725 24.835 ;
        RECT 116.505 24.335 117.745 24.505 ;
        RECT 116.505 24.205 116.675 24.335 ;
        RECT 114.965 23.875 116.675 24.205 ;
        RECT 116.870 23.955 117.325 24.165 ;
        RECT 114.605 23.535 116.395 23.705 ;
        RECT 116.870 23.625 117.085 23.955 ;
        RECT 117.555 23.750 117.745 24.335 ;
        RECT 118.045 24.325 120.750 24.495 ;
        RECT 118.045 23.955 118.375 24.325 ;
        RECT 120.375 24.155 120.750 24.325 ;
        RECT 121.445 24.440 121.715 25.345 ;
        RECT 121.885 24.755 122.215 25.515 ;
        RECT 122.395 24.585 122.565 25.345 ;
        RECT 118.585 23.955 118.915 24.155 ;
        RECT 119.195 23.955 119.545 24.155 ;
        RECT 119.845 23.955 120.175 24.125 ;
        RECT 120.375 23.985 120.755 24.155 ;
        RECT 120.375 23.955 120.750 23.985 ;
        RECT 118.730 23.785 118.915 23.955 ;
        RECT 119.925 23.785 120.095 23.955 ;
        RECT 117.555 23.685 118.550 23.750 ;
        RECT 117.415 23.580 118.550 23.685 ;
        RECT 118.730 23.615 120.095 23.785 ;
        RECT 114.795 22.965 115.125 23.365 ;
        RECT 115.635 22.965 115.965 23.365 ;
        RECT 116.635 22.965 117.165 23.445 ;
        RECT 117.415 23.175 117.745 23.580 ;
        RECT 118.380 23.445 118.550 23.580 ;
        RECT 117.915 22.965 118.200 23.410 ;
        RECT 118.380 23.275 119.545 23.445 ;
        RECT 120.555 22.965 120.725 23.785 ;
        RECT 121.445 23.640 121.615 24.440 ;
        RECT 121.900 24.415 122.565 24.585 ;
        RECT 122.825 24.425 124.035 25.515 ;
        RECT 128.760 25.150 128.930 25.780 ;
        RECT 129.500 25.980 129.830 26.060 ;
        RECT 130.070 25.980 130.240 27.260 ;
        RECT 130.510 26.220 130.680 27.580 ;
        RECT 129.500 25.780 130.240 25.980 ;
        RECT 129.500 25.720 129.830 25.780 ;
        RECT 129.200 24.830 129.370 25.610 ;
        RECT 130.070 25.150 130.240 25.780 ;
        RECT 130.810 25.980 131.140 26.060 ;
        RECT 131.380 25.980 131.550 27.260 ;
        RECT 131.820 26.220 131.990 27.580 ;
        RECT 132.980 27.310 133.820 27.700 ;
        RECT 141.030 27.590 141.230 28.180 ;
        RECT 151.770 28.030 152.630 31.660 ;
        RECT 141.840 27.860 152.630 28.030 ;
        RECT 141.030 27.420 143.880 27.590 ;
        RECT 132.980 27.140 140.860 27.310 ;
        RECT 132.980 26.350 133.820 27.140 ;
        RECT 141.030 26.830 141.230 27.420 ;
        RECT 136.320 26.660 141.230 26.830 ;
        RECT 141.030 26.450 141.230 26.660 ;
        RECT 132.980 26.180 140.860 26.350 ;
        RECT 130.810 25.780 131.550 25.980 ;
        RECT 130.810 25.720 131.140 25.780 ;
        RECT 130.510 24.830 130.680 25.610 ;
        RECT 131.380 25.150 131.550 25.780 ;
        RECT 132.120 25.720 132.450 26.060 ;
        RECT 132.980 25.790 133.820 26.180 ;
        RECT 141.030 26.120 141.360 26.450 ;
        RECT 132.980 25.620 140.860 25.790 ;
        RECT 131.820 24.830 131.990 25.610 ;
        RECT 132.980 24.830 133.820 25.620 ;
        RECT 141.030 25.520 141.360 25.850 ;
        RECT 138.320 25.140 141.230 25.310 ;
        RECT 121.900 24.270 122.070 24.415 ;
        RECT 121.785 23.940 122.070 24.270 ;
        RECT 121.900 23.685 122.070 23.940 ;
        RECT 122.305 23.865 122.635 24.235 ;
        RECT 122.825 23.885 123.345 24.425 ;
        RECT 123.515 23.715 124.035 24.255 ;
        RECT 128.510 23.980 132.460 24.830 ;
        RECT 132.980 24.660 140.860 24.830 ;
        RECT 132.980 24.270 133.820 24.660 ;
        RECT 141.030 24.550 141.230 25.140 ;
        RECT 151.770 24.990 152.630 27.860 ;
        RECT 141.470 24.820 152.630 24.990 ;
        RECT 141.030 24.380 148.510 24.550 ;
        RECT 132.980 24.100 140.860 24.270 ;
        RECT 121.445 23.135 121.705 23.640 ;
        RECT 121.900 23.515 122.565 23.685 ;
        RECT 121.885 22.965 122.215 23.345 ;
        RECT 122.395 23.135 122.565 23.515 ;
        RECT 122.825 22.965 124.035 23.715 ;
        RECT 92.380 22.795 124.120 22.965 ;
        RECT 92.465 22.045 93.675 22.795 ;
        RECT 93.845 22.250 99.190 22.795 ;
        RECT 99.365 22.250 104.710 22.795 ;
        RECT 104.885 22.250 110.230 22.795 ;
        RECT 92.465 21.505 92.985 22.045 ;
        RECT 93.155 21.335 93.675 21.875 ;
        RECT 95.430 21.420 95.770 22.250 ;
        RECT 92.465 20.245 93.675 21.335 ;
        RECT 97.250 20.680 97.600 21.930 ;
        RECT 100.950 21.420 101.290 22.250 ;
        RECT 102.770 20.680 103.120 21.930 ;
        RECT 106.470 21.420 106.810 22.250 ;
        RECT 110.405 22.025 112.995 22.795 ;
        RECT 113.805 22.415 114.135 22.795 ;
        RECT 114.305 22.245 114.495 22.625 ;
        RECT 114.665 22.435 114.995 22.795 ;
        RECT 114.095 22.055 114.495 22.245 ;
        RECT 115.215 22.225 115.405 22.625 ;
        RECT 114.665 22.055 115.405 22.225 ;
        RECT 108.290 20.680 108.640 21.930 ;
        RECT 110.405 21.505 111.615 22.025 ;
        RECT 111.785 21.335 112.995 21.855 ;
        RECT 93.845 20.245 99.190 20.680 ;
        RECT 99.365 20.245 104.710 20.680 ;
        RECT 104.885 20.245 110.230 20.680 ;
        RECT 110.405 20.245 112.995 21.335 ;
        RECT 113.635 20.245 113.925 21.215 ;
        RECT 114.095 20.415 114.325 22.055 ;
        RECT 114.665 21.885 114.835 22.055 ;
        RECT 114.495 21.190 114.835 21.885 ;
        RECT 115.005 21.470 115.330 21.885 ;
        RECT 115.780 21.555 116.160 22.515 ;
        RECT 116.345 22.315 116.675 22.795 ;
        RECT 116.350 21.555 116.665 22.130 ;
        RECT 116.845 22.045 118.055 22.795 ;
        RECT 118.225 22.070 118.515 22.795 ;
        RECT 119.145 22.075 119.485 22.585 ;
        RECT 116.845 21.505 117.365 22.045 ;
        RECT 117.535 21.335 118.055 21.875 ;
        RECT 114.495 20.960 115.330 21.190 ;
        RECT 114.495 20.245 114.825 20.660 ;
        RECT 115.015 20.415 115.330 20.960 ;
        RECT 115.500 20.945 116.615 21.210 ;
        RECT 115.500 20.415 115.725 20.945 ;
        RECT 115.895 20.245 116.225 20.755 ;
        RECT 116.395 20.415 116.615 20.945 ;
        RECT 116.845 20.245 118.055 21.335 ;
        RECT 118.225 20.245 118.515 21.410 ;
        RECT 119.145 20.675 119.405 22.075 ;
        RECT 119.655 21.995 119.925 22.795 ;
        RECT 119.580 21.555 119.910 21.805 ;
        RECT 120.105 21.555 120.385 22.525 ;
        RECT 120.565 21.555 120.865 22.525 ;
        RECT 121.045 21.555 121.395 22.520 ;
        RECT 121.615 22.295 122.110 22.625 ;
        RECT 119.595 21.385 119.910 21.555 ;
        RECT 121.615 21.385 121.785 22.295 ;
        RECT 119.595 21.215 121.785 21.385 ;
        RECT 119.145 20.415 119.485 20.675 ;
        RECT 119.655 20.245 119.985 21.045 ;
        RECT 120.450 20.415 120.700 21.215 ;
        RECT 120.885 20.245 121.215 20.965 ;
        RECT 121.435 20.415 121.685 21.215 ;
        RECT 121.955 20.805 122.195 22.115 ;
        RECT 122.825 22.045 124.035 22.795 ;
        RECT 128.520 22.660 132.450 23.520 ;
        RECT 132.980 23.310 133.820 24.100 ;
        RECT 141.030 23.790 141.230 24.380 ;
        RECT 138.320 23.620 141.230 23.790 ;
        RECT 141.030 23.410 141.230 23.620 ;
        RECT 132.980 23.140 140.860 23.310 ;
        RECT 122.825 21.335 123.345 21.875 ;
        RECT 123.515 21.505 124.035 22.045 ;
        RECT 121.855 20.245 122.190 20.625 ;
        RECT 122.825 20.245 124.035 21.335 ;
        RECT 128.240 21.060 128.570 21.130 ;
        RECT 128.760 21.060 128.930 22.340 ;
        RECT 129.200 21.300 129.370 22.660 ;
        RECT 128.240 20.860 128.930 21.060 ;
        RECT 128.240 20.790 128.570 20.860 ;
        RECT 92.380 20.075 124.120 20.245 ;
        RECT 128.760 20.230 128.930 20.860 ;
        RECT 129.500 21.060 129.830 21.140 ;
        RECT 130.070 21.060 130.240 22.340 ;
        RECT 130.510 21.300 130.680 22.660 ;
        RECT 129.500 20.860 130.240 21.060 ;
        RECT 129.500 20.800 129.830 20.860 ;
        RECT 92.465 18.985 93.675 20.075 ;
        RECT 93.845 19.640 99.190 20.075 ;
        RECT 99.365 19.640 104.710 20.075 ;
        RECT 92.465 18.275 92.985 18.815 ;
        RECT 93.155 18.445 93.675 18.985 ;
        RECT 92.465 17.525 93.675 18.275 ;
        RECT 95.430 18.070 95.770 18.900 ;
        RECT 97.250 18.390 97.600 19.640 ;
        RECT 100.950 18.070 101.290 18.900 ;
        RECT 102.770 18.390 103.120 19.640 ;
        RECT 105.345 18.910 105.635 20.075 ;
        RECT 105.805 19.640 111.150 20.075 ;
        RECT 93.845 17.525 99.190 18.070 ;
        RECT 99.365 17.525 104.710 18.070 ;
        RECT 105.345 17.525 105.635 18.250 ;
        RECT 107.390 18.070 107.730 18.900 ;
        RECT 109.210 18.390 109.560 19.640 ;
        RECT 111.325 18.985 112.995 20.075 ;
        RECT 113.635 19.355 113.965 20.075 ;
        RECT 114.135 19.105 114.305 19.905 ;
        RECT 114.475 19.355 114.805 20.075 ;
        RECT 114.975 19.105 115.145 19.905 ;
        RECT 115.315 19.355 115.645 20.075 ;
        RECT 115.815 19.525 115.985 19.905 ;
        RECT 116.155 19.695 116.485 20.075 ;
        RECT 116.755 19.525 116.925 19.905 ;
        RECT 117.095 19.695 117.425 20.075 ;
        RECT 117.595 19.525 117.765 19.905 ;
        RECT 117.935 19.695 118.265 20.075 ;
        RECT 118.435 19.695 121.265 19.865 ;
        RECT 118.435 19.525 118.605 19.695 ;
        RECT 115.815 19.355 118.605 19.525 ;
        RECT 119.675 19.515 120.845 19.525 ;
        RECT 118.820 19.355 120.845 19.515 ;
        RECT 118.820 19.345 119.740 19.355 ;
        RECT 118.820 19.105 118.990 19.345 ;
        RECT 121.015 19.195 121.265 19.695 ;
        RECT 111.325 18.295 112.075 18.815 ;
        RECT 112.245 18.465 112.995 18.985 ;
        RECT 113.660 18.935 115.145 19.105 ;
        RECT 115.340 18.935 118.990 19.105 ;
        RECT 105.805 17.525 111.150 18.070 ;
        RECT 111.325 17.525 112.995 18.295 ;
        RECT 113.660 18.245 113.880 18.935 ;
        RECT 115.340 18.765 115.510 18.935 ;
        RECT 114.110 18.435 115.510 18.765 ;
        RECT 115.750 18.515 116.645 18.735 ;
        RECT 116.875 18.515 117.570 18.765 ;
        RECT 117.820 18.515 118.615 18.765 ;
        RECT 113.660 18.075 115.145 18.245 ;
        RECT 113.635 17.525 113.965 17.905 ;
        RECT 114.135 17.695 114.305 18.075 ;
        RECT 114.475 17.525 114.805 17.905 ;
        RECT 114.975 17.695 115.145 18.075 ;
        RECT 115.815 18.095 117.425 18.265 ;
        RECT 118.820 18.245 118.990 18.935 ;
        RECT 119.170 18.515 120.320 19.065 ;
        RECT 120.570 18.735 120.765 19.075 ;
        RECT 121.445 19.000 121.715 19.905 ;
        RECT 121.885 19.315 122.215 20.075 ;
        RECT 122.395 19.145 122.565 19.905 ;
        RECT 120.570 18.515 121.250 18.735 ;
        RECT 115.315 17.525 115.645 17.905 ;
        RECT 115.815 17.695 115.985 18.095 ;
        RECT 117.935 18.075 119.965 18.245 ;
        RECT 120.175 18.085 121.185 18.255 ;
        RECT 120.175 17.905 120.345 18.085 ;
        RECT 116.155 17.525 116.485 17.905 ;
        RECT 116.675 17.735 118.685 17.905 ;
        RECT 119.210 17.735 120.345 17.905 ;
        RECT 120.175 17.695 120.345 17.735 ;
        RECT 120.515 17.525 120.845 17.905 ;
        RECT 121.015 17.695 121.185 18.085 ;
        RECT 121.445 18.200 121.615 19.000 ;
        RECT 121.900 18.975 122.565 19.145 ;
        RECT 122.825 18.985 124.035 20.075 ;
        RECT 129.200 19.900 129.370 20.690 ;
        RECT 130.070 20.230 130.240 20.860 ;
        RECT 130.810 21.060 131.140 21.140 ;
        RECT 131.380 21.060 131.550 22.340 ;
        RECT 131.820 21.300 131.990 22.660 ;
        RECT 132.980 22.450 133.820 23.140 ;
        RECT 141.030 23.080 141.360 23.410 ;
        RECT 141.030 22.580 141.360 22.910 ;
        RECT 151.770 22.450 152.630 24.820 ;
        RECT 132.980 22.280 140.860 22.450 ;
        RECT 141.470 22.280 152.630 22.450 ;
        RECT 132.980 21.490 133.820 22.280 ;
        RECT 138.320 21.800 149.010 21.970 ;
        RECT 132.980 21.320 140.860 21.490 ;
        RECT 130.810 20.860 131.550 21.060 ;
        RECT 130.810 20.800 131.140 20.860 ;
        RECT 130.510 19.900 130.680 20.690 ;
        RECT 131.380 20.230 131.550 20.860 ;
        RECT 132.120 20.800 132.450 21.140 ;
        RECT 131.820 19.900 131.990 20.690 ;
        RECT 132.980 20.170 133.820 21.320 ;
        RECT 141.030 21.170 141.230 21.800 ;
        RECT 151.770 21.490 152.630 22.280 ;
        RECT 141.470 21.320 152.630 21.490 ;
        RECT 141.030 20.840 141.360 21.170 ;
        RECT 141.030 20.340 141.360 20.670 ;
        RECT 151.770 20.210 152.630 21.320 ;
        RECT 132.980 20.000 140.860 20.170 ;
        RECT 141.470 20.040 152.630 20.210 ;
        RECT 128.520 19.050 132.450 19.900 ;
        RECT 121.900 18.830 122.070 18.975 ;
        RECT 121.785 18.500 122.070 18.830 ;
        RECT 121.900 18.245 122.070 18.500 ;
        RECT 122.305 18.425 122.635 18.795 ;
        RECT 122.825 18.445 123.345 18.985 ;
        RECT 123.515 18.275 124.035 18.815 ;
        RECT 121.445 17.695 121.705 18.200 ;
        RECT 121.900 18.075 122.565 18.245 ;
        RECT 121.885 17.525 122.215 17.905 ;
        RECT 122.395 17.695 122.565 18.075 ;
        RECT 122.825 17.525 124.035 18.275 ;
        RECT 128.520 17.740 132.450 18.600 ;
        RECT 92.380 17.355 124.120 17.525 ;
        RECT 92.465 16.605 93.675 17.355 ;
        RECT 93.845 16.810 99.190 17.355 ;
        RECT 99.365 16.810 104.710 17.355 ;
        RECT 104.885 16.810 110.230 17.355 ;
        RECT 110.405 16.810 115.750 17.355 ;
        RECT 92.465 16.065 92.985 16.605 ;
        RECT 93.155 15.895 93.675 16.435 ;
        RECT 95.430 15.980 95.770 16.810 ;
        RECT 92.465 14.805 93.675 15.895 ;
        RECT 97.250 15.240 97.600 16.490 ;
        RECT 100.950 15.980 101.290 16.810 ;
        RECT 102.770 15.240 103.120 16.490 ;
        RECT 106.470 15.980 106.810 16.810 ;
        RECT 108.290 15.240 108.640 16.490 ;
        RECT 111.990 15.980 112.330 16.810 ;
        RECT 115.925 16.705 116.185 17.185 ;
        RECT 116.355 16.815 116.605 17.355 ;
        RECT 113.810 15.240 114.160 16.490 ;
        RECT 115.925 15.675 116.095 16.705 ;
        RECT 116.775 16.650 116.995 17.135 ;
        RECT 116.265 16.055 116.495 16.450 ;
        RECT 116.665 16.225 116.995 16.650 ;
        RECT 117.165 16.975 118.055 17.145 ;
        RECT 117.165 16.250 117.335 16.975 ;
        RECT 117.505 16.420 118.055 16.805 ;
        RECT 118.225 16.630 118.515 17.355 ;
        RECT 119.155 16.955 119.485 17.355 ;
        RECT 119.655 16.785 119.825 17.055 ;
        RECT 119.995 16.955 120.325 17.355 ;
        RECT 120.500 16.795 120.765 17.055 ;
        RECT 121.015 16.865 121.275 17.355 ;
        RECT 120.500 16.785 120.855 16.795 ;
        RECT 117.165 16.180 118.055 16.250 ;
        RECT 117.160 16.155 118.055 16.180 ;
        RECT 117.150 16.140 118.055 16.155 ;
        RECT 117.145 16.125 118.055 16.140 ;
        RECT 117.135 16.120 118.055 16.125 ;
        RECT 117.130 16.110 118.055 16.120 ;
        RECT 117.125 16.100 118.055 16.110 ;
        RECT 117.115 16.095 118.055 16.100 ;
        RECT 117.105 16.085 118.055 16.095 ;
        RECT 117.095 16.080 118.055 16.085 ;
        RECT 117.095 16.075 117.430 16.080 ;
        RECT 117.080 16.070 117.430 16.075 ;
        RECT 117.065 16.060 117.430 16.070 ;
        RECT 117.040 16.055 117.430 16.060 ;
        RECT 116.265 16.050 117.430 16.055 ;
        RECT 116.265 16.015 117.400 16.050 ;
        RECT 116.265 15.990 117.365 16.015 ;
        RECT 116.265 15.960 117.335 15.990 ;
        RECT 116.265 15.930 117.315 15.960 ;
        RECT 116.265 15.900 117.295 15.930 ;
        RECT 116.265 15.890 117.225 15.900 ;
        RECT 116.265 15.880 117.200 15.890 ;
        RECT 116.265 15.865 117.180 15.880 ;
        RECT 116.265 15.850 117.160 15.865 ;
        RECT 116.370 15.840 117.155 15.850 ;
        RECT 116.370 15.805 117.140 15.840 ;
        RECT 93.845 14.805 99.190 15.240 ;
        RECT 99.365 14.805 104.710 15.240 ;
        RECT 104.885 14.805 110.230 15.240 ;
        RECT 110.405 14.805 115.750 15.240 ;
        RECT 115.925 14.975 116.200 15.675 ;
        RECT 116.370 15.555 117.125 15.805 ;
        RECT 117.295 15.485 117.625 15.730 ;
        RECT 117.795 15.630 118.055 16.080 ;
        RECT 117.440 15.460 117.625 15.485 ;
        RECT 117.440 15.360 118.055 15.460 ;
        RECT 116.370 14.805 116.625 15.350 ;
        RECT 116.795 14.975 117.275 15.315 ;
        RECT 117.450 14.805 118.055 15.360 ;
        RECT 118.225 14.805 118.515 15.970 ;
        RECT 119.145 15.775 119.405 16.785 ;
        RECT 119.655 16.615 120.855 16.785 ;
        RECT 119.665 16.195 120.115 16.365 ;
        RECT 119.145 14.805 119.405 15.605 ;
        RECT 119.665 14.990 119.905 16.195 ;
        RECT 120.285 16.025 120.515 16.445 ;
        RECT 120.075 15.825 120.515 16.025 ;
        RECT 120.685 15.945 120.855 16.615 ;
        RECT 121.025 16.115 121.275 16.695 ;
        RECT 121.445 16.680 121.705 17.185 ;
        RECT 121.885 16.975 122.215 17.355 ;
        RECT 122.395 16.805 122.565 17.185 ;
        RECT 120.075 14.990 120.330 15.825 ;
        RECT 120.685 15.775 121.270 15.945 ;
        RECT 120.935 14.990 121.270 15.775 ;
        RECT 121.445 15.880 121.625 16.680 ;
        RECT 121.900 16.635 122.565 16.805 ;
        RECT 121.900 16.380 122.070 16.635 ;
        RECT 122.825 16.605 124.035 17.355 ;
        RECT 121.795 16.050 122.070 16.380 ;
        RECT 122.295 16.085 122.635 16.455 ;
        RECT 121.900 15.905 122.070 16.050 ;
        RECT 121.445 14.975 121.715 15.880 ;
        RECT 121.900 15.735 122.575 15.905 ;
        RECT 121.885 14.805 122.215 15.565 ;
        RECT 122.395 14.975 122.575 15.735 ;
        RECT 122.825 15.895 123.345 16.435 ;
        RECT 123.515 16.065 124.035 16.605 ;
        RECT 128.240 16.140 128.570 16.210 ;
        RECT 128.760 16.140 128.930 17.420 ;
        RECT 129.200 16.380 129.370 17.740 ;
        RECT 128.240 15.940 128.930 16.140 ;
        RECT 122.825 14.805 124.035 15.895 ;
        RECT 128.240 15.870 128.570 15.940 ;
        RECT 128.760 15.310 128.930 15.940 ;
        RECT 129.500 16.140 129.830 16.220 ;
        RECT 130.070 16.140 130.240 17.420 ;
        RECT 130.510 16.380 130.680 17.740 ;
        RECT 129.500 15.940 130.240 16.140 ;
        RECT 129.500 15.880 129.830 15.940 ;
        RECT 129.200 14.980 129.370 15.770 ;
        RECT 130.070 15.310 130.240 15.940 ;
        RECT 130.810 16.140 131.140 16.220 ;
        RECT 131.380 16.140 131.550 17.420 ;
        RECT 131.820 16.380 131.990 17.740 ;
        RECT 132.980 17.150 133.820 20.000 ;
        RECT 139.320 19.560 149.510 19.730 ;
        RECT 141.030 18.950 141.230 19.560 ;
        RECT 151.770 19.250 152.630 20.040 ;
        RECT 141.470 19.080 152.630 19.250 ;
        RECT 141.030 18.620 141.360 18.950 ;
        RECT 141.030 18.120 141.360 18.450 ;
        RECT 151.770 17.950 152.630 19.080 ;
        RECT 141.410 17.780 152.630 17.950 ;
        RECT 141.030 17.300 151.450 17.470 ;
        RECT 132.980 16.980 140.800 17.150 ;
        RECT 130.810 15.940 131.550 16.140 ;
        RECT 130.810 15.880 131.140 15.940 ;
        RECT 130.510 14.980 130.680 15.770 ;
        RECT 131.380 15.310 131.550 15.940 ;
        RECT 132.120 15.880 132.450 16.220 ;
        RECT 131.820 14.980 131.990 15.770 ;
        RECT 92.380 14.635 124.120 14.805 ;
        RECT 92.465 13.545 93.675 14.635 ;
        RECT 93.845 14.200 99.190 14.635 ;
        RECT 99.365 14.200 104.710 14.635 ;
        RECT 92.465 12.835 92.985 13.375 ;
        RECT 93.155 13.005 93.675 13.545 ;
        RECT 92.465 12.085 93.675 12.835 ;
        RECT 95.430 12.630 95.770 13.460 ;
        RECT 97.250 12.950 97.600 14.200 ;
        RECT 100.950 12.630 101.290 13.460 ;
        RECT 102.770 12.950 103.120 14.200 ;
        RECT 105.345 13.470 105.635 14.635 ;
        RECT 105.805 14.200 111.150 14.635 ;
        RECT 93.845 12.085 99.190 12.630 ;
        RECT 99.365 12.085 104.710 12.630 ;
        RECT 105.345 12.085 105.635 12.810 ;
        RECT 107.390 12.630 107.730 13.460 ;
        RECT 109.210 12.950 109.560 14.200 ;
        RECT 111.325 13.545 114.835 14.635 ;
        RECT 111.325 12.855 112.975 13.375 ;
        RECT 113.145 13.025 114.835 13.545 ;
        RECT 115.015 13.495 115.345 14.635 ;
        RECT 115.875 13.665 116.205 14.450 ;
        RECT 115.525 13.495 116.205 13.665 ;
        RECT 116.420 13.845 116.955 14.465 ;
        RECT 115.005 13.075 115.355 13.325 ;
        RECT 115.525 12.895 115.695 13.495 ;
        RECT 115.865 13.075 116.215 13.325 ;
        RECT 105.805 12.085 111.150 12.630 ;
        RECT 111.325 12.085 114.835 12.855 ;
        RECT 115.015 12.085 115.285 12.895 ;
        RECT 115.455 12.255 115.785 12.895 ;
        RECT 115.955 12.085 116.195 12.895 ;
        RECT 116.420 12.825 116.735 13.845 ;
        RECT 117.125 13.835 117.455 14.635 ;
        RECT 118.685 13.915 119.145 14.465 ;
        RECT 119.335 13.915 119.665 14.635 ;
        RECT 117.940 13.665 118.330 13.840 ;
        RECT 116.905 13.495 118.330 13.665 ;
        RECT 116.905 12.995 117.075 13.495 ;
        RECT 116.420 12.255 117.035 12.825 ;
        RECT 117.325 12.765 117.590 13.325 ;
        RECT 117.760 12.595 117.930 13.495 ;
        RECT 118.100 12.765 118.455 13.325 ;
        RECT 117.205 12.085 117.420 12.595 ;
        RECT 117.650 12.265 117.930 12.595 ;
        RECT 118.110 12.085 118.350 12.595 ;
        RECT 118.685 12.545 118.935 13.915 ;
        RECT 119.865 13.745 120.165 14.295 ;
        RECT 120.335 13.965 120.615 14.635 ;
        RECT 119.225 13.575 120.165 13.745 ;
        RECT 119.225 13.325 119.395 13.575 ;
        RECT 120.535 13.325 120.800 13.685 ;
        RECT 119.105 12.995 119.395 13.325 ;
        RECT 119.565 13.075 119.905 13.325 ;
        RECT 120.125 13.075 120.800 13.325 ;
        RECT 121.445 13.560 121.715 14.465 ;
        RECT 121.885 13.875 122.215 14.635 ;
        RECT 122.395 13.705 122.575 14.465 ;
        RECT 119.225 12.905 119.395 12.995 ;
        RECT 119.225 12.715 120.615 12.905 ;
        RECT 118.685 12.255 119.245 12.545 ;
        RECT 119.415 12.085 119.665 12.545 ;
        RECT 120.285 12.355 120.615 12.715 ;
        RECT 121.445 12.760 121.625 13.560 ;
        RECT 121.900 13.535 122.575 13.705 ;
        RECT 122.825 13.545 124.035 14.635 ;
        RECT 128.520 14.140 132.450 14.980 ;
        RECT 121.900 13.390 122.070 13.535 ;
        RECT 121.795 13.060 122.070 13.390 ;
        RECT 121.900 12.805 122.070 13.060 ;
        RECT 122.295 12.985 122.635 13.355 ;
        RECT 122.825 13.005 123.345 13.545 ;
        RECT 123.515 12.835 124.035 13.375 ;
        RECT 121.445 12.255 121.705 12.760 ;
        RECT 121.900 12.635 122.565 12.805 ;
        RECT 121.885 12.085 122.215 12.465 ;
        RECT 122.395 12.255 122.565 12.635 ;
        RECT 122.825 12.085 124.035 12.835 ;
        RECT 128.520 12.820 132.450 13.680 ;
        RECT 92.380 11.915 124.120 12.085 ;
        RECT 92.465 11.165 93.675 11.915 ;
        RECT 93.845 11.370 99.190 11.915 ;
        RECT 99.365 11.370 104.710 11.915 ;
        RECT 104.885 11.370 110.230 11.915 ;
        RECT 110.405 11.370 115.750 11.915 ;
        RECT 92.465 10.625 92.985 11.165 ;
        RECT 93.155 10.455 93.675 10.995 ;
        RECT 95.430 10.540 95.770 11.370 ;
        RECT 92.465 9.365 93.675 10.455 ;
        RECT 97.250 9.800 97.600 11.050 ;
        RECT 100.950 10.540 101.290 11.370 ;
        RECT 102.770 9.800 103.120 11.050 ;
        RECT 106.470 10.540 106.810 11.370 ;
        RECT 108.290 9.800 108.640 11.050 ;
        RECT 111.990 10.540 112.330 11.370 ;
        RECT 115.925 11.145 117.595 11.915 ;
        RECT 118.225 11.190 118.515 11.915 ;
        RECT 118.685 11.145 122.195 11.915 ;
        RECT 122.825 11.165 124.035 11.915 ;
        RECT 113.810 9.800 114.160 11.050 ;
        RECT 115.925 10.625 116.675 11.145 ;
        RECT 116.845 10.455 117.595 10.975 ;
        RECT 118.685 10.625 120.335 11.145 ;
        RECT 93.845 9.365 99.190 9.800 ;
        RECT 99.365 9.365 104.710 9.800 ;
        RECT 104.885 9.365 110.230 9.800 ;
        RECT 110.405 9.365 115.750 9.800 ;
        RECT 115.925 9.365 117.595 10.455 ;
        RECT 118.225 9.365 118.515 10.530 ;
        RECT 120.505 10.455 122.195 10.975 ;
        RECT 118.685 9.365 122.195 10.455 ;
        RECT 122.825 10.455 123.345 10.995 ;
        RECT 123.515 10.625 124.035 11.165 ;
        RECT 128.240 11.220 128.570 11.280 ;
        RECT 128.760 11.220 128.930 12.500 ;
        RECT 129.200 11.460 129.370 12.820 ;
        RECT 128.240 11.020 128.930 11.220 ;
        RECT 128.240 10.940 128.570 11.020 ;
        RECT 122.825 9.365 124.035 10.455 ;
        RECT 128.760 10.390 128.930 11.020 ;
        RECT 129.500 11.220 129.830 11.300 ;
        RECT 130.070 11.220 130.240 12.500 ;
        RECT 130.510 11.460 130.680 12.820 ;
        RECT 129.500 11.020 130.240 11.220 ;
        RECT 129.500 10.960 129.830 11.020 ;
        RECT 129.200 10.070 129.370 10.850 ;
        RECT 130.070 10.390 130.240 11.020 ;
        RECT 130.810 11.220 131.140 11.300 ;
        RECT 131.380 11.220 131.550 12.500 ;
        RECT 131.820 11.460 131.990 12.820 ;
        RECT 132.980 11.610 133.820 16.980 ;
        RECT 141.030 16.710 141.230 17.300 ;
        RECT 151.770 16.990 152.630 17.780 ;
        RECT 141.410 16.820 152.630 16.990 ;
        RECT 139.760 16.540 141.230 16.710 ;
        RECT 141.030 15.950 141.230 16.540 ;
        RECT 151.770 16.430 152.630 16.820 ;
        RECT 141.410 16.260 152.630 16.430 ;
        RECT 141.030 15.780 151.450 15.950 ;
        RECT 141.030 15.130 141.230 15.780 ;
        RECT 151.770 15.470 152.630 16.260 ;
        RECT 141.410 15.300 152.630 15.470 ;
        RECT 141.030 14.800 141.360 15.130 ;
        RECT 141.030 14.300 141.360 14.630 ;
        RECT 151.770 14.130 152.630 15.300 ;
        RECT 141.410 13.960 152.630 14.130 ;
        RECT 141.030 13.480 151.450 13.650 ;
        RECT 141.030 12.690 141.220 13.480 ;
        RECT 151.770 13.170 152.630 13.960 ;
        RECT 141.410 13.000 152.630 13.170 ;
        RECT 141.030 12.520 151.450 12.690 ;
        RECT 141.030 12.130 141.220 12.520 ;
        RECT 141.030 11.960 151.450 12.130 ;
        RECT 141.030 11.940 141.240 11.960 ;
        RECT 132.980 11.440 140.800 11.610 ;
        RECT 130.810 11.020 131.550 11.220 ;
        RECT 130.810 10.960 131.140 11.020 ;
        RECT 130.510 10.070 130.680 10.850 ;
        RECT 131.380 10.390 131.550 11.020 ;
        RECT 132.120 10.960 132.450 11.300 ;
        RECT 131.820 10.070 131.990 10.850 ;
        RECT 92.380 9.195 124.120 9.365 ;
        RECT 128.520 9.220 132.450 10.070 ;
        RECT 92.465 8.105 93.675 9.195 ;
        RECT 93.845 8.760 99.190 9.195 ;
        RECT 99.365 8.760 104.710 9.195 ;
        RECT 92.465 7.395 92.985 7.935 ;
        RECT 93.155 7.565 93.675 8.105 ;
        RECT 92.465 6.645 93.675 7.395 ;
        RECT 95.430 7.190 95.770 8.020 ;
        RECT 97.250 7.510 97.600 8.760 ;
        RECT 100.950 7.190 101.290 8.020 ;
        RECT 102.770 7.510 103.120 8.760 ;
        RECT 105.345 8.030 105.635 9.195 ;
        RECT 105.805 8.760 111.150 9.195 ;
        RECT 111.325 8.760 116.670 9.195 ;
        RECT 93.845 6.645 99.190 7.190 ;
        RECT 99.365 6.645 104.710 7.190 ;
        RECT 105.345 6.645 105.635 7.370 ;
        RECT 107.390 7.190 107.730 8.020 ;
        RECT 109.210 7.510 109.560 8.760 ;
        RECT 112.910 7.190 113.250 8.020 ;
        RECT 114.730 7.510 115.080 8.760 ;
        RECT 116.845 8.105 118.055 9.195 ;
        RECT 116.845 7.395 117.365 7.935 ;
        RECT 117.535 7.565 118.055 8.105 ;
        RECT 118.225 8.030 118.515 9.195 ;
        RECT 118.685 8.105 121.275 9.195 ;
        RECT 118.685 7.415 119.895 7.935 ;
        RECT 120.065 7.585 121.275 8.105 ;
        RECT 121.445 8.120 121.715 9.025 ;
        RECT 121.885 8.435 122.215 9.195 ;
        RECT 122.395 8.265 122.575 9.025 ;
        RECT 105.805 6.645 111.150 7.190 ;
        RECT 111.325 6.645 116.670 7.190 ;
        RECT 116.845 6.645 118.055 7.395 ;
        RECT 118.225 6.645 118.515 7.370 ;
        RECT 118.685 6.645 121.275 7.415 ;
        RECT 121.445 7.320 121.625 8.120 ;
        RECT 121.900 8.095 122.575 8.265 ;
        RECT 122.825 8.105 124.035 9.195 ;
        RECT 121.900 7.950 122.070 8.095 ;
        RECT 121.795 7.620 122.070 7.950 ;
        RECT 121.900 7.365 122.070 7.620 ;
        RECT 122.295 7.545 122.635 7.915 ;
        RECT 122.825 7.565 123.345 8.105 ;
        RECT 123.515 7.395 124.035 7.935 ;
        RECT 128.520 7.900 132.450 8.760 ;
        RECT 132.980 8.010 133.820 11.440 ;
        RECT 141.040 11.170 141.240 11.940 ;
        RECT 151.770 11.650 152.630 13.000 ;
        RECT 141.410 11.480 152.630 11.650 ;
        RECT 140.290 11.000 151.450 11.170 ;
        RECT 141.040 10.130 141.240 11.000 ;
        RECT 151.770 10.690 152.630 11.480 ;
        RECT 141.410 10.520 152.630 10.690 ;
        RECT 141.040 9.960 151.450 10.130 ;
        RECT 141.040 9.170 141.240 9.960 ;
        RECT 151.770 9.650 152.630 10.520 ;
        RECT 141.410 9.480 152.630 9.650 ;
        RECT 141.040 9.000 151.450 9.170 ;
        RECT 141.040 8.350 141.240 9.000 ;
        RECT 151.770 8.690 152.630 9.480 ;
        RECT 141.410 8.520 152.630 8.690 ;
        RECT 141.040 8.020 141.370 8.350 ;
        RECT 151.770 8.020 152.630 8.520 ;
        RECT 121.445 6.815 121.705 7.320 ;
        RECT 121.900 7.195 122.565 7.365 ;
        RECT 121.885 6.645 122.215 7.025 ;
        RECT 122.395 6.815 122.565 7.195 ;
        RECT 122.825 6.645 124.035 7.395 ;
        RECT 92.380 6.475 124.120 6.645 ;
        RECT 128.240 6.300 128.570 6.360 ;
        RECT 128.760 6.300 128.930 7.580 ;
        RECT 129.200 6.540 129.370 7.900 ;
        RECT 128.240 6.100 128.930 6.300 ;
        RECT 128.240 6.020 128.570 6.100 ;
        RECT 128.760 5.470 128.930 6.100 ;
        RECT 129.500 6.300 129.830 6.380 ;
        RECT 130.070 6.300 130.240 7.580 ;
        RECT 130.510 6.540 130.680 7.900 ;
        RECT 129.500 6.100 130.240 6.300 ;
        RECT 129.500 6.040 129.830 6.100 ;
        RECT 129.200 5.140 129.370 5.930 ;
        RECT 130.070 5.470 130.240 6.100 ;
        RECT 130.810 6.300 131.140 6.380 ;
        RECT 131.380 6.300 131.550 7.580 ;
        RECT 131.820 6.540 131.990 7.900 ;
        RECT 130.810 6.100 131.550 6.300 ;
        RECT 130.810 6.040 131.140 6.100 ;
        RECT 130.510 5.140 130.680 5.930 ;
        RECT 131.380 5.470 131.550 6.100 ;
        RECT 132.120 6.040 132.450 6.380 ;
        RECT 131.820 5.140 131.990 5.930 ;
        RECT 128.520 4.300 132.450 5.140 ;
      LAYER met1 ;
        RECT 126.550 38.310 152.610 38.320 ;
        RECT 126.550 38.290 152.630 38.310 ;
        RECT 107.900 37.420 152.630 38.290 ;
        RECT 126.550 37.410 152.630 37.420 ;
        RECT 92.380 36.240 124.120 36.720 ;
        RECT 120.970 34.820 121.290 35.080 ;
        RECT 122.350 34.820 122.670 35.080 ;
        RECT 120.050 34.140 120.370 34.400 ;
        RECT 121.445 34.340 121.735 34.385 ;
        RECT 122.810 34.340 123.130 34.400 ;
        RECT 121.445 34.200 123.130 34.340 ;
        RECT 121.445 34.155 121.735 34.200 ;
        RECT 122.810 34.140 123.130 34.200 ;
        RECT 92.380 33.520 124.120 34.000 ;
        RECT 127.200 33.380 127.950 37.410 ;
        RECT 128.730 36.090 128.960 37.090 ;
        RECT 129.170 36.090 129.400 37.090 ;
        RECT 130.040 36.090 130.270 37.090 ;
        RECT 130.480 36.090 130.710 37.090 ;
        RECT 131.350 36.090 131.580 37.090 ;
        RECT 131.790 36.090 132.020 37.090 ;
        RECT 128.240 35.560 128.570 35.900 ;
        RECT 132.120 35.570 132.450 35.910 ;
        RECT 128.730 35.020 128.960 35.440 ;
        RECT 129.170 35.020 129.400 35.440 ;
        RECT 130.040 35.020 130.270 35.440 ;
        RECT 130.480 35.020 130.710 35.440 ;
        RECT 131.350 35.020 131.580 35.440 ;
        RECT 131.790 35.020 132.020 35.440 ;
        RECT 132.450 34.670 133.910 34.680 ;
        RECT 128.520 33.840 133.910 34.670 ;
        RECT 128.520 33.830 132.450 33.840 ;
        RECT 132.900 33.630 133.910 33.840 ;
        RECT 127.200 33.370 132.440 33.380 ;
        RECT 127.200 32.520 132.450 33.370 ;
        RECT 92.380 30.800 124.120 31.280 ;
        RECT 122.350 29.380 122.670 29.640 ;
        RECT 121.430 28.700 121.750 28.960 ;
        RECT 92.380 28.080 124.120 28.560 ;
        RECT 127.200 28.440 127.950 32.520 ;
        RECT 128.520 32.510 132.450 32.520 ;
        RECT 128.730 31.170 128.960 32.170 ;
        RECT 129.170 31.170 129.400 32.170 ;
        RECT 130.040 31.170 130.270 32.170 ;
        RECT 130.480 31.170 130.710 32.170 ;
        RECT 131.350 31.170 131.580 32.170 ;
        RECT 131.790 31.170 132.020 32.170 ;
        RECT 128.240 30.620 128.570 30.960 ;
        RECT 132.120 30.650 132.450 30.990 ;
        RECT 128.730 30.100 128.960 30.520 ;
        RECT 129.170 30.100 129.400 30.520 ;
        RECT 130.040 30.100 130.270 30.520 ;
        RECT 130.480 30.100 130.710 30.520 ;
        RECT 131.350 30.100 131.580 30.520 ;
        RECT 131.790 30.100 132.020 30.520 ;
        RECT 132.980 29.750 133.820 33.630 ;
        RECT 134.170 33.190 140.840 33.420 ;
        RECT 141.030 33.120 141.360 33.450 ;
        RECT 134.170 32.710 140.840 32.940 ;
        RECT 134.170 32.230 140.840 32.460 ;
        RECT 134.170 31.670 140.840 31.900 ;
        RECT 141.490 31.630 141.960 31.860 ;
        RECT 134.170 31.190 140.840 31.420 ;
        RECT 141.490 31.190 141.960 31.420 ;
        RECT 134.170 30.710 140.840 30.940 ;
        RECT 134.170 30.150 140.840 30.380 ;
        RECT 128.520 28.910 133.820 29.750 ;
        RECT 134.170 29.670 140.840 29.900 ;
        RECT 134.170 29.190 140.840 29.420 ;
        RECT 141.030 29.160 141.360 29.490 ;
        RECT 119.130 27.880 119.450 27.940 ;
        RECT 120.050 27.880 120.370 27.940 ;
        RECT 120.525 27.880 120.815 27.925 ;
        RECT 116.000 27.740 120.815 27.880 ;
        RECT 116.000 27.585 116.140 27.740 ;
        RECT 119.130 27.680 119.450 27.740 ;
        RECT 120.050 27.680 120.370 27.740 ;
        RECT 120.525 27.695 120.815 27.740 ;
        RECT 115.925 27.355 116.215 27.585 ;
        RECT 117.005 27.540 117.295 27.585 ;
        RECT 121.905 27.540 122.195 27.585 ;
        RECT 117.005 27.400 120.280 27.540 ;
        RECT 117.005 27.355 117.295 27.400 ;
        RECT 119.605 27.015 119.895 27.245 ;
        RECT 117.765 26.520 118.055 26.565 ;
        RECT 119.680 26.520 119.820 27.015 ;
        RECT 120.140 26.920 120.280 27.400 ;
        RECT 121.060 27.400 122.195 27.540 ;
        RECT 121.060 27.245 121.200 27.400 ;
        RECT 121.905 27.355 122.195 27.400 ;
        RECT 127.200 27.580 132.450 28.440 ;
        RECT 120.985 27.015 121.275 27.245 ;
        RECT 121.430 27.000 121.750 27.260 ;
        RECT 122.365 27.200 122.655 27.245 ;
        RECT 122.810 27.200 123.130 27.260 ;
        RECT 122.365 27.060 123.130 27.200 ;
        RECT 122.365 27.015 122.655 27.060 ;
        RECT 122.810 27.000 123.130 27.060 ;
        RECT 120.050 26.860 120.370 26.920 ;
        RECT 121.520 26.860 121.660 27.000 ;
        RECT 120.050 26.720 121.660 26.860 ;
        RECT 120.050 26.660 120.370 26.720 ;
        RECT 117.765 26.380 119.820 26.520 ;
        RECT 117.765 26.335 118.055 26.380 ;
        RECT 116.845 26.180 117.135 26.225 ;
        RECT 117.290 26.180 117.610 26.240 ;
        RECT 116.845 26.040 117.610 26.180 ;
        RECT 116.845 25.995 117.135 26.040 ;
        RECT 117.290 25.980 117.610 26.040 ;
        RECT 118.670 25.980 118.990 26.240 ;
        RECT 92.380 25.360 124.120 25.840 ;
        RECT 103.490 24.820 103.810 24.880 ;
        RECT 114.545 24.820 114.835 24.865 ;
        RECT 103.490 24.680 114.835 24.820 ;
        RECT 103.490 24.620 103.810 24.680 ;
        RECT 114.545 24.635 114.835 24.680 ;
        RECT 119.130 23.940 119.450 24.200 ;
        RECT 120.510 23.940 120.830 24.200 ;
        RECT 122.350 23.940 122.670 24.200 ;
        RECT 114.990 23.800 115.310 23.860 ;
        RECT 116.845 23.800 117.135 23.845 ;
        RECT 114.990 23.660 117.135 23.800 ;
        RECT 114.990 23.600 115.310 23.660 ;
        RECT 116.845 23.615 117.135 23.660 ;
        RECT 117.290 23.800 117.610 23.860 ;
        RECT 118.685 23.800 118.975 23.845 ;
        RECT 120.970 23.800 121.290 23.860 ;
        RECT 122.810 23.800 123.130 23.860 ;
        RECT 117.290 23.660 123.130 23.800 ;
        RECT 117.290 23.600 117.610 23.660 ;
        RECT 118.685 23.615 118.975 23.660 ;
        RECT 120.970 23.600 121.290 23.660 ;
        RECT 122.810 23.600 123.130 23.660 ;
        RECT 127.200 23.520 127.950 27.580 ;
        RECT 128.730 26.240 128.960 27.240 ;
        RECT 129.170 26.240 129.400 27.240 ;
        RECT 130.040 26.240 130.270 27.240 ;
        RECT 130.480 26.240 130.710 27.240 ;
        RECT 131.350 26.240 131.580 27.240 ;
        RECT 131.790 26.240 132.020 27.240 ;
        RECT 128.240 25.710 128.570 26.050 ;
        RECT 132.120 25.720 132.450 26.060 ;
        RECT 128.730 25.170 128.960 25.590 ;
        RECT 129.170 25.170 129.400 25.590 ;
        RECT 130.040 25.170 130.270 25.590 ;
        RECT 130.480 25.170 130.710 25.590 ;
        RECT 131.350 25.170 131.580 25.590 ;
        RECT 131.790 25.170 132.020 25.590 ;
        RECT 132.980 24.830 133.820 28.910 ;
        RECT 136.340 28.630 140.840 28.860 ;
        RECT 141.030 28.560 141.360 28.890 ;
        RECT 136.340 28.150 140.840 28.380 ;
        RECT 136.340 27.670 140.840 27.900 ;
        RECT 141.860 27.830 143.860 28.060 ;
        RECT 141.860 27.390 143.860 27.620 ;
        RECT 136.340 27.110 140.840 27.340 ;
        RECT 136.340 26.630 140.840 26.860 ;
        RECT 136.340 26.150 140.840 26.380 ;
        RECT 141.030 26.120 141.360 26.450 ;
        RECT 138.340 25.590 140.840 25.820 ;
        RECT 141.030 25.520 141.360 25.850 ;
        RECT 138.340 25.110 140.840 25.340 ;
        RECT 128.510 23.990 133.820 24.830 ;
        RECT 138.340 24.630 140.840 24.860 ;
        RECT 141.490 24.790 148.490 25.020 ;
        RECT 141.490 24.350 148.490 24.580 ;
        RECT 138.340 24.070 140.840 24.300 ;
        RECT 128.510 23.980 132.460 23.990 ;
        RECT 121.430 23.260 121.750 23.520 ;
        RECT 92.380 22.640 124.120 23.120 ;
        RECT 127.200 22.660 132.450 23.520 ;
        RECT 119.590 22.440 119.910 22.500 ;
        RECT 120.065 22.440 120.355 22.485 ;
        RECT 121.430 22.440 121.750 22.500 ;
        RECT 119.590 22.300 121.750 22.440 ;
        RECT 119.590 22.240 119.910 22.300 ;
        RECT 120.065 22.255 120.355 22.300 ;
        RECT 121.430 22.240 121.750 22.300 ;
        RECT 110.390 22.100 110.710 22.160 ;
        RECT 114.085 22.100 114.375 22.145 ;
        RECT 110.390 21.960 114.375 22.100 ;
        RECT 110.390 21.900 110.710 21.960 ;
        RECT 114.085 21.915 114.375 21.960 ;
        RECT 115.925 22.100 116.215 22.145 ;
        RECT 116.830 22.100 117.150 22.160 ;
        RECT 119.145 22.100 119.435 22.145 ;
        RECT 115.925 21.960 119.435 22.100 ;
        RECT 115.925 21.915 116.215 21.960 ;
        RECT 116.830 21.900 117.150 21.960 ;
        RECT 119.145 21.915 119.435 21.960 ;
        RECT 120.970 21.900 121.290 22.160 ;
        RECT 114.990 21.560 115.310 21.820 ;
        RECT 116.385 21.575 116.675 21.805 ;
        RECT 120.050 21.760 120.370 21.820 ;
        RECT 120.525 21.760 120.815 21.805 ;
        RECT 120.050 21.620 120.815 21.760 ;
        RECT 115.910 21.420 116.230 21.480 ;
        RECT 116.460 21.420 116.600 21.575 ;
        RECT 120.050 21.560 120.370 21.620 ;
        RECT 120.525 21.575 120.815 21.620 ;
        RECT 115.910 21.280 116.600 21.420 ;
        RECT 119.130 21.420 119.450 21.480 ;
        RECT 121.905 21.420 122.195 21.465 ;
        RECT 119.130 21.280 122.195 21.420 ;
        RECT 115.910 21.220 116.230 21.280 ;
        RECT 119.130 21.220 119.450 21.280 ;
        RECT 121.905 21.235 122.195 21.280 ;
        RECT 92.380 19.920 124.120 20.400 ;
        RECT 120.510 19.720 120.830 19.780 ;
        RECT 121.445 19.720 121.735 19.765 ;
        RECT 120.510 19.580 121.735 19.720 ;
        RECT 120.510 19.520 120.830 19.580 ;
        RECT 121.445 19.535 121.735 19.580 ;
        RECT 118.670 19.040 118.990 19.100 ;
        RECT 119.145 19.040 119.435 19.085 ;
        RECT 118.670 18.900 119.435 19.040 ;
        RECT 118.670 18.840 118.990 18.900 ;
        RECT 119.145 18.855 119.435 18.900 ;
        RECT 116.370 18.500 116.690 18.760 ;
        RECT 116.830 18.500 117.150 18.760 ;
        RECT 117.750 18.500 118.070 18.760 ;
        RECT 120.510 18.700 120.830 18.760 ;
        RECT 122.365 18.700 122.655 18.745 ;
        RECT 120.510 18.560 122.655 18.700 ;
        RECT 120.510 18.500 120.830 18.560 ;
        RECT 122.365 18.515 122.655 18.560 ;
        RECT 127.200 18.600 127.950 22.660 ;
        RECT 128.730 21.320 128.960 22.320 ;
        RECT 129.170 21.320 129.400 22.320 ;
        RECT 130.040 21.320 130.270 22.320 ;
        RECT 130.480 21.320 130.710 22.320 ;
        RECT 131.350 21.320 131.580 22.320 ;
        RECT 131.790 21.320 132.020 22.320 ;
        RECT 128.240 20.790 128.570 21.130 ;
        RECT 132.120 20.800 132.450 21.140 ;
        RECT 128.730 20.250 128.960 20.670 ;
        RECT 129.170 20.250 129.400 20.670 ;
        RECT 130.040 20.250 130.270 20.670 ;
        RECT 130.480 20.250 130.710 20.670 ;
        RECT 131.350 20.250 131.580 20.670 ;
        RECT 131.790 20.250 132.020 20.670 ;
        RECT 132.980 19.900 133.820 23.990 ;
        RECT 138.340 23.590 140.840 23.820 ;
        RECT 138.340 23.110 140.840 23.340 ;
        RECT 141.030 23.080 141.360 23.410 ;
        RECT 141.030 22.580 141.360 22.910 ;
        RECT 138.340 22.250 140.840 22.480 ;
        RECT 141.490 22.250 148.990 22.480 ;
        RECT 138.340 21.770 140.840 22.000 ;
        RECT 141.490 21.770 148.990 22.000 ;
        RECT 138.340 21.290 140.840 21.520 ;
        RECT 141.490 21.290 148.990 21.520 ;
        RECT 141.030 20.840 141.360 21.170 ;
        RECT 141.030 20.340 141.360 20.670 ;
        RECT 139.340 19.970 140.840 20.200 ;
        RECT 141.490 20.010 149.490 20.240 ;
        RECT 128.520 19.060 133.820 19.900 ;
        RECT 139.340 19.530 140.840 19.760 ;
        RECT 141.490 19.530 149.490 19.760 ;
        RECT 128.520 19.050 132.450 19.060 ;
        RECT 113.610 18.160 113.930 18.420 ;
        RECT 127.200 17.740 132.450 18.600 ;
        RECT 92.380 17.200 124.120 17.680 ;
        RECT 114.990 17.000 115.310 17.060 ;
        RECT 116.830 17.045 117.150 17.060 ;
        RECT 115.925 17.000 116.215 17.045 ;
        RECT 114.990 16.860 116.215 17.000 ;
        RECT 114.990 16.800 115.310 16.860 ;
        RECT 115.925 16.815 116.215 16.860 ;
        RECT 116.765 16.815 117.150 17.045 ;
        RECT 116.830 16.800 117.150 16.815 ;
        RECT 120.510 16.800 120.830 17.060 ;
        RECT 117.750 16.660 118.070 16.720 ;
        RECT 117.750 16.520 120.280 16.660 ;
        RECT 117.750 16.460 118.070 16.520 ;
        RECT 119.590 16.120 119.910 16.380 ;
        RECT 120.140 16.025 120.280 16.520 ;
        RECT 120.985 16.320 121.275 16.365 ;
        RECT 121.430 16.320 121.750 16.380 ;
        RECT 120.985 16.180 121.750 16.320 ;
        RECT 120.985 16.135 121.275 16.180 ;
        RECT 121.430 16.120 121.750 16.180 ;
        RECT 122.350 16.120 122.670 16.380 ;
        RECT 119.145 15.795 119.435 16.025 ;
        RECT 120.065 15.980 120.355 16.025 ;
        RECT 120.065 15.840 121.660 15.980 ;
        RECT 120.065 15.795 120.355 15.840 ;
        RECT 119.220 15.640 119.360 15.795 ;
        RECT 120.510 15.640 120.830 15.700 ;
        RECT 121.520 15.685 121.660 15.840 ;
        RECT 119.220 15.500 120.830 15.640 ;
        RECT 120.510 15.440 120.830 15.500 ;
        RECT 121.445 15.455 121.735 15.685 ;
        RECT 116.845 15.300 117.135 15.345 ;
        RECT 120.970 15.300 121.290 15.360 ;
        RECT 116.845 15.160 121.290 15.300 ;
        RECT 116.845 15.115 117.135 15.160 ;
        RECT 120.970 15.100 121.290 15.160 ;
        RECT 92.380 14.480 124.120 14.960 ;
        RECT 115.910 14.080 116.230 14.340 ;
        RECT 116.370 14.080 116.690 14.340 ;
        RECT 121.430 14.080 121.750 14.340 ;
        RECT 116.000 13.600 116.140 14.080 ;
        RECT 121.520 13.600 121.660 14.080 ;
        RECT 116.000 13.460 117.520 13.600 ;
        RECT 117.380 13.305 117.520 13.460 ;
        RECT 119.680 13.460 121.660 13.600 ;
        RECT 127.200 13.680 127.950 17.740 ;
        RECT 128.730 16.400 128.960 17.400 ;
        RECT 129.170 16.400 129.400 17.400 ;
        RECT 130.040 16.400 130.270 17.400 ;
        RECT 130.480 16.400 130.710 17.400 ;
        RECT 131.350 16.400 131.580 17.400 ;
        RECT 131.790 16.400 132.020 17.400 ;
        RECT 128.240 15.870 128.570 16.210 ;
        RECT 132.120 15.880 132.450 16.220 ;
        RECT 128.730 15.330 128.960 15.750 ;
        RECT 129.170 15.330 129.400 15.750 ;
        RECT 130.040 15.330 130.270 15.750 ;
        RECT 130.480 15.330 130.710 15.750 ;
        RECT 131.350 15.330 131.580 15.750 ;
        RECT 131.790 15.330 132.020 15.750 ;
        RECT 132.980 14.990 133.820 19.060 ;
        RECT 141.490 19.050 149.490 19.280 ;
        RECT 141.030 18.620 141.360 18.950 ;
        RECT 141.030 18.120 141.360 18.450 ;
        RECT 141.430 17.750 151.430 17.980 ;
        RECT 141.430 17.270 151.430 17.500 ;
        RECT 139.780 16.950 140.780 17.180 ;
        RECT 141.430 16.790 151.430 17.020 ;
        RECT 139.780 16.510 140.780 16.740 ;
        RECT 141.430 16.230 151.430 16.460 ;
        RECT 141.430 15.750 151.430 15.980 ;
        RECT 141.430 15.270 151.430 15.500 ;
        RECT 132.450 14.980 133.820 14.990 ;
        RECT 128.520 14.150 133.820 14.980 ;
        RECT 141.030 14.800 141.360 15.130 ;
        RECT 141.030 14.300 141.360 14.630 ;
        RECT 128.520 14.140 132.450 14.150 ;
        RECT 119.680 13.305 119.820 13.460 ;
        RECT 115.005 13.075 115.295 13.305 ;
        RECT 115.925 13.075 116.215 13.305 ;
        RECT 117.305 13.075 117.595 13.305 ;
        RECT 119.605 13.260 119.895 13.305 ;
        RECT 117.840 13.120 119.895 13.260 ;
        RECT 115.080 12.580 115.220 13.075 ;
        RECT 116.000 12.920 116.140 13.075 ;
        RECT 117.840 12.920 117.980 13.120 ;
        RECT 119.605 13.075 119.895 13.120 ;
        RECT 120.510 13.260 120.830 13.320 ;
        RECT 121.430 13.260 121.750 13.320 ;
        RECT 120.510 13.120 121.750 13.260 ;
        RECT 120.510 13.060 120.830 13.120 ;
        RECT 121.430 13.060 121.750 13.120 ;
        RECT 122.350 13.060 122.670 13.320 ;
        RECT 116.000 12.780 117.980 12.920 ;
        RECT 118.225 12.920 118.515 12.965 ;
        RECT 118.685 12.920 118.975 12.965 ;
        RECT 118.225 12.780 118.975 12.920 ;
        RECT 118.225 12.735 118.515 12.780 ;
        RECT 118.685 12.735 118.975 12.780 ;
        RECT 120.600 12.580 120.740 13.060 ;
        RECT 115.080 12.440 120.740 12.580 ;
        RECT 127.200 12.820 132.450 13.680 ;
        RECT 92.380 11.760 124.120 12.240 ;
        RECT 92.380 9.040 124.120 9.520 ;
        RECT 121.430 8.640 121.750 8.900 ;
        RECT 127.200 8.760 127.950 12.820 ;
        RECT 128.730 11.480 128.960 12.480 ;
        RECT 129.170 11.480 129.400 12.480 ;
        RECT 130.040 11.480 130.270 12.480 ;
        RECT 130.480 11.480 130.710 12.480 ;
        RECT 131.350 11.480 131.580 12.480 ;
        RECT 131.790 11.480 132.020 12.480 ;
        RECT 128.240 10.940 128.570 11.280 ;
        RECT 132.120 10.960 132.450 11.300 ;
        RECT 128.730 10.410 128.960 10.830 ;
        RECT 129.170 10.410 129.400 10.830 ;
        RECT 130.040 10.410 130.270 10.830 ;
        RECT 130.480 10.410 130.710 10.830 ;
        RECT 131.350 10.410 131.580 10.830 ;
        RECT 131.790 10.410 132.020 10.830 ;
        RECT 132.980 10.070 133.820 14.150 ;
        RECT 141.430 13.930 151.430 14.160 ;
        RECT 141.430 13.450 151.430 13.680 ;
        RECT 141.430 12.970 151.430 13.200 ;
        RECT 141.430 12.490 151.430 12.720 ;
        RECT 141.430 11.930 151.430 12.160 ;
        RECT 140.310 11.410 140.780 11.640 ;
        RECT 141.430 11.450 151.430 11.680 ;
        RECT 140.310 10.970 140.780 11.200 ;
        RECT 141.430 10.970 151.430 11.200 ;
        RECT 141.430 10.490 151.430 10.720 ;
        RECT 128.520 9.230 133.820 10.070 ;
        RECT 141.430 9.930 151.430 10.160 ;
        RECT 141.430 9.450 151.430 9.680 ;
        RECT 128.520 9.220 132.450 9.230 ;
        RECT 127.200 7.900 132.450 8.760 ;
        RECT 122.350 7.620 122.670 7.880 ;
        RECT 92.380 6.320 124.120 6.800 ;
        RECT 128.730 6.560 128.960 7.560 ;
        RECT 129.170 6.560 129.400 7.560 ;
        RECT 130.040 6.560 130.270 7.560 ;
        RECT 130.480 6.560 130.710 7.560 ;
        RECT 131.350 6.560 131.580 7.560 ;
        RECT 131.790 6.560 132.020 7.560 ;
        RECT 128.240 6.020 128.570 6.360 ;
        RECT 132.120 6.040 132.450 6.380 ;
        RECT 128.730 5.490 128.960 5.910 ;
        RECT 129.170 5.490 129.400 5.910 ;
        RECT 130.040 5.490 130.270 5.910 ;
        RECT 130.480 5.490 130.710 5.910 ;
        RECT 131.350 5.490 131.580 5.910 ;
        RECT 131.790 5.490 132.020 5.910 ;
        RECT 132.980 5.140 133.820 9.230 ;
        RECT 141.430 8.970 151.430 9.200 ;
        RECT 141.430 8.490 151.430 8.720 ;
        RECT 141.040 8.020 141.370 8.350 ;
        RECT 151.770 8.020 152.630 37.410 ;
        RECT 111.200 4.300 133.820 5.140 ;
      LAYER met2 ;
        RECT 107.900 37.420 109.500 38.290 ;
        RECT 107.930 36.295 109.470 36.665 ;
        RECT 120.990 36.635 121.270 37.005 ;
        RECT 121.060 35.110 121.200 36.635 ;
        RECT 125.900 35.900 126.240 38.360 ;
        RECT 125.900 35.560 128.570 35.900 ;
        RECT 132.120 35.570 140.820 35.910 ;
        RECT 121.000 34.790 121.260 35.110 ;
        RECT 122.380 34.790 122.640 35.110 ;
        RECT 110.410 33.915 110.690 34.285 ;
        RECT 120.080 34.110 120.340 34.430 ;
        RECT 122.440 34.285 122.580 34.790 ;
        RECT 107.930 30.855 109.470 31.225 ;
        RECT 107.930 25.415 109.470 25.785 ;
        RECT 103.520 24.590 103.780 24.910 ;
        RECT 103.580 22.045 103.720 24.590 ;
        RECT 110.480 22.190 110.620 33.915 ;
        RECT 111.230 33.575 112.770 33.945 ;
        RECT 111.230 28.135 112.770 28.505 ;
        RECT 120.140 27.970 120.280 34.110 ;
        RECT 122.370 33.915 122.650 34.285 ;
        RECT 122.840 34.110 123.100 34.430 ;
        RECT 122.380 29.350 122.640 29.670 ;
        RECT 121.460 28.670 121.720 28.990 ;
        RECT 122.440 28.845 122.580 29.350 ;
        RECT 119.160 27.650 119.420 27.970 ;
        RECT 120.080 27.650 120.340 27.970 ;
        RECT 117.320 25.950 117.580 26.270 ;
        RECT 118.700 25.950 118.960 26.270 ;
        RECT 117.380 23.890 117.520 25.950 ;
        RECT 115.020 23.570 115.280 23.890 ;
        RECT 117.320 23.570 117.580 23.890 ;
        RECT 111.230 22.695 112.770 23.065 ;
        RECT 103.510 21.675 103.790 22.045 ;
        RECT 110.420 21.870 110.680 22.190 ;
        RECT 115.080 21.850 115.220 23.570 ;
        RECT 116.860 21.870 117.120 22.190 ;
        RECT 115.020 21.530 115.280 21.850 ;
        RECT 107.930 19.975 109.470 20.345 ;
        RECT 113.640 18.130 113.900 18.450 ;
        RECT 111.230 17.255 112.770 17.625 ;
        RECT 107.930 14.535 109.470 14.905 ;
        RECT 111.230 11.815 112.770 12.185 ;
        RECT 113.700 10.485 113.840 18.130 ;
        RECT 115.080 17.090 115.220 21.530 ;
        RECT 115.940 21.190 116.200 21.510 ;
        RECT 115.020 16.770 115.280 17.090 ;
        RECT 116.000 14.370 116.140 21.190 ;
        RECT 116.920 18.790 117.060 21.870 ;
        RECT 118.760 19.130 118.900 25.950 ;
        RECT 119.220 24.230 119.360 27.650 ;
        RECT 121.520 27.290 121.660 28.670 ;
        RECT 122.370 28.475 122.650 28.845 ;
        RECT 122.900 27.290 123.040 34.110 ;
        RECT 126.010 30.960 126.350 32.930 ;
        RECT 126.010 30.620 128.570 30.960 ;
        RECT 132.120 30.650 140.350 30.990 ;
        RECT 121.460 26.970 121.720 27.290 ;
        RECT 122.840 26.970 123.100 27.290 ;
        RECT 120.080 26.630 120.340 26.950 ;
        RECT 119.160 23.910 119.420 24.230 ;
        RECT 119.220 21.510 119.360 23.910 ;
        RECT 119.620 22.210 119.880 22.530 ;
        RECT 119.160 21.190 119.420 21.510 ;
        RECT 118.700 18.810 118.960 19.130 ;
        RECT 116.400 18.470 116.660 18.790 ;
        RECT 116.860 18.470 117.120 18.790 ;
        RECT 117.780 18.470 118.040 18.790 ;
        RECT 116.460 14.370 116.600 18.470 ;
        RECT 116.920 17.090 117.060 18.470 ;
        RECT 116.860 16.770 117.120 17.090 ;
        RECT 117.840 16.750 117.980 18.470 ;
        RECT 117.780 16.430 118.040 16.750 ;
        RECT 119.680 16.410 119.820 22.210 ;
        RECT 120.140 21.850 120.280 26.630 ;
        RECT 120.540 23.910 120.800 24.230 ;
        RECT 122.380 23.910 122.640 24.230 ;
        RECT 120.080 21.530 120.340 21.850 ;
        RECT 120.600 19.810 120.740 23.910 ;
        RECT 121.000 23.570 121.260 23.890 ;
        RECT 121.060 22.190 121.200 23.570 ;
        RECT 121.460 23.230 121.720 23.550 ;
        RECT 122.440 23.405 122.580 23.910 ;
        RECT 122.900 23.890 123.040 26.970 ;
        RECT 126.010 26.050 126.350 27.490 ;
        RECT 140.020 26.450 140.350 30.650 ;
        RECT 140.490 29.490 140.820 35.570 ;
        RECT 141.030 33.370 141.360 33.450 ;
        RECT 141.030 33.200 141.680 33.370 ;
        RECT 141.030 33.120 141.360 33.200 ;
        RECT 140.490 29.160 141.360 29.490 ;
        RECT 141.030 28.810 141.360 28.890 ;
        RECT 141.510 28.810 141.680 33.200 ;
        RECT 141.030 28.640 141.680 28.810 ;
        RECT 141.030 28.560 141.360 28.640 ;
        RECT 140.020 26.120 141.360 26.450 ;
        RECT 126.010 25.710 128.570 26.050 ;
        RECT 132.120 25.720 139.880 26.060 ;
        RECT 122.840 23.570 123.100 23.890 ;
        RECT 139.550 23.410 139.880 25.720 ;
        RECT 141.030 25.770 141.360 25.850 ;
        RECT 141.510 25.770 141.680 28.640 ;
        RECT 141.030 25.600 141.680 25.770 ;
        RECT 141.030 25.520 141.360 25.600 ;
        RECT 121.520 22.530 121.660 23.230 ;
        RECT 122.370 23.035 122.650 23.405 ;
        RECT 139.550 23.080 141.360 23.410 ;
        RECT 141.030 22.830 141.360 22.910 ;
        RECT 141.510 22.830 141.680 25.600 ;
        RECT 141.030 22.660 141.680 22.830 ;
        RECT 141.030 22.580 141.360 22.660 ;
        RECT 121.460 22.210 121.720 22.530 ;
        RECT 121.000 21.870 121.260 22.190 ;
        RECT 126.010 21.130 126.350 22.060 ;
        RECT 126.010 20.790 128.570 21.130 ;
        RECT 132.120 20.840 141.360 21.170 ;
        RECT 132.120 20.800 132.450 20.840 ;
        RECT 141.030 20.590 141.360 20.670 ;
        RECT 141.510 20.590 141.680 22.660 ;
        RECT 141.030 20.420 141.680 20.590 ;
        RECT 141.030 20.340 141.360 20.420 ;
        RECT 120.540 19.490 120.800 19.810 ;
        RECT 120.540 18.470 120.800 18.790 ;
        RECT 140.490 18.620 141.360 18.950 ;
        RECT 120.600 17.090 120.740 18.470 ;
        RECT 120.540 16.770 120.800 17.090 ;
        RECT 119.620 16.090 119.880 16.410 ;
        RECT 121.460 16.090 121.720 16.410 ;
        RECT 122.370 16.235 122.650 16.605 ;
        RECT 122.380 16.090 122.640 16.235 ;
        RECT 126.010 16.210 126.350 16.580 ;
        RECT 140.490 16.220 140.820 18.620 ;
        RECT 141.030 18.370 141.360 18.450 ;
        RECT 141.510 18.370 141.680 20.420 ;
        RECT 141.030 18.200 141.680 18.370 ;
        RECT 141.030 18.120 141.360 18.200 ;
        RECT 120.540 15.410 120.800 15.730 ;
        RECT 115.940 14.050 116.200 14.370 ;
        RECT 116.400 14.050 116.660 14.370 ;
        RECT 120.600 13.350 120.740 15.410 ;
        RECT 121.000 15.130 121.260 15.390 ;
        RECT 121.520 15.130 121.660 16.090 ;
        RECT 126.010 15.870 128.570 16.210 ;
        RECT 132.120 15.880 140.820 16.220 ;
        RECT 121.000 15.070 121.660 15.130 ;
        RECT 121.060 14.990 121.660 15.070 ;
        RECT 121.520 14.370 121.660 14.990 ;
        RECT 140.490 14.800 141.360 15.130 ;
        RECT 121.460 14.050 121.720 14.370 ;
        RECT 120.540 13.030 120.800 13.350 ;
        RECT 121.460 13.030 121.720 13.350 ;
        RECT 122.380 13.030 122.640 13.350 ;
        RECT 113.630 10.115 113.910 10.485 ;
        RECT 107.930 9.095 109.470 9.465 ;
        RECT 108.110 3.840 108.390 9.095 ;
        RECT 121.520 8.930 121.660 13.030 ;
        RECT 122.440 12.525 122.580 13.030 ;
        RECT 122.370 12.155 122.650 12.525 ;
        RECT 140.490 11.300 140.820 14.800 ;
        RECT 141.030 14.550 141.360 14.630 ;
        RECT 141.510 14.550 141.680 18.200 ;
        RECT 141.030 14.380 143.620 14.550 ;
        RECT 141.030 14.300 141.360 14.380 ;
        RECT 126.010 10.940 128.570 11.280 ;
        RECT 132.120 10.960 140.820 11.300 ;
        RECT 126.010 10.790 126.350 10.940 ;
        RECT 121.460 8.610 121.720 8.930 ;
        RECT 122.380 7.590 122.640 7.910 ;
        RECT 122.440 7.085 122.580 7.590 ;
        RECT 111.230 6.375 112.770 6.745 ;
        RECT 122.370 6.715 122.650 7.085 ;
        RECT 141.040 6.380 141.370 8.350 ;
        RECT 126.010 6.020 128.570 6.360 ;
        RECT 132.120 6.040 141.370 6.380 ;
        RECT 126.010 5.380 126.350 6.020 ;
        RECT 111.200 4.300 112.800 5.140 ;
        RECT 143.240 2.470 143.620 14.380 ;
      LAYER met3 ;
        RECT 85.280 9.920 85.780 41.970 ;
        RECT 87.120 22.160 87.620 41.970 ;
        RECT 89.620 34.400 90.120 41.970 ;
        RECT 107.900 37.420 109.500 38.290 ;
        RECT 124.975 37.880 126.975 38.480 ;
        RECT 120.965 36.970 121.295 36.985 ;
        RECT 125.810 36.970 126.110 37.880 ;
        RECT 120.965 36.670 126.110 36.970 ;
        RECT 120.965 36.655 121.295 36.670 ;
        RECT 107.910 36.315 109.490 36.645 ;
        RECT 89.620 34.250 91.620 34.400 ;
        RECT 110.385 34.250 110.715 34.265 ;
        RECT 89.620 33.950 110.715 34.250 ;
        RECT 89.620 33.800 91.620 33.950 ;
        RECT 110.385 33.935 110.715 33.950 ;
        RECT 122.345 34.250 122.675 34.265 ;
        RECT 122.345 33.950 126.110 34.250 ;
        RECT 122.345 33.935 122.675 33.950 ;
        RECT 111.210 33.595 112.790 33.925 ;
        RECT 125.810 33.040 126.110 33.950 ;
        RECT 124.975 32.440 126.975 33.040 ;
        RECT 107.910 30.875 109.490 31.205 ;
        RECT 122.345 28.810 122.675 28.825 ;
        RECT 122.345 28.510 126.110 28.810 ;
        RECT 122.345 28.495 122.675 28.510 ;
        RECT 111.210 28.155 112.790 28.485 ;
        RECT 125.810 27.600 126.110 28.510 ;
        RECT 124.975 27.000 126.975 27.600 ;
        RECT 107.910 25.435 109.490 25.765 ;
        RECT 122.345 23.370 122.675 23.385 ;
        RECT 122.345 23.070 126.110 23.370 ;
        RECT 122.345 23.055 122.675 23.070 ;
        RECT 111.210 22.715 112.790 23.045 ;
        RECT 125.810 22.160 126.110 23.070 ;
        RECT 87.120 22.010 91.630 22.160 ;
        RECT 103.485 22.010 103.815 22.025 ;
        RECT 87.120 21.710 103.815 22.010 ;
        RECT 87.120 21.560 91.630 21.710 ;
        RECT 103.485 21.695 103.815 21.710 ;
        RECT 124.975 21.560 126.975 22.160 ;
        RECT 107.910 19.995 109.490 20.325 ;
        RECT 111.210 17.275 112.790 17.605 ;
        RECT 122.345 16.570 122.675 16.585 ;
        RECT 124.975 16.570 126.975 16.720 ;
        RECT 122.345 16.270 126.975 16.570 ;
        RECT 122.345 16.255 122.675 16.270 ;
        RECT 124.890 16.120 126.975 16.270 ;
        RECT 124.890 16.100 126.110 16.120 ;
        RECT 107.910 14.555 109.490 14.885 ;
        RECT 122.345 12.490 122.675 12.505 ;
        RECT 122.345 12.190 126.110 12.490 ;
        RECT 122.345 12.175 122.675 12.190 ;
        RECT 111.210 11.835 112.790 12.165 ;
        RECT 125.810 11.280 126.110 12.190 ;
        RECT 124.975 10.680 126.975 11.280 ;
        RECT 113.605 10.450 113.935 10.465 ;
        RECT 101.890 10.150 113.935 10.450 ;
        RECT 85.280 9.770 91.620 9.920 ;
        RECT 101.890 9.770 102.190 10.150 ;
        RECT 113.605 10.135 113.935 10.150 ;
        RECT 85.280 9.470 102.190 9.770 ;
        RECT 85.280 9.320 91.620 9.470 ;
        RECT 107.910 9.115 109.490 9.445 ;
        RECT 122.345 7.050 122.675 7.065 ;
        RECT 122.345 6.750 126.110 7.050 ;
        RECT 122.345 6.735 122.675 6.750 ;
        RECT 111.210 6.395 112.790 6.725 ;
        RECT 125.810 5.840 126.110 6.750 ;
        RECT 124.975 5.240 126.975 5.840 ;
        RECT 111.200 4.300 112.800 5.140 ;
        RECT 143.220 2.390 152.530 2.890 ;
      LAYER met4 ;
        RECT 30.670 223.780 30.970 224.760 ;
        RECT 33.430 223.780 33.730 224.760 ;
        RECT 36.190 223.780 36.490 224.760 ;
        RECT 38.950 223.780 39.250 224.760 ;
        RECT 41.710 223.780 42.010 224.760 ;
        RECT 44.470 223.780 44.770 224.760 ;
        RECT 47.230 223.780 47.530 224.760 ;
        RECT 49.990 223.780 50.290 224.760 ;
        RECT 52.750 223.780 53.050 224.760 ;
        RECT 55.510 223.780 55.810 224.760 ;
        RECT 58.270 223.780 58.570 224.760 ;
        RECT 61.030 223.780 61.330 224.760 ;
        RECT 63.790 223.780 64.090 224.760 ;
        RECT 66.550 223.780 66.850 224.760 ;
        RECT 69.310 223.780 69.610 224.760 ;
        RECT 72.070 223.780 72.370 224.760 ;
        RECT 74.830 223.780 75.130 224.760 ;
        RECT 77.590 223.780 77.890 224.760 ;
        RECT 80.350 223.780 80.650 224.760 ;
        RECT 83.110 223.780 83.410 224.760 ;
        RECT 85.870 223.780 86.170 224.760 ;
        RECT 5.670 223.770 86.170 223.780 ;
        RECT 4.000 223.480 86.170 223.770 ;
        RECT 4.000 220.760 6.000 223.480 ;
        RECT 88.630 222.150 88.930 224.760 ;
        RECT 85.270 221.850 88.930 222.150 ;
        RECT 85.280 41.470 85.780 221.850 ;
        RECT 91.390 220.750 91.690 224.760 ;
        RECT 87.120 220.450 91.690 220.750 ;
        RECT 87.120 41.470 87.620 220.450 ;
        RECT 94.150 219.580 94.450 224.760 ;
        RECT 89.620 219.280 94.450 219.580 ;
        RECT 89.620 41.470 90.120 219.280 ;
        RECT 6.000 38.750 112.800 40.770 ;
        RECT 1.000 4.240 3.000 5.000 ;
        RECT 107.900 4.240 109.500 38.290 ;
        RECT 111.200 4.300 112.800 38.750 ;
        RECT 1.000 2.220 109.500 4.240 ;
        RECT 151.810 1.000 152.710 2.970 ;
  END
END tt_um_emmersonv_tiq_adc
END LIBRARY

