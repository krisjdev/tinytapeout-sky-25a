VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_cw_vref
  CLASS BLOCK ;
  FOREIGN tt_um_cw_vref ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 4.640000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNADIFFAREA 4.640000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 320.000000 ;
    ANTENNADIFFAREA 9.280000 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 969.314453 ;
    ANTENNADIFFAREA 952.880676 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1730.705933 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    USE POWER ;
    ANTENNAGATEAREA 969.314453 ;
    ANTENNADIFFAREA 952.880676 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.600 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.600 5.000 5.200 220.760 ;
    END
  END VGND
  PIN VAPWR
    USE POWER ;
    ANTENNAGATEAREA 2912.000000 ;
    ANTENNADIFFAREA 2005.394531 ;
    PORT
      LAYER met4 ;
        RECT 6.200 5.000 7.800 220.760 ;
    END
  END VAPWR
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  OBS
      LAYER nwell ;
        RECT 3.250 220.980 103.675 223.480 ;
        RECT 3.250 5.750 5.750 220.980 ;
        RECT 8.935 180.290 45.725 212.250 ;
        RECT 48.860 187.290 56.700 210.740 ;
      LAYER pwell ;
        RECT 9.140 168.330 52.250 178.810 ;
      LAYER nwell ;
        RECT 62.865 170.855 99.075 217.105 ;
        RECT 101.175 182.070 103.675 220.980 ;
        RECT 108.240 216.015 153.520 220.985 ;
        RECT 108.240 203.045 153.520 214.015 ;
      LAYER pwell ;
        RECT 108.440 184.690 153.320 201.100 ;
      LAYER nwell ;
        RECT 164.960 200.075 239.400 201.680 ;
      LAYER pwell ;
        RECT 165.155 198.875 166.525 199.685 ;
        RECT 166.535 198.875 167.905 199.685 ;
        RECT 171.160 199.555 172.505 199.785 ;
        RECT 167.925 198.875 170.665 199.555 ;
        RECT 170.675 198.875 172.505 199.555 ;
        RECT 172.515 198.875 178.025 199.685 ;
        RECT 178.045 198.960 178.475 199.745 ;
        RECT 178.980 199.555 180.325 199.785 ;
        RECT 178.495 198.875 180.325 199.555 ;
        RECT 180.335 198.875 185.845 199.685 ;
        RECT 185.855 198.875 187.685 199.685 ;
        RECT 188.155 199.555 189.500 199.785 ;
        RECT 188.155 198.875 189.985 199.555 ;
        RECT 190.925 198.960 191.355 199.745 ;
        RECT 191.375 198.875 196.885 199.685 ;
        RECT 197.815 199.555 199.160 199.785 ;
        RECT 197.815 198.875 199.645 199.555 ;
        RECT 199.655 198.875 203.325 199.685 ;
        RECT 203.805 198.960 204.235 199.745 ;
        RECT 204.255 198.875 207.005 199.685 ;
        RECT 207.475 199.555 208.820 199.785 ;
        RECT 207.475 198.875 209.305 199.555 ;
        RECT 209.315 198.875 214.825 199.685 ;
        RECT 214.835 198.875 216.665 199.685 ;
        RECT 216.685 198.960 217.115 199.745 ;
        RECT 217.135 198.875 219.875 199.555 ;
        RECT 219.895 198.875 225.405 199.685 ;
        RECT 225.415 198.875 226.785 199.685 ;
        RECT 227.280 199.555 228.625 199.785 ;
        RECT 226.795 198.875 228.625 199.555 ;
        RECT 229.565 198.960 229.995 199.745 ;
        RECT 230.015 198.875 235.525 199.685 ;
        RECT 236.480 199.555 237.825 199.785 ;
        RECT 235.995 198.875 237.825 199.555 ;
        RECT 237.835 198.875 239.205 199.685 ;
        RECT 165.295 198.665 165.465 198.875 ;
        RECT 166.675 198.665 166.845 198.875 ;
        RECT 170.355 198.685 170.525 198.875 ;
        RECT 170.815 198.685 170.985 198.875 ;
        RECT 172.195 198.665 172.365 198.855 ;
        RECT 172.655 198.685 172.825 198.875 ;
        RECT 177.715 198.665 177.885 198.855 ;
        RECT 178.635 198.685 178.805 198.875 ;
        RECT 180.475 198.685 180.645 198.875 ;
        RECT 183.235 198.665 183.405 198.855 ;
        RECT 185.995 198.685 186.165 198.875 ;
        RECT 187.830 198.715 187.950 198.825 ;
        RECT 188.755 198.665 188.925 198.855 ;
        RECT 189.675 198.685 189.845 198.875 ;
        RECT 190.145 198.720 190.305 198.830 ;
        RECT 190.590 198.715 190.710 198.825 ;
        RECT 191.515 198.665 191.685 198.875 ;
        RECT 197.035 198.665 197.205 198.855 ;
        RECT 199.335 198.685 199.505 198.875 ;
        RECT 199.795 198.685 199.965 198.875 ;
        RECT 202.555 198.665 202.725 198.855 ;
        RECT 203.470 198.715 203.590 198.825 ;
        RECT 204.395 198.685 204.565 198.875 ;
        RECT 207.150 198.715 207.270 198.825 ;
        RECT 208.075 198.665 208.245 198.855 ;
        RECT 208.995 198.685 209.165 198.875 ;
        RECT 209.455 198.685 209.625 198.875 ;
        RECT 213.595 198.665 213.765 198.855 ;
        RECT 214.975 198.685 215.145 198.875 ;
        RECT 216.350 198.715 216.470 198.825 ;
        RECT 217.275 198.665 217.445 198.875 ;
        RECT 220.035 198.685 220.205 198.875 ;
        RECT 222.795 198.665 222.965 198.855 ;
        RECT 225.555 198.685 225.725 198.875 ;
        RECT 226.935 198.685 227.105 198.875 ;
        RECT 228.315 198.665 228.485 198.855 ;
        RECT 228.785 198.720 228.945 198.830 ;
        RECT 230.155 198.685 230.325 198.875 ;
        RECT 233.835 198.665 234.005 198.855 ;
        RECT 235.670 198.715 235.790 198.825 ;
        RECT 236.135 198.685 236.305 198.875 ;
        RECT 237.510 198.715 237.630 198.825 ;
        RECT 238.895 198.665 239.065 198.875 ;
        RECT 165.155 197.855 166.525 198.665 ;
        RECT 166.535 197.855 172.045 198.665 ;
        RECT 172.055 197.855 177.565 198.665 ;
        RECT 177.575 197.855 183.085 198.665 ;
        RECT 183.095 197.855 188.605 198.665 ;
        RECT 188.615 197.855 190.445 198.665 ;
        RECT 190.925 197.795 191.355 198.580 ;
        RECT 191.375 197.855 196.885 198.665 ;
        RECT 196.895 197.855 202.405 198.665 ;
        RECT 202.415 197.855 207.925 198.665 ;
        RECT 207.935 197.855 213.445 198.665 ;
        RECT 213.455 197.855 216.205 198.665 ;
        RECT 216.685 197.795 217.115 198.580 ;
        RECT 217.135 197.855 222.645 198.665 ;
        RECT 222.655 197.855 228.165 198.665 ;
        RECT 228.175 197.855 233.685 198.665 ;
        RECT 233.695 197.855 237.365 198.665 ;
        RECT 237.835 197.855 239.205 198.665 ;
      LAYER nwell ;
        RECT 164.960 194.635 239.400 197.465 ;
      LAYER pwell ;
        RECT 165.155 193.435 166.525 194.245 ;
        RECT 166.535 193.435 172.045 194.245 ;
        RECT 172.055 193.435 177.565 194.245 ;
        RECT 178.045 193.520 178.475 194.305 ;
        RECT 178.495 193.435 184.005 194.245 ;
        RECT 184.015 193.435 187.685 194.245 ;
        RECT 187.695 193.435 189.065 194.245 ;
        RECT 189.075 193.435 191.825 194.345 ;
        RECT 191.835 193.435 195.505 194.245 ;
        RECT 195.525 193.435 196.875 194.345 ;
        RECT 196.895 193.435 202.405 194.245 ;
        RECT 202.415 193.435 203.785 194.245 ;
        RECT 203.805 193.520 204.235 194.305 ;
        RECT 204.255 193.435 209.765 194.245 ;
        RECT 209.775 193.435 215.285 194.245 ;
        RECT 215.295 193.435 220.805 194.245 ;
        RECT 220.815 193.435 226.325 194.245 ;
        RECT 226.335 193.435 229.085 194.245 ;
        RECT 229.565 193.520 229.995 194.305 ;
        RECT 230.015 193.435 235.525 194.245 ;
        RECT 235.535 193.435 237.365 194.245 ;
        RECT 237.835 193.435 239.205 194.245 ;
        RECT 165.295 193.225 165.465 193.435 ;
        RECT 166.675 193.225 166.845 193.435 ;
        RECT 172.195 193.225 172.365 193.435 ;
        RECT 174.030 193.275 174.150 193.385 ;
        RECT 175.415 193.225 175.585 193.415 ;
        RECT 175.870 193.275 175.990 193.385 ;
        RECT 177.255 193.225 177.425 193.415 ;
        RECT 177.710 193.275 177.830 193.385 ;
        RECT 178.175 193.225 178.345 193.415 ;
        RECT 178.635 193.245 178.805 193.435 ;
        RECT 165.155 192.415 166.525 193.225 ;
        RECT 166.535 192.415 172.045 193.225 ;
        RECT 172.055 192.415 173.885 193.225 ;
        RECT 174.355 192.445 175.725 193.225 ;
        RECT 176.195 192.445 177.565 193.225 ;
        RECT 178.035 192.315 180.785 193.225 ;
        RECT 180.940 193.195 181.110 193.415 ;
        RECT 183.700 193.225 183.870 193.415 ;
        RECT 184.155 193.245 184.325 193.435 ;
        RECT 187.385 193.270 187.545 193.380 ;
        RECT 187.835 193.245 188.005 193.435 ;
        RECT 182.600 193.195 183.545 193.225 ;
        RECT 180.795 192.515 183.545 193.195 ;
        RECT 182.600 192.315 183.545 192.515 ;
        RECT 183.555 192.315 187.210 193.225 ;
        RECT 188.300 193.195 188.470 193.415 ;
        RECT 189.215 193.245 189.385 193.435 ;
        RECT 191.525 193.270 191.685 193.380 ;
        RECT 191.975 193.245 192.145 193.435 ;
        RECT 192.440 193.225 192.610 193.415 ;
        RECT 195.655 193.245 195.825 193.435 ;
        RECT 196.115 193.225 196.285 193.415 ;
        RECT 197.035 193.245 197.205 193.435 ;
        RECT 198.870 193.275 198.990 193.385 ;
        RECT 199.335 193.225 199.505 193.415 ;
        RECT 202.095 193.225 202.265 193.415 ;
        RECT 202.555 193.245 202.725 193.435 ;
        RECT 204.395 193.245 204.565 193.435 ;
        RECT 207.615 193.225 207.785 193.415 ;
        RECT 209.915 193.245 210.085 193.435 ;
        RECT 213.135 193.225 213.305 193.415 ;
        RECT 215.435 193.245 215.605 193.435 ;
        RECT 217.275 193.225 217.445 193.415 ;
        RECT 220.955 193.245 221.125 193.435 ;
        RECT 222.795 193.225 222.965 193.415 ;
        RECT 226.475 193.245 226.645 193.435 ;
        RECT 228.315 193.225 228.485 193.415 ;
        RECT 229.230 193.275 229.350 193.385 ;
        RECT 230.155 193.245 230.325 193.435 ;
        RECT 233.835 193.225 234.005 193.415 ;
        RECT 235.675 193.245 235.845 193.435 ;
        RECT 237.510 193.275 237.630 193.385 ;
        RECT 238.895 193.225 239.065 193.435 ;
        RECT 189.960 193.195 190.905 193.225 ;
        RECT 188.155 192.515 190.905 193.195 ;
        RECT 189.960 192.315 190.905 192.515 ;
        RECT 190.925 192.355 191.355 193.140 ;
        RECT 192.295 192.315 195.950 193.225 ;
        RECT 195.975 192.415 198.725 193.225 ;
        RECT 199.195 192.315 201.945 193.225 ;
        RECT 201.955 192.415 207.465 193.225 ;
        RECT 207.475 192.415 212.985 193.225 ;
        RECT 212.995 192.415 216.665 193.225 ;
        RECT 216.685 192.355 217.115 193.140 ;
        RECT 217.135 192.415 222.645 193.225 ;
        RECT 222.655 192.415 228.165 193.225 ;
        RECT 228.175 192.415 233.685 193.225 ;
        RECT 233.695 192.415 237.365 193.225 ;
        RECT 237.835 192.415 239.205 193.225 ;
      LAYER nwell ;
        RECT 164.960 189.195 239.400 192.025 ;
      LAYER pwell ;
        RECT 165.155 187.995 166.525 188.805 ;
        RECT 166.535 187.995 167.905 188.775 ;
        RECT 167.915 187.995 171.585 188.805 ;
        RECT 171.595 187.995 172.965 188.775 ;
        RECT 173.115 187.995 176.565 188.905 ;
        RECT 176.655 187.995 178.025 188.775 ;
        RECT 178.045 188.080 178.475 188.865 ;
        RECT 178.495 187.995 181.245 188.905 ;
        RECT 181.715 187.995 183.085 188.775 ;
        RECT 183.555 187.995 184.925 188.775 ;
        RECT 185.395 187.995 186.765 188.775 ;
        RECT 187.235 187.995 188.605 188.775 ;
        RECT 188.615 187.995 189.985 188.775 ;
        RECT 191.800 188.705 192.745 188.905 ;
        RECT 189.995 188.025 192.745 188.705 ;
        RECT 165.295 187.785 165.465 187.995 ;
        RECT 166.685 187.975 166.855 187.995 ;
        RECT 166.675 187.805 166.855 187.975 ;
        RECT 168.055 187.805 168.225 187.995 ;
        RECT 166.675 187.785 166.845 187.805 ;
        RECT 168.515 187.785 168.685 187.975 ;
        RECT 169.895 187.785 170.065 187.975 ;
        RECT 171.275 187.785 171.445 187.975 ;
        RECT 171.735 187.805 171.905 187.995 ;
        RECT 176.335 187.785 176.505 187.995 ;
        RECT 176.795 187.805 176.965 187.995 ;
        RECT 178.635 187.805 178.805 187.995 ;
        RECT 180.015 187.785 180.185 187.975 ;
        RECT 181.395 187.945 181.565 187.975 ;
        RECT 180.485 187.830 180.645 187.940 ;
        RECT 181.390 187.835 181.565 187.945 ;
        RECT 181.395 187.785 181.565 187.835 ;
        RECT 182.775 187.785 182.945 187.995 ;
        RECT 183.230 187.835 183.350 187.945 ;
        RECT 183.695 187.805 183.865 187.995 ;
        RECT 185.075 187.945 185.245 187.975 ;
        RECT 185.070 187.835 185.245 187.945 ;
        RECT 185.075 187.785 185.245 187.835 ;
        RECT 185.535 187.785 185.705 187.995 ;
        RECT 186.915 187.945 187.085 187.975 ;
        RECT 186.910 187.835 187.085 187.945 ;
        RECT 186.915 187.785 187.085 187.835 ;
        RECT 187.375 187.805 187.545 187.995 ;
        RECT 165.155 186.975 166.525 187.785 ;
        RECT 166.535 186.975 168.365 187.785 ;
        RECT 168.375 187.005 169.745 187.785 ;
        RECT 169.755 187.005 171.125 187.785 ;
        RECT 171.135 187.105 172.965 187.785 ;
        RECT 171.620 186.875 172.965 187.105 ;
        RECT 173.115 186.875 176.565 187.785 ;
        RECT 176.795 186.875 180.245 187.785 ;
        RECT 181.255 187.005 182.625 187.785 ;
        RECT 182.635 187.005 184.005 187.785 ;
        RECT 184.015 187.005 185.385 187.785 ;
        RECT 185.395 187.005 186.765 187.785 ;
        RECT 186.775 187.005 188.145 187.785 ;
        RECT 188.300 187.755 188.470 187.975 ;
        RECT 189.675 187.805 189.845 187.995 ;
        RECT 190.140 187.805 190.310 188.025 ;
        RECT 191.800 187.995 192.745 188.025 ;
        RECT 192.755 187.995 194.125 188.775 ;
        RECT 194.135 187.995 197.790 188.905 ;
        RECT 197.815 187.995 199.185 188.775 ;
        RECT 199.195 187.995 202.865 188.805 ;
        RECT 203.805 188.080 204.235 188.865 ;
        RECT 204.255 187.995 207.925 188.805 ;
        RECT 208.395 187.995 211.145 188.905 ;
        RECT 211.155 187.995 216.665 188.805 ;
        RECT 216.675 187.995 222.185 188.805 ;
        RECT 222.195 187.995 225.865 188.805 ;
        RECT 226.335 187.995 229.085 188.905 ;
        RECT 229.565 188.080 229.995 188.865 ;
        RECT 230.015 187.995 231.385 188.775 ;
        RECT 231.395 187.995 232.765 188.775 ;
        RECT 232.775 187.995 234.145 188.775 ;
        RECT 234.155 187.995 237.825 188.805 ;
        RECT 237.835 187.995 239.205 188.805 ;
        RECT 191.525 187.830 191.685 187.940 ;
        RECT 192.440 187.785 192.610 187.975 ;
        RECT 192.895 187.805 193.065 187.995 ;
        RECT 194.280 187.805 194.450 187.995 ;
        RECT 196.120 187.785 196.290 187.975 ;
        RECT 198.875 187.805 199.045 187.995 ;
        RECT 199.335 187.805 199.505 187.995 ;
        RECT 199.800 187.785 199.970 187.975 ;
        RECT 203.025 187.840 203.185 187.950 ;
        RECT 203.475 187.785 203.645 187.975 ;
        RECT 204.395 187.805 204.565 187.995 ;
        RECT 208.070 187.835 208.190 187.945 ;
        RECT 208.535 187.805 208.705 187.995 ;
        RECT 208.995 187.785 209.165 187.975 ;
        RECT 210.835 187.785 211.005 187.975 ;
        RECT 211.295 187.805 211.465 187.995 ;
        RECT 212.215 187.785 212.385 187.975 ;
        RECT 213.595 187.785 213.765 187.975 ;
        RECT 214.975 187.785 215.145 187.975 ;
        RECT 216.350 187.835 216.470 187.945 ;
        RECT 216.815 187.805 216.985 187.995 ;
        RECT 217.275 187.785 217.445 187.975 ;
        RECT 220.035 187.785 220.205 187.975 ;
        RECT 222.335 187.785 222.505 187.995 ;
        RECT 222.795 187.785 222.965 187.975 ;
        RECT 226.010 187.835 226.130 187.945 ;
        RECT 226.475 187.805 226.645 187.995 ;
        RECT 229.230 187.835 229.350 187.945 ;
        RECT 231.075 187.805 231.245 187.995 ;
        RECT 231.535 187.805 231.705 187.995 ;
        RECT 233.835 187.805 234.005 187.995 ;
        RECT 234.295 187.805 234.465 187.995 ;
        RECT 234.755 187.785 234.925 187.975 ;
        RECT 236.135 187.785 236.305 187.975 ;
        RECT 237.515 187.785 237.685 187.975 ;
        RECT 238.895 187.785 239.065 187.995 ;
        RECT 189.960 187.755 190.905 187.785 ;
        RECT 188.155 187.075 190.905 187.755 ;
        RECT 189.960 186.875 190.905 187.075 ;
        RECT 190.925 186.915 191.355 187.700 ;
        RECT 192.295 186.875 195.950 187.785 ;
        RECT 195.975 186.875 199.630 187.785 ;
        RECT 199.655 186.875 203.310 187.785 ;
        RECT 203.335 186.975 208.845 187.785 ;
        RECT 208.855 187.105 210.685 187.785 ;
        RECT 209.340 186.875 210.685 187.105 ;
        RECT 210.695 187.005 212.065 187.785 ;
        RECT 212.075 187.005 213.445 187.785 ;
        RECT 213.455 187.005 214.825 187.785 ;
        RECT 214.835 187.005 216.205 187.785 ;
        RECT 216.685 186.915 217.115 187.700 ;
        RECT 217.135 186.875 219.885 187.785 ;
        RECT 219.895 187.005 221.265 187.785 ;
        RECT 221.275 187.005 222.645 187.785 ;
        RECT 222.655 187.615 224.415 187.785 ;
        RECT 222.655 187.570 224.910 187.615 ;
        RECT 222.655 187.535 225.850 187.570 ;
        RECT 227.210 187.535 232.305 187.785 ;
        RECT 222.655 187.105 232.305 187.535 ;
        RECT 223.980 186.935 227.210 187.105 ;
        RECT 224.920 186.890 227.210 186.935 ;
        RECT 225.860 186.855 227.210 186.890 ;
        RECT 230.285 186.875 232.305 187.105 ;
        RECT 232.315 186.875 235.065 187.785 ;
        RECT 235.075 187.005 236.445 187.785 ;
        RECT 236.455 187.005 237.825 187.785 ;
        RECT 237.835 186.975 239.205 187.785 ;
        RECT 230.285 186.855 231.205 186.875 ;
      LAYER nwell ;
        RECT 164.960 183.755 239.400 186.585 ;
      LAYER pwell ;
        RECT 208.575 183.465 209.495 183.485 ;
        RECT 165.155 182.555 166.525 183.365 ;
        RECT 166.535 182.555 167.905 183.335 ;
        RECT 167.915 182.555 169.285 183.335 ;
        RECT 169.295 182.555 170.665 183.335 ;
        RECT 170.815 182.555 174.265 183.465 ;
        RECT 174.370 182.555 178.025 183.465 ;
        RECT 178.045 182.640 178.475 183.425 ;
        RECT 178.510 182.555 182.165 183.465 ;
        RECT 182.315 182.555 185.765 183.465 ;
        RECT 186.775 182.555 188.145 183.335 ;
        RECT 189.960 183.265 190.905 183.465 ;
        RECT 192.720 183.265 193.665 183.465 ;
        RECT 188.155 182.585 190.905 183.265 ;
        RECT 190.915 182.585 193.665 183.265 ;
        RECT 165.295 182.345 165.465 182.555 ;
        RECT 166.675 182.345 166.845 182.555 ;
        RECT 168.055 182.365 168.225 182.555 ;
        RECT 168.515 182.345 168.685 182.535 ;
        RECT 169.435 182.365 169.605 182.555 ;
        RECT 169.895 182.345 170.065 182.535 ;
        RECT 174.035 182.365 174.205 182.555 ;
        RECT 174.955 182.345 175.125 182.535 ;
        RECT 177.710 182.365 177.880 182.555 ;
        RECT 178.635 182.345 178.805 182.535 ;
      LAYER nwell ;
        RECT 101.175 179.570 156.750 182.070 ;
      LAYER pwell ;
        RECT 165.155 181.535 166.525 182.345 ;
        RECT 166.535 181.665 168.365 182.345 ;
        RECT 168.375 181.565 169.745 182.345 ;
        RECT 169.755 181.535 171.585 182.345 ;
        RECT 171.735 181.435 175.185 182.345 ;
        RECT 175.415 181.435 178.865 182.345 ;
        RECT 178.955 182.315 179.900 182.345 ;
        RECT 181.390 182.315 181.560 182.535 ;
        RECT 181.850 182.500 182.020 182.555 ;
        RECT 181.850 182.390 182.025 182.500 ;
        RECT 181.850 182.365 182.020 182.390 ;
        RECT 183.050 182.345 183.220 182.535 ;
        RECT 185.535 182.365 185.705 182.555 ;
        RECT 186.005 182.400 186.165 182.510 ;
        RECT 186.915 182.365 187.085 182.555 ;
        RECT 187.190 182.345 187.360 182.535 ;
        RECT 188.300 182.365 188.470 182.585 ;
        RECT 189.960 182.555 190.905 182.585 ;
        RECT 191.060 182.365 191.230 182.585 ;
        RECT 192.720 182.555 193.665 182.585 ;
        RECT 194.595 183.235 195.525 183.465 ;
        RECT 194.595 182.555 198.495 183.235 ;
        RECT 198.735 182.555 201.475 183.235 ;
        RECT 201.955 182.555 203.325 183.335 ;
        RECT 203.805 182.640 204.235 183.425 ;
        RECT 204.255 182.555 205.625 183.335 ;
        RECT 206.095 182.555 207.465 183.335 ;
        RECT 207.475 183.235 209.495 183.465 ;
        RECT 212.570 183.450 213.920 183.485 ;
        RECT 223.100 183.450 224.450 183.485 ;
        RECT 212.570 183.405 214.860 183.450 ;
        RECT 222.160 183.405 224.450 183.450 ;
        RECT 212.570 183.235 215.800 183.405 ;
        RECT 207.475 182.805 217.125 183.235 ;
        RECT 207.475 182.555 212.570 182.805 ;
        RECT 213.930 182.770 217.125 182.805 ;
        RECT 214.870 182.725 217.125 182.770 ;
        RECT 215.365 182.555 217.125 182.725 ;
        RECT 217.135 182.555 218.505 183.335 ;
        RECT 218.515 182.555 219.885 183.335 ;
        RECT 221.220 183.235 224.450 183.405 ;
        RECT 227.525 183.465 228.445 183.485 ;
        RECT 227.525 183.235 229.545 183.465 ;
        RECT 219.895 182.805 229.545 183.235 ;
        RECT 219.895 182.770 223.090 182.805 ;
        RECT 219.895 182.725 222.150 182.770 ;
        RECT 219.895 182.555 221.655 182.725 ;
        RECT 224.450 182.555 229.545 182.805 ;
        RECT 229.565 182.640 229.995 183.425 ;
        RECT 230.015 182.555 231.385 183.335 ;
        RECT 231.395 182.555 232.765 183.335 ;
        RECT 232.775 182.555 234.145 183.335 ;
        RECT 234.155 182.555 235.525 183.335 ;
        RECT 235.535 182.555 236.905 183.335 ;
        RECT 237.835 182.555 239.205 183.365 ;
        RECT 191.525 182.390 191.685 182.500 ;
        RECT 193.825 182.400 193.985 182.510 ;
        RECT 195.010 182.365 195.180 182.555 ;
        RECT 195.840 182.345 196.010 182.535 ;
        RECT 196.850 182.345 197.020 182.535 ;
        RECT 198.875 182.365 199.045 182.555 ;
        RECT 200.990 182.345 201.160 182.535 ;
        RECT 201.630 182.395 201.750 182.505 ;
        RECT 203.015 182.365 203.185 182.555 ;
        RECT 203.470 182.395 203.590 182.505 ;
        RECT 204.395 182.365 204.565 182.555 ;
        RECT 205.775 182.505 205.945 182.535 ;
        RECT 204.865 182.390 205.025 182.500 ;
        RECT 205.770 182.395 205.945 182.505 ;
        RECT 205.775 182.345 205.945 182.395 ;
        RECT 206.235 182.365 206.405 182.555 ;
        RECT 216.355 182.345 216.525 182.535 ;
        RECT 216.815 182.365 216.985 182.555 ;
        RECT 218.195 182.365 218.365 182.555 ;
        RECT 218.655 182.365 218.825 182.555 ;
        RECT 220.035 182.365 220.205 182.555 ;
        RECT 225.095 182.345 225.265 182.535 ;
        RECT 225.555 182.345 225.725 182.535 ;
        RECT 226.935 182.345 227.105 182.535 ;
        RECT 230.155 182.365 230.325 182.555 ;
        RECT 232.455 182.365 232.625 182.555 ;
        RECT 233.835 182.365 234.005 182.555 ;
        RECT 235.215 182.365 235.385 182.555 ;
        RECT 236.595 182.365 236.765 182.555 ;
        RECT 237.065 182.400 237.225 182.510 ;
        RECT 237.515 182.345 237.685 182.535 ;
        RECT 238.895 182.345 239.065 182.555 ;
        RECT 178.955 181.635 181.705 182.315 ;
        RECT 182.635 181.665 186.535 182.345 ;
        RECT 186.775 181.665 190.675 182.345 ;
        RECT 178.955 181.435 179.900 181.635 ;
        RECT 182.635 181.435 183.565 181.665 ;
        RECT 186.775 181.435 187.705 181.665 ;
        RECT 190.925 181.475 191.355 182.260 ;
        RECT 192.525 181.665 196.425 182.345 ;
        RECT 195.495 181.435 196.425 181.665 ;
        RECT 196.435 181.665 200.335 182.345 ;
        RECT 200.575 181.665 204.475 182.345 ;
        RECT 196.435 181.435 197.365 181.665 ;
        RECT 200.575 181.435 201.505 181.665 ;
        RECT 205.635 181.565 207.005 182.345 ;
        RECT 207.015 182.095 212.110 182.345 ;
        RECT 214.905 182.175 216.665 182.345 ;
        RECT 214.410 182.130 216.665 182.175 ;
        RECT 213.470 182.095 216.665 182.130 ;
        RECT 207.015 181.665 216.665 182.095 ;
        RECT 207.015 181.435 209.035 181.665 ;
        RECT 208.115 181.415 209.035 181.435 ;
        RECT 212.110 181.495 215.340 181.665 ;
        RECT 212.110 181.450 214.400 181.495 ;
        RECT 216.685 181.475 217.115 182.260 ;
        RECT 217.135 181.665 225.405 182.345 ;
        RECT 212.110 181.415 213.460 181.450 ;
        RECT 217.135 181.435 218.585 181.665 ;
        RECT 225.415 181.535 226.785 182.345 ;
        RECT 226.795 182.175 228.555 182.345 ;
        RECT 226.795 182.130 229.050 182.175 ;
        RECT 226.795 182.095 229.990 182.130 ;
        RECT 231.350 182.095 236.445 182.345 ;
        RECT 226.795 181.665 236.445 182.095 ;
        RECT 228.120 181.495 231.350 181.665 ;
        RECT 229.060 181.450 231.350 181.495 ;
        RECT 230.000 181.415 231.350 181.450 ;
        RECT 234.425 181.435 236.445 181.665 ;
        RECT 236.455 181.565 237.825 182.345 ;
        RECT 237.835 181.535 239.205 182.345 ;
        RECT 234.425 181.415 235.345 181.435 ;
        RECT 9.140 147.810 51.970 168.220 ;
      LAYER nwell ;
        RECT 63.050 164.975 97.990 167.475 ;
      LAYER pwell ;
        RECT 9.600 134.835 20.550 138.315 ;
        RECT 23.425 135.385 58.475 143.515 ;
      LAYER nwell ;
        RECT 63.050 135.035 65.550 164.975 ;
        RECT 69.300 160.385 91.740 161.225 ;
        RECT 69.300 139.625 70.140 160.385 ;
      LAYER pwell ;
        RECT 71.090 158.670 89.950 159.435 ;
        RECT 71.090 156.220 71.855 158.670 ;
        RECT 74.305 156.220 75.575 158.670 ;
        RECT 78.025 156.220 79.295 158.670 ;
        RECT 81.745 156.220 83.015 158.670 ;
        RECT 85.465 156.220 86.735 158.670 ;
        RECT 89.185 156.220 89.950 158.670 ;
        RECT 71.090 154.950 89.950 156.220 ;
        RECT 71.090 152.500 71.855 154.950 ;
        RECT 74.305 152.500 75.575 154.950 ;
        RECT 78.025 152.500 79.295 154.950 ;
        RECT 81.745 152.500 83.015 154.950 ;
        RECT 85.465 152.500 86.735 154.950 ;
        RECT 89.185 152.500 89.950 154.950 ;
        RECT 71.090 151.230 89.950 152.500 ;
        RECT 71.090 148.780 71.855 151.230 ;
        RECT 74.305 148.780 75.575 151.230 ;
        RECT 78.025 148.780 79.295 151.230 ;
        RECT 81.745 148.780 83.015 151.230 ;
        RECT 85.465 148.780 86.735 151.230 ;
        RECT 89.185 148.780 89.950 151.230 ;
        RECT 71.090 147.510 89.950 148.780 ;
        RECT 71.090 145.060 71.855 147.510 ;
        RECT 74.305 145.060 75.575 147.510 ;
        RECT 78.025 145.060 79.295 147.510 ;
        RECT 81.745 145.060 83.015 147.510 ;
        RECT 85.465 145.060 86.735 147.510 ;
        RECT 89.185 145.060 89.950 147.510 ;
        RECT 71.090 143.790 89.950 145.060 ;
        RECT 71.090 141.340 71.855 143.790 ;
        RECT 74.305 141.340 75.575 143.790 ;
        RECT 78.025 141.340 79.295 143.790 ;
        RECT 81.745 141.340 83.015 143.790 ;
        RECT 85.465 141.340 86.735 143.790 ;
        RECT 89.185 141.340 89.950 143.790 ;
        RECT 71.090 140.575 89.950 141.340 ;
      LAYER nwell ;
        RECT 90.900 139.625 91.740 160.385 ;
        RECT 69.300 138.785 91.740 139.625 ;
        RECT 95.490 135.035 97.990 164.975 ;
      LAYER pwell ;
        RECT 102.550 158.280 111.160 172.690 ;
        RECT 114.030 166.235 151.540 176.715 ;
      LAYER nwell ;
        RECT 102.350 141.345 111.360 156.335 ;
        RECT 115.985 139.690 149.475 158.060 ;
        RECT 63.050 132.535 97.990 135.035 ;
        RECT 138.080 129.720 145.960 134.690 ;
      LAYER pwell ;
        RECT 138.280 124.290 145.760 128.770 ;
      LAYER nwell ;
        RECT 10.025 41.635 128.935 124.285 ;
      LAYER pwell ;
        RECT 10.225 9.090 74.495 39.430 ;
        RECT 79.865 9.090 128.735 39.430 ;
      LAYER nwell ;
        RECT 135.120 13.460 149.570 109.050 ;
        RECT 154.250 5.750 156.750 179.570 ;
        RECT 164.960 178.315 239.400 181.145 ;
      LAYER pwell ;
        RECT 208.115 178.025 209.035 178.045 ;
        RECT 165.155 177.115 166.525 177.925 ;
        RECT 167.455 177.115 168.825 177.895 ;
        RECT 168.835 177.115 170.665 177.795 ;
        RECT 170.815 177.115 174.265 178.025 ;
        RECT 174.365 177.115 177.105 177.795 ;
        RECT 178.045 177.200 178.475 177.985 ;
        RECT 178.495 177.825 179.440 178.025 ;
        RECT 178.495 177.145 181.245 177.825 ;
        RECT 178.495 177.115 179.440 177.145 ;
        RECT 165.295 176.925 165.465 177.115 ;
        RECT 166.685 176.960 166.845 177.070 ;
        RECT 167.595 176.925 167.765 177.115 ;
        RECT 168.975 176.925 169.145 177.115 ;
        RECT 174.035 176.925 174.205 177.115 ;
        RECT 176.795 176.925 176.965 177.115 ;
        RECT 177.265 176.960 177.425 177.070 ;
        RECT 180.930 176.925 181.100 177.145 ;
        RECT 181.255 177.115 182.625 177.895 ;
        RECT 182.635 177.795 183.565 178.025 ;
        RECT 182.635 177.115 186.535 177.795 ;
        RECT 186.775 177.115 188.145 177.895 ;
        RECT 188.155 177.115 189.525 177.895 ;
        RECT 189.535 177.115 190.905 177.895 ;
        RECT 190.925 177.200 191.355 177.985 ;
        RECT 191.835 177.115 193.205 177.895 ;
        RECT 193.215 177.115 194.585 177.895 ;
        RECT 194.595 177.115 195.965 177.895 ;
        RECT 195.975 177.795 196.905 178.025 ;
        RECT 195.975 177.115 199.875 177.795 ;
        RECT 201.035 177.115 202.405 177.895 ;
        RECT 202.415 177.115 203.785 177.895 ;
        RECT 203.805 177.200 204.235 177.985 ;
        RECT 204.715 177.115 206.085 177.895 ;
        RECT 207.015 177.795 209.035 178.025 ;
        RECT 212.110 178.010 213.460 178.045 ;
        RECT 223.100 178.010 224.450 178.045 ;
        RECT 212.110 177.965 214.400 178.010 ;
        RECT 212.110 177.795 215.340 177.965 ;
        RECT 207.015 177.365 216.665 177.795 ;
        RECT 207.015 177.115 212.110 177.365 ;
        RECT 213.470 177.330 216.665 177.365 ;
        RECT 214.410 177.285 216.665 177.330 ;
        RECT 214.905 177.115 216.665 177.285 ;
        RECT 216.685 177.200 217.115 177.985 ;
        RECT 222.160 177.965 224.450 178.010 ;
        RECT 217.135 177.115 218.505 177.895 ;
        RECT 218.515 177.115 219.885 177.895 ;
        RECT 221.220 177.795 224.450 177.965 ;
        RECT 227.525 178.025 228.445 178.045 ;
        RECT 227.525 177.795 229.545 178.025 ;
        RECT 219.895 177.365 229.545 177.795 ;
        RECT 219.895 177.330 223.090 177.365 ;
        RECT 219.895 177.285 222.150 177.330 ;
        RECT 219.895 177.115 221.655 177.285 ;
        RECT 224.450 177.115 229.545 177.365 ;
        RECT 229.565 177.200 229.995 177.985 ;
        RECT 230.015 177.115 231.385 177.895 ;
        RECT 231.395 177.115 232.765 177.895 ;
        RECT 232.775 177.115 234.145 177.895 ;
        RECT 234.155 177.115 235.525 177.895 ;
        RECT 235.535 177.115 236.905 177.895 ;
        RECT 237.835 177.115 239.205 177.925 ;
        RECT 181.395 176.925 181.565 177.115 ;
        RECT 183.050 176.925 183.220 177.115 ;
        RECT 187.835 176.925 188.005 177.115 ;
        RECT 189.215 176.925 189.385 177.115 ;
        RECT 189.675 176.925 189.845 177.115 ;
        RECT 191.510 176.955 191.630 177.065 ;
        RECT 191.975 176.925 192.145 177.115 ;
        RECT 194.275 176.925 194.445 177.115 ;
        RECT 194.735 176.925 194.905 177.115 ;
        RECT 196.390 176.925 196.560 177.115 ;
        RECT 200.265 176.960 200.425 177.070 ;
        RECT 201.175 176.925 201.345 177.115 ;
        RECT 202.555 176.925 202.725 177.115 ;
        RECT 204.390 176.955 204.510 177.065 ;
        RECT 204.855 176.925 205.025 177.115 ;
        RECT 206.245 176.960 206.405 177.070 ;
        RECT 216.355 176.925 216.525 177.115 ;
        RECT 217.275 176.925 217.445 177.115 ;
        RECT 218.655 176.925 218.825 177.115 ;
        RECT 220.035 176.925 220.205 177.115 ;
        RECT 231.075 176.925 231.245 177.115 ;
        RECT 232.455 176.925 232.625 177.115 ;
        RECT 233.835 176.925 234.005 177.115 ;
        RECT 235.215 176.925 235.385 177.115 ;
        RECT 236.595 176.925 236.765 177.115 ;
        RECT 237.065 176.960 237.225 177.070 ;
        RECT 238.895 176.925 239.065 177.115 ;
        RECT 162.240 106.320 162.410 106.510 ;
        RECT 163.615 106.370 163.735 106.480 ;
        RECT 165.460 106.320 165.630 106.510 ;
        RECT 165.930 106.365 166.090 106.475 ;
        RECT 166.840 106.360 167.010 106.510 ;
        RECT 162.100 105.510 163.470 106.320 ;
        RECT 163.940 105.640 165.770 106.320 ;
        RECT 163.940 105.410 165.285 105.640 ;
        RECT 166.720 105.410 167.610 106.360 ;
        RECT 170.060 106.320 170.230 106.510 ;
        RECT 171.900 106.320 172.070 106.510 ;
        RECT 174.660 106.320 174.830 106.510 ;
        RECT 175.575 106.370 175.695 106.480 ;
        RECT 176.040 106.320 176.210 106.510 ;
        RECT 177.880 106.320 178.050 106.510 ;
        RECT 182.020 106.320 182.190 106.510 ;
        RECT 182.480 106.320 182.650 106.510 ;
        RECT 185.700 106.320 185.870 106.510 ;
        RECT 186.160 106.320 186.330 106.510 ;
        RECT 190.760 106.320 190.930 106.510 ;
        RECT 191.220 106.320 191.390 106.510 ;
        RECT 194.900 106.320 195.070 106.510 ;
        RECT 195.360 106.320 195.530 106.510 ;
        RECT 198.580 106.320 198.750 106.510 ;
        RECT 199.040 106.320 199.210 106.510 ;
        RECT 203.640 106.320 203.810 106.510 ;
        RECT 204.100 106.320 204.270 106.510 ;
        RECT 207.135 106.320 207.305 106.510 ;
        RECT 211.010 106.365 211.170 106.475 ;
        RECT 213.300 106.320 213.470 106.510 ;
        RECT 216.520 106.320 216.690 106.510 ;
        RECT 216.980 106.320 217.150 106.510 ;
        RECT 218.360 106.320 218.530 106.510 ;
        RECT 220.200 106.320 220.370 106.510 ;
        RECT 222.960 106.320 223.130 106.510 ;
        RECT 224.800 106.320 224.970 106.510 ;
        RECT 227.095 106.370 227.215 106.480 ;
        RECT 229.860 106.320 230.030 106.510 ;
        RECT 230.320 106.320 230.490 106.510 ;
        RECT 232.160 106.320 232.330 106.510 ;
        RECT 234.000 106.320 234.170 106.510 ;
        RECT 236.770 106.365 236.930 106.475 ;
        RECT 237.680 106.320 237.850 106.510 ;
        RECT 240.255 106.320 240.425 106.510 ;
        RECT 247.525 106.320 247.695 106.510 ;
        RECT 250.560 106.320 250.730 106.510 ;
        RECT 251.020 106.320 251.190 106.510 ;
        RECT 255.160 106.320 255.330 106.510 ;
        RECT 257.920 106.320 258.090 106.510 ;
        RECT 259.760 106.320 259.930 106.510 ;
        RECT 260.230 106.365 260.390 106.475 ;
        RECT 263.440 106.320 263.610 106.510 ;
        RECT 263.900 106.320 264.070 106.510 ;
        RECT 267.120 106.320 267.290 106.510 ;
        RECT 267.590 106.365 267.750 106.475 ;
        RECT 270.800 106.320 270.970 106.510 ;
        RECT 273.560 106.320 273.730 106.510 ;
        RECT 275.400 106.320 275.570 106.510 ;
        RECT 277.240 106.320 277.410 106.510 ;
        RECT 277.695 106.370 277.815 106.480 ;
        RECT 280.920 106.320 281.090 106.510 ;
        RECT 282.760 106.320 282.930 106.510 ;
        RECT 285.520 106.320 285.690 106.510 ;
        RECT 287.360 106.320 287.530 106.510 ;
        RECT 289.200 106.320 289.370 106.510 ;
        RECT 290.580 106.320 290.750 106.510 ;
        RECT 293.800 106.320 293.970 106.510 ;
        RECT 294.260 106.320 294.430 106.510 ;
        RECT 296.110 106.365 296.270 106.475 ;
        RECT 299.320 106.320 299.490 106.510 ;
        RECT 301.160 106.320 301.330 106.510 ;
        RECT 301.620 106.320 301.790 106.510 ;
        RECT 303.455 106.370 303.575 106.480 ;
        RECT 304.380 106.320 304.550 106.510 ;
        RECT 308.520 106.320 308.690 106.510 ;
        RECT 308.990 106.365 309.150 106.475 ;
        RECT 310.820 106.320 310.990 106.510 ;
        RECT 167.630 105.640 170.370 106.320 ;
        RECT 170.380 105.640 172.210 106.320 ;
        RECT 172.230 105.640 174.970 106.320 ;
        RECT 170.380 105.410 171.725 105.640 ;
        RECT 174.990 105.450 175.420 106.235 ;
        RECT 175.900 105.640 177.730 106.320 ;
        RECT 177.740 105.640 179.570 106.320 ;
        RECT 179.590 105.640 182.330 106.320 ;
        RECT 182.340 105.640 184.170 106.320 ;
        RECT 176.385 105.410 177.730 105.640 ;
        RECT 178.225 105.410 179.570 105.640 ;
        RECT 182.825 105.410 184.170 105.640 ;
        RECT 184.180 105.640 186.010 106.320 ;
        RECT 186.020 105.640 187.850 106.320 ;
        RECT 184.180 105.410 185.525 105.640 ;
        RECT 186.505 105.410 187.850 105.640 ;
        RECT 187.870 105.450 188.300 106.235 ;
        RECT 188.330 105.640 191.070 106.320 ;
        RECT 191.080 105.510 192.450 106.320 ;
        RECT 192.470 105.640 195.210 106.320 ;
        RECT 195.220 105.640 197.050 106.320 ;
        RECT 195.705 105.410 197.050 105.640 ;
        RECT 197.060 105.640 198.890 106.320 ;
        RECT 198.900 105.640 200.730 106.320 ;
        RECT 197.060 105.410 198.405 105.640 ;
        RECT 199.385 105.410 200.730 105.640 ;
        RECT 200.750 105.450 201.180 106.235 ;
        RECT 201.210 105.640 203.950 106.320 ;
        RECT 203.960 105.640 206.700 106.320 ;
        RECT 206.720 105.640 210.620 106.320 ;
        RECT 211.780 105.640 213.610 106.320 ;
        RECT 206.720 105.410 207.650 105.640 ;
        RECT 211.780 105.410 213.125 105.640 ;
        RECT 213.630 105.450 214.060 106.235 ;
        RECT 214.090 105.640 216.830 106.320 ;
        RECT 216.840 105.510 218.210 106.320 ;
        RECT 218.220 105.640 220.050 106.320 ;
        RECT 220.060 105.640 222.800 106.320 ;
        RECT 222.820 105.640 224.650 106.320 ;
        RECT 224.660 105.640 226.490 106.320 ;
        RECT 218.705 105.410 220.050 105.640 ;
        RECT 223.305 105.410 224.650 105.640 ;
        RECT 225.145 105.410 226.490 105.640 ;
        RECT 226.510 105.450 226.940 106.235 ;
        RECT 227.430 105.640 230.170 106.320 ;
        RECT 230.180 105.640 232.010 106.320 ;
        RECT 232.020 105.640 233.850 106.320 ;
        RECT 233.860 105.640 236.600 106.320 ;
        RECT 237.540 105.640 239.370 106.320 ;
        RECT 230.665 105.410 232.010 105.640 ;
        RECT 232.505 105.410 233.850 105.640 ;
        RECT 238.025 105.410 239.370 105.640 ;
        RECT 239.390 105.450 239.820 106.235 ;
        RECT 239.840 105.640 243.740 106.320 ;
        RECT 244.210 105.640 248.110 106.320 ;
        RECT 248.130 105.640 250.870 106.320 ;
        RECT 239.840 105.410 240.770 105.640 ;
        RECT 247.180 105.410 248.110 105.640 ;
        RECT 250.880 105.510 252.250 106.320 ;
        RECT 252.270 105.450 252.700 106.235 ;
        RECT 252.730 105.640 255.470 106.320 ;
        RECT 255.490 105.640 258.230 106.320 ;
        RECT 258.240 105.640 260.070 106.320 ;
        RECT 261.010 105.640 263.750 106.320 ;
        RECT 258.240 105.410 259.585 105.640 ;
        RECT 263.760 105.510 265.130 106.320 ;
        RECT 265.150 105.450 265.580 106.235 ;
        RECT 265.600 105.640 267.430 106.320 ;
        RECT 268.370 105.640 271.110 106.320 ;
        RECT 271.130 105.640 273.870 106.320 ;
        RECT 273.880 105.640 275.710 106.320 ;
        RECT 275.720 105.640 277.550 106.320 ;
        RECT 265.600 105.410 266.945 105.640 ;
        RECT 273.880 105.410 275.225 105.640 ;
        RECT 275.720 105.410 277.065 105.640 ;
        RECT 278.030 105.450 278.460 106.235 ;
        RECT 278.490 105.640 281.230 106.320 ;
        RECT 281.240 105.640 283.070 106.320 ;
        RECT 283.090 105.640 285.830 106.320 ;
        RECT 285.840 105.640 287.670 106.320 ;
        RECT 287.680 105.640 289.510 106.320 ;
        RECT 281.240 105.410 282.585 105.640 ;
        RECT 285.840 105.410 287.185 105.640 ;
        RECT 287.680 105.410 289.025 105.640 ;
        RECT 289.520 105.540 290.890 106.320 ;
        RECT 290.910 105.450 291.340 106.235 ;
        RECT 291.370 105.640 294.110 106.320 ;
        RECT 294.120 105.640 295.950 106.320 ;
        RECT 296.890 105.640 299.630 106.320 ;
        RECT 299.640 105.640 301.470 106.320 ;
        RECT 301.480 105.640 303.310 106.320 ;
        RECT 294.605 105.410 295.950 105.640 ;
        RECT 299.640 105.410 300.985 105.640 ;
        RECT 301.965 105.410 303.310 105.640 ;
        RECT 303.790 105.450 304.220 106.235 ;
        RECT 304.240 105.640 306.980 106.320 ;
        RECT 307.000 105.640 308.830 106.320 ;
        RECT 307.000 105.410 308.345 105.640 ;
        RECT 309.760 105.510 311.130 106.320 ;
      LAYER nwell ;
        RECT 161.905 102.290 311.325 105.120 ;
      LAYER pwell ;
        RECT 162.100 101.090 163.470 101.900 ;
        RECT 163.480 101.090 165.310 101.900 ;
        RECT 169.830 101.770 170.760 101.990 ;
        RECT 173.590 101.770 174.930 102.000 ;
        RECT 165.320 101.090 174.930 101.770 ;
        RECT 174.990 101.175 175.420 101.960 ;
        RECT 175.440 101.770 176.370 102.000 ;
        RECT 179.580 101.770 180.925 102.000 ;
        RECT 185.930 101.770 186.860 101.990 ;
        RECT 189.690 101.770 191.030 102.000 ;
        RECT 195.590 101.770 196.520 101.990 ;
        RECT 199.350 101.770 200.690 102.000 ;
        RECT 175.440 101.090 179.340 101.770 ;
        RECT 179.580 101.090 181.410 101.770 ;
        RECT 181.420 101.090 191.030 101.770 ;
        RECT 191.080 101.090 200.690 101.770 ;
        RECT 200.750 101.175 201.180 101.960 ;
        RECT 201.660 101.090 203.030 101.870 ;
        RECT 203.525 101.770 204.870 102.000 ;
        RECT 209.850 101.770 210.780 101.990 ;
        RECT 213.610 101.770 214.530 102.000 ;
        RECT 221.810 101.770 222.740 101.990 ;
        RECT 225.570 101.770 226.490 102.000 ;
        RECT 203.040 101.090 204.870 101.770 ;
        RECT 205.340 101.090 214.530 101.770 ;
        RECT 214.550 101.090 217.290 101.770 ;
        RECT 217.300 101.090 226.490 101.770 ;
        RECT 226.510 101.175 226.940 101.960 ;
        RECT 231.470 101.770 232.400 101.990 ;
        RECT 235.230 101.770 236.150 102.000 ;
        RECT 226.960 101.090 236.150 101.770 ;
        RECT 236.160 101.770 237.505 102.000 ;
        RECT 242.970 101.770 243.900 101.990 ;
        RECT 246.730 101.770 247.650 102.000 ;
        RECT 236.160 101.090 237.990 101.770 ;
        RECT 238.460 101.090 247.650 101.770 ;
        RECT 247.670 101.090 250.410 101.770 ;
        RECT 250.420 101.090 251.790 101.870 ;
        RECT 252.270 101.175 252.700 101.960 ;
        RECT 252.720 101.770 254.065 102.000 ;
        RECT 252.720 101.090 254.550 101.770 ;
        RECT 255.480 101.090 258.690 102.000 ;
        RECT 258.700 101.090 262.355 102.000 ;
        RECT 262.380 101.090 265.590 102.000 ;
        RECT 265.600 101.770 266.945 102.000 ;
        RECT 265.600 101.090 267.430 101.770 ;
        RECT 267.440 101.090 268.810 101.900 ;
        RECT 268.820 101.770 269.740 102.000 ;
        RECT 272.570 101.770 273.500 101.990 ;
        RECT 268.820 101.090 278.010 101.770 ;
        RECT 278.030 101.175 278.460 101.960 ;
        RECT 281.680 101.770 282.610 102.000 ;
        RECT 278.710 101.090 282.610 101.770 ;
        RECT 282.620 101.770 283.965 102.000 ;
        RECT 289.430 101.770 290.360 101.990 ;
        RECT 293.190 101.770 294.530 102.000 ;
        RECT 282.620 101.090 284.450 101.770 ;
        RECT 284.920 101.090 294.530 101.770 ;
        RECT 294.580 101.770 295.500 102.000 ;
        RECT 298.330 101.770 299.260 101.990 ;
        RECT 294.580 101.090 303.770 101.770 ;
        RECT 303.790 101.175 304.220 101.960 ;
        RECT 304.725 101.770 306.070 102.000 ;
        RECT 304.240 101.090 306.070 101.770 ;
        RECT 307.000 101.090 309.740 101.770 ;
        RECT 309.760 101.090 311.130 101.900 ;
        RECT 162.240 100.880 162.410 101.090 ;
        RECT 163.620 100.880 163.790 101.090 ;
        RECT 165.460 100.880 165.630 101.090 ;
        RECT 168.220 100.880 168.390 101.070 ;
        RECT 168.680 100.880 168.850 101.070 ;
        RECT 175.855 100.900 176.025 101.090 ;
        RECT 178.155 100.880 178.325 101.070 ;
        RECT 181.100 100.900 181.270 101.090 ;
        RECT 181.560 100.900 181.730 101.090 ;
        RECT 182.020 100.880 182.190 101.070 ;
        RECT 183.395 100.930 183.515 101.040 ;
        RECT 184.135 100.880 184.305 101.070 ;
        RECT 188.460 100.880 188.630 101.070 ;
        RECT 191.220 100.900 191.390 101.090 ;
        RECT 201.065 100.880 201.235 101.070 ;
        RECT 201.335 100.930 201.455 101.040 ;
        RECT 201.800 100.900 201.970 101.090 ;
        RECT 203.180 100.900 203.350 101.090 ;
        RECT 205.015 100.930 205.135 101.040 ;
        RECT 205.480 100.900 205.650 101.090 ;
        RECT 210.540 100.880 210.710 101.070 ;
        RECT 211.920 100.880 212.090 101.070 ;
        RECT 212.380 100.880 212.550 101.070 ;
        RECT 214.230 100.925 214.390 101.035 ;
        RECT 215.140 100.880 215.310 101.070 ;
        RECT 216.980 100.880 217.150 101.090 ;
        RECT 217.440 100.900 217.610 101.090 ;
        RECT 218.830 100.925 218.990 101.035 ;
        RECT 219.740 100.920 219.910 101.070 ;
        RECT 220.670 100.925 220.830 101.035 ;
        RECT 162.100 100.070 163.470 100.880 ;
        RECT 163.480 100.070 165.310 100.880 ;
        RECT 165.320 100.100 166.690 100.880 ;
        RECT 166.700 100.200 168.530 100.880 ;
        RECT 168.540 100.200 177.730 100.880 ;
        RECT 166.700 99.970 168.045 100.200 ;
        RECT 173.050 99.980 173.980 100.200 ;
        RECT 176.810 99.970 177.730 100.200 ;
        RECT 177.740 100.200 181.640 100.880 ;
        RECT 177.740 99.970 178.670 100.200 ;
        RECT 181.880 100.100 183.250 100.880 ;
        RECT 183.720 100.200 187.620 100.880 ;
        RECT 183.720 99.970 184.650 100.200 ;
        RECT 187.870 100.010 188.300 100.795 ;
        RECT 188.320 100.200 197.510 100.880 ;
        RECT 197.750 100.200 201.650 100.880 ;
        RECT 192.830 99.980 193.760 100.200 ;
        RECT 196.590 99.970 197.510 100.200 ;
        RECT 200.720 99.970 201.650 100.200 ;
        RECT 201.660 100.200 210.850 100.880 ;
        RECT 201.660 99.970 202.580 100.200 ;
        RECT 205.410 99.980 206.340 100.200 ;
        RECT 210.860 100.100 212.230 100.880 ;
        RECT 212.240 100.070 213.610 100.880 ;
        RECT 213.630 100.010 214.060 100.795 ;
        RECT 215.000 100.200 216.830 100.880 ;
        RECT 216.840 100.200 218.670 100.880 ;
        RECT 215.485 99.970 216.830 100.200 ;
        RECT 217.325 99.970 218.670 100.200 ;
        RECT 219.620 99.970 220.510 100.920 ;
        RECT 221.855 100.880 222.025 101.070 ;
        RECT 225.720 100.880 225.890 101.070 ;
        RECT 227.100 100.900 227.270 101.090 ;
        RECT 229.400 100.880 229.570 101.070 ;
        RECT 230.135 100.880 230.305 101.070 ;
        RECT 234.000 100.880 234.170 101.070 ;
        RECT 237.680 100.900 237.850 101.090 ;
        RECT 238.135 100.930 238.255 101.040 ;
        RECT 238.600 100.900 238.770 101.090 ;
        RECT 240.900 100.880 241.070 101.070 ;
        RECT 241.360 100.880 241.530 101.070 ;
        RECT 243.195 100.930 243.315 101.040 ;
        RECT 250.100 100.900 250.270 101.090 ;
        RECT 251.480 100.900 251.650 101.090 ;
        RECT 251.935 100.930 252.055 101.040 ;
        RECT 252.400 100.880 252.570 101.070 ;
        RECT 252.870 100.925 253.030 101.035 ;
        RECT 253.780 100.880 253.950 101.070 ;
        RECT 254.240 100.900 254.410 101.090 ;
        RECT 254.710 100.935 254.870 101.045 ;
        RECT 255.620 100.900 255.790 101.090 ;
        RECT 257.000 100.880 257.170 101.070 ;
        RECT 258.845 100.880 259.015 101.090 ;
        RECT 262.520 101.040 262.690 101.090 ;
        RECT 262.515 100.930 262.690 101.040 ;
        RECT 262.520 100.900 262.690 100.930 ;
        RECT 262.980 100.900 263.150 101.070 ;
        RECT 263.000 100.880 263.150 100.900 ;
        RECT 265.740 100.880 265.910 101.070 ;
        RECT 267.120 100.900 267.290 101.090 ;
        RECT 267.580 100.900 267.750 101.090 ;
        RECT 271.260 100.880 271.430 101.070 ;
        RECT 277.700 100.900 277.870 101.090 ;
        RECT 280.460 100.880 280.630 101.070 ;
        RECT 281.840 100.880 282.010 101.070 ;
        RECT 282.025 100.900 282.195 101.090 ;
        RECT 284.140 100.900 284.310 101.090 ;
        RECT 284.595 100.930 284.715 101.040 ;
        RECT 285.060 100.900 285.230 101.090 ;
        RECT 291.510 100.925 291.670 101.035 ;
        RECT 292.420 100.880 292.590 101.070 ;
        RECT 302.355 100.880 302.525 101.070 ;
        RECT 303.460 100.900 303.630 101.090 ;
        RECT 304.380 100.900 304.550 101.090 ;
        RECT 306.220 100.880 306.390 101.070 ;
        RECT 307.140 100.900 307.310 101.090 ;
        RECT 308.060 100.880 308.230 101.070 ;
        RECT 310.820 100.880 310.990 101.090 ;
        RECT 221.440 100.200 225.340 100.880 ;
        RECT 221.440 99.970 222.370 100.200 ;
        RECT 225.580 100.070 228.330 100.880 ;
        RECT 228.340 100.100 229.710 100.880 ;
        RECT 229.720 100.200 233.620 100.880 ;
        RECT 229.720 99.970 230.650 100.200 ;
        RECT 233.860 100.070 239.370 100.880 ;
        RECT 239.390 100.010 239.820 100.795 ;
        RECT 239.840 100.100 241.210 100.880 ;
        RECT 241.220 100.070 243.050 100.880 ;
        RECT 243.520 100.200 252.710 100.880 ;
        RECT 243.520 99.970 244.440 100.200 ;
        RECT 247.270 99.980 248.200 100.200 ;
        RECT 253.640 99.970 256.850 100.880 ;
        RECT 256.860 100.070 258.690 100.880 ;
        RECT 258.700 99.970 262.355 100.880 ;
        RECT 263.000 100.060 264.930 100.880 ;
        RECT 263.980 99.970 264.930 100.060 ;
        RECT 265.150 100.010 265.580 100.795 ;
        RECT 265.600 100.070 271.110 100.880 ;
        RECT 271.120 100.200 280.310 100.880 ;
        RECT 275.630 99.980 276.560 100.200 ;
        RECT 279.390 99.970 280.310 100.200 ;
        RECT 280.320 100.100 281.690 100.880 ;
        RECT 281.700 100.200 290.890 100.880 ;
        RECT 286.210 99.980 287.140 100.200 ;
        RECT 289.970 99.970 290.890 100.200 ;
        RECT 290.910 100.010 291.340 100.795 ;
        RECT 292.280 100.200 301.890 100.880 ;
        RECT 296.790 99.980 297.720 100.200 ;
        RECT 300.550 99.970 301.890 100.200 ;
        RECT 301.940 100.200 305.840 100.880 ;
        RECT 306.080 100.200 307.910 100.880 ;
        RECT 307.920 100.200 309.750 100.880 ;
        RECT 301.940 99.970 302.870 100.200 ;
        RECT 306.565 99.970 307.910 100.200 ;
        RECT 308.405 99.970 309.750 100.200 ;
        RECT 309.760 100.070 311.130 100.880 ;
      LAYER nwell ;
        RECT 161.905 96.850 311.325 99.680 ;
      LAYER pwell ;
        RECT 162.100 95.650 163.470 96.460 ;
        RECT 163.480 95.650 168.990 96.460 ;
        RECT 169.920 95.650 171.290 96.430 ;
        RECT 171.300 95.650 172.670 96.430 ;
        RECT 172.680 95.650 174.050 96.430 ;
        RECT 174.990 95.735 175.420 96.520 ;
        RECT 175.440 96.330 176.370 96.560 ;
        RECT 175.440 95.650 179.340 96.330 ;
        RECT 179.580 95.650 183.250 96.460 ;
        RECT 187.770 96.330 188.700 96.550 ;
        RECT 191.530 96.330 192.870 96.560 ;
        RECT 183.260 95.650 192.870 96.330 ;
        RECT 192.920 95.650 194.290 96.430 ;
        RECT 194.300 95.650 195.670 96.460 ;
        RECT 195.680 96.330 196.610 96.560 ;
        RECT 195.680 95.650 199.580 96.330 ;
        RECT 200.750 95.735 201.180 96.520 ;
        RECT 201.200 95.650 203.950 96.560 ;
        RECT 207.620 96.330 208.550 96.560 ;
        RECT 204.650 95.650 208.550 96.330 ;
        RECT 208.560 95.650 211.310 96.560 ;
        RECT 211.320 95.650 214.990 96.460 ;
        RECT 215.920 95.650 217.290 96.430 ;
        RECT 218.220 95.650 221.430 96.560 ;
        RECT 221.440 95.650 224.650 96.560 ;
        RECT 224.660 95.650 226.490 96.460 ;
        RECT 226.510 95.735 226.940 96.520 ;
        RECT 226.960 95.650 230.170 96.560 ;
        RECT 230.180 95.650 233.850 96.460 ;
        RECT 234.780 95.650 237.990 96.560 ;
        RECT 238.000 95.650 241.655 96.560 ;
        RECT 241.680 95.650 247.190 96.460 ;
        RECT 247.200 95.650 250.870 96.460 ;
        RECT 250.880 95.650 252.250 96.460 ;
        RECT 252.270 95.735 252.700 96.520 ;
        RECT 252.720 95.650 254.550 96.460 ;
        RECT 254.560 95.650 257.770 96.560 ;
        RECT 257.780 95.650 261.435 96.560 ;
        RECT 261.460 95.650 264.670 96.560 ;
        RECT 266.485 96.360 267.430 96.560 ;
        RECT 264.680 95.680 267.430 96.360 ;
        RECT 162.240 95.440 162.410 95.650 ;
        RECT 163.620 95.460 163.790 95.650 ;
        RECT 165.920 95.440 166.090 95.630 ;
        RECT 166.380 95.440 166.550 95.630 ;
        RECT 168.215 95.490 168.335 95.600 ;
        RECT 168.680 95.440 168.850 95.630 ;
        RECT 169.150 95.495 169.310 95.605 ;
        RECT 170.980 95.460 171.150 95.650 ;
        RECT 172.360 95.460 172.530 95.650 ;
        RECT 173.740 95.460 173.910 95.650 ;
        RECT 174.210 95.495 174.370 95.605 ;
        RECT 175.855 95.460 176.025 95.650 ;
        RECT 177.880 95.440 178.050 95.630 ;
        RECT 179.720 95.460 179.890 95.650 ;
        RECT 183.400 95.440 183.570 95.650 ;
        RECT 187.080 95.440 187.250 95.630 ;
        RECT 187.535 95.490 187.655 95.600 ;
        RECT 188.735 95.440 188.905 95.630 ;
        RECT 193.520 95.440 193.690 95.630 ;
        RECT 193.980 95.440 194.150 95.650 ;
        RECT 194.440 95.460 194.610 95.650 ;
        RECT 196.095 95.460 196.265 95.650 ;
        RECT 199.500 95.440 199.670 95.630 ;
        RECT 199.970 95.495 200.130 95.605 ;
        RECT 201.340 95.460 201.510 95.650 ;
        RECT 202.260 95.440 202.430 95.630 ;
        RECT 202.720 95.440 202.890 95.630 ;
        RECT 204.095 95.490 204.215 95.600 ;
        RECT 207.965 95.460 208.135 95.650 ;
        RECT 208.240 95.440 208.410 95.630 ;
        RECT 208.700 95.460 208.870 95.650 ;
        RECT 211.460 95.460 211.630 95.650 ;
        RECT 214.220 95.440 214.390 95.630 ;
        RECT 215.150 95.495 215.310 95.605 ;
        RECT 216.060 95.460 216.230 95.650 ;
        RECT 216.985 95.440 217.155 95.630 ;
        RECT 217.450 95.495 217.610 95.605 ;
        RECT 218.360 95.460 218.530 95.650 ;
        RECT 162.100 94.630 163.470 95.440 ;
        RECT 163.490 94.760 166.230 95.440 ;
        RECT 166.240 94.630 168.070 95.440 ;
        RECT 168.540 94.760 177.730 95.440 ;
        RECT 173.050 94.540 173.980 94.760 ;
        RECT 176.810 94.530 177.730 94.760 ;
        RECT 177.740 94.630 183.250 95.440 ;
        RECT 183.260 94.630 186.010 95.440 ;
        RECT 186.020 94.660 187.390 95.440 ;
        RECT 187.870 94.570 188.300 95.355 ;
        RECT 188.320 94.760 192.220 95.440 ;
        RECT 188.320 94.530 189.250 94.760 ;
        RECT 192.460 94.660 193.830 95.440 ;
        RECT 193.840 94.630 199.350 95.440 ;
        RECT 199.360 94.630 201.190 95.440 ;
        RECT 201.200 94.660 202.570 95.440 ;
        RECT 202.580 94.630 208.090 95.440 ;
        RECT 208.100 94.630 213.610 95.440 ;
        RECT 213.630 94.570 214.060 95.355 ;
        RECT 214.080 94.630 216.830 95.440 ;
        RECT 216.840 94.530 220.495 95.440 ;
        RECT 220.655 95.410 220.825 95.630 ;
        RECT 224.340 95.460 224.510 95.650 ;
        RECT 224.800 95.460 224.970 95.650 ;
        RECT 226.175 95.440 226.345 95.630 ;
        RECT 221.855 95.410 222.810 95.440 ;
        RECT 220.530 94.730 222.810 95.410 ;
        RECT 221.855 94.530 222.810 94.730 ;
        RECT 222.820 94.530 226.490 95.440 ;
        RECT 226.645 95.410 226.815 95.630 ;
        RECT 227.100 95.460 227.270 95.650 ;
        RECT 229.400 95.440 229.570 95.630 ;
        RECT 230.320 95.460 230.490 95.650 ;
        RECT 234.010 95.495 234.170 95.605 ;
        RECT 234.920 95.460 235.090 95.650 ;
        RECT 235.845 95.440 236.015 95.630 ;
        RECT 238.145 95.460 238.315 95.650 ;
        RECT 239.985 95.440 240.155 95.630 ;
        RECT 241.820 95.460 241.990 95.650 ;
        RECT 246.420 95.440 246.590 95.630 ;
        RECT 246.880 95.440 247.050 95.630 ;
        RECT 247.340 95.460 247.510 95.650 ;
        RECT 251.020 95.460 251.190 95.650 ;
        RECT 252.400 95.440 252.570 95.630 ;
        RECT 252.860 95.460 253.030 95.650 ;
        RECT 254.700 95.460 254.870 95.650 ;
        RECT 257.925 95.440 258.095 95.650 ;
        RECT 261.600 95.440 261.770 95.650 ;
        RECT 264.825 95.600 264.995 95.680 ;
        RECT 266.485 95.650 267.430 95.680 ;
        RECT 267.440 95.650 272.950 96.460 ;
        RECT 273.420 95.650 274.790 96.430 ;
        RECT 274.800 95.650 277.550 96.460 ;
        RECT 278.030 95.735 278.460 96.520 ;
        RECT 278.480 96.330 279.410 96.560 ;
        RECT 282.620 96.330 283.550 96.560 ;
        RECT 286.760 96.330 287.690 96.560 ;
        RECT 291.820 96.330 292.750 96.560 ;
        RECT 299.620 96.330 300.550 96.560 ;
        RECT 278.480 95.650 282.380 96.330 ;
        RECT 282.620 95.650 286.520 96.330 ;
        RECT 286.760 95.650 290.660 96.330 ;
        RECT 291.820 95.650 295.720 96.330 ;
        RECT 296.650 95.650 300.550 96.330 ;
        RECT 300.560 95.650 301.930 96.430 ;
        RECT 301.940 95.650 303.310 96.430 ;
        RECT 303.790 95.735 304.220 96.520 ;
        RECT 304.240 95.650 307.910 96.460 ;
        RECT 308.405 96.330 309.750 96.560 ;
        RECT 307.920 95.650 309.750 96.330 ;
        RECT 309.760 95.650 311.130 96.460 ;
        RECT 264.815 95.490 264.995 95.600 ;
        RECT 264.825 95.460 264.995 95.490 ;
        RECT 265.740 95.440 265.910 95.630 ;
        RECT 267.580 95.460 267.750 95.650 ;
        RECT 271.260 95.440 271.430 95.630 ;
        RECT 273.095 95.490 273.215 95.600 ;
        RECT 274.480 95.460 274.650 95.650 ;
        RECT 274.940 95.460 275.110 95.650 ;
        RECT 276.790 95.485 276.950 95.595 ;
        RECT 277.695 95.490 277.815 95.600 ;
        RECT 278.895 95.460 279.065 95.650 ;
        RECT 280.000 95.440 280.170 95.630 ;
        RECT 282.760 95.440 282.930 95.630 ;
        RECT 283.035 95.460 283.205 95.650 ;
        RECT 284.140 95.440 284.310 95.630 ;
        RECT 284.600 95.440 284.770 95.630 ;
        RECT 287.175 95.460 287.345 95.650 ;
        RECT 288.280 95.440 288.450 95.630 ;
        RECT 289.660 95.440 289.830 95.630 ;
        RECT 291.050 95.495 291.210 95.605 ;
        RECT 292.235 95.460 292.405 95.650 ;
        RECT 296.095 95.490 296.215 95.600 ;
        RECT 299.965 95.460 300.135 95.650 ;
        RECT 300.240 95.440 300.410 95.630 ;
        RECT 300.700 95.440 300.870 95.650 ;
        RECT 303.000 95.460 303.170 95.650 ;
        RECT 303.455 95.490 303.575 95.600 ;
        RECT 304.380 95.460 304.550 95.650 ;
        RECT 308.060 95.460 308.230 95.650 ;
        RECT 310.820 95.440 310.990 95.650 ;
        RECT 228.305 95.410 229.250 95.440 ;
        RECT 226.500 94.730 229.250 95.410 ;
        RECT 228.305 94.530 229.250 94.730 ;
        RECT 229.260 94.630 234.770 95.440 ;
        RECT 235.700 94.530 239.355 95.440 ;
        RECT 239.390 94.570 239.820 95.355 ;
        RECT 239.840 94.530 243.495 95.440 ;
        RECT 243.520 94.530 246.730 95.440 ;
        RECT 246.740 94.630 252.250 95.440 ;
        RECT 252.260 94.630 257.770 95.440 ;
        RECT 257.780 94.530 261.435 95.440 ;
        RECT 261.460 94.530 264.670 95.440 ;
        RECT 265.150 94.570 265.580 95.355 ;
        RECT 265.600 94.630 271.110 95.440 ;
        RECT 271.120 94.630 276.630 95.440 ;
        RECT 277.560 94.530 280.310 95.440 ;
        RECT 280.320 94.530 283.070 95.440 ;
        RECT 283.080 94.660 284.450 95.440 ;
        RECT 284.460 94.630 288.130 95.440 ;
        RECT 288.140 94.630 289.510 95.440 ;
        RECT 289.520 94.660 290.890 95.440 ;
        RECT 290.910 94.570 291.340 95.355 ;
        RECT 291.360 94.760 300.550 95.440 ;
        RECT 300.560 94.760 309.750 95.440 ;
        RECT 291.360 94.530 292.280 94.760 ;
        RECT 295.110 94.540 296.040 94.760 ;
        RECT 305.070 94.540 306.000 94.760 ;
        RECT 308.830 94.530 309.750 94.760 ;
        RECT 309.760 94.630 311.130 95.440 ;
      LAYER nwell ;
        RECT 161.905 91.410 311.325 94.240 ;
      LAYER pwell ;
        RECT 162.100 90.210 163.470 91.020 ;
        RECT 163.480 90.210 165.310 91.020 ;
        RECT 169.830 90.890 170.760 91.110 ;
        RECT 173.590 90.890 174.930 91.120 ;
        RECT 165.320 90.210 174.930 90.890 ;
        RECT 174.990 90.295 175.420 91.080 ;
        RECT 175.440 90.890 176.370 91.120 ;
        RECT 175.440 90.210 179.340 90.890 ;
        RECT 179.580 90.210 183.250 91.020 ;
        RECT 186.920 90.890 187.850 91.120 ;
        RECT 183.950 90.210 187.850 90.890 ;
        RECT 188.780 90.890 189.710 91.120 ;
        RECT 193.840 90.890 194.770 91.120 ;
        RECT 188.780 90.210 192.680 90.890 ;
        RECT 193.840 90.210 197.740 90.890 ;
        RECT 197.990 90.210 200.730 90.890 ;
        RECT 200.750 90.295 201.180 91.080 ;
        RECT 201.200 90.210 202.570 91.020 ;
        RECT 202.580 90.890 203.510 91.120 ;
        RECT 202.580 90.210 206.480 90.890 ;
        RECT 206.720 90.210 209.470 91.120 ;
        RECT 209.480 90.210 212.230 91.020 ;
        RECT 162.240 90.000 162.410 90.210 ;
        RECT 163.620 90.000 163.790 90.210 ;
        RECT 165.000 90.000 165.170 90.190 ;
        RECT 165.460 90.020 165.630 90.210 ;
        RECT 166.380 90.000 166.550 90.190 ;
        RECT 175.855 90.020 176.025 90.210 ;
        RECT 176.040 90.000 176.210 90.190 ;
        RECT 179.720 90.020 179.890 90.210 ;
        RECT 183.395 90.050 183.515 90.160 ;
        RECT 185.710 90.045 185.870 90.155 ;
        RECT 187.265 90.020 187.435 90.210 ;
        RECT 187.540 90.000 187.710 90.190 ;
        RECT 188.010 90.055 188.170 90.165 ;
        RECT 189.195 90.020 189.365 90.210 ;
        RECT 189.380 90.000 189.550 90.190 ;
        RECT 189.840 90.000 190.010 90.190 ;
        RECT 193.070 90.055 193.230 90.165 ;
        RECT 194.255 90.020 194.425 90.210 ;
        RECT 199.050 90.045 199.210 90.155 ;
        RECT 199.960 90.000 200.130 90.190 ;
        RECT 200.420 90.020 200.590 90.210 ;
        RECT 201.340 90.000 201.510 90.210 ;
        RECT 202.995 90.020 203.165 90.210 ;
        RECT 206.860 90.020 207.030 90.210 ;
        RECT 209.620 90.020 209.790 90.210 ;
        RECT 211.000 90.000 211.170 90.190 ;
        RECT 212.700 90.170 213.590 91.120 ;
        RECT 216.615 90.890 217.750 91.120 ;
        RECT 214.540 90.210 217.750 90.890 ;
        RECT 217.760 90.210 219.590 91.020 ;
        RECT 219.600 90.890 220.735 91.120 ;
        RECT 219.600 90.210 222.810 90.890 ;
        RECT 212.375 90.050 212.495 90.160 ;
        RECT 212.850 90.045 213.010 90.155 ;
        RECT 213.300 90.020 213.470 90.170 ;
        RECT 213.770 90.055 213.930 90.165 ;
        RECT 214.220 90.000 214.390 90.190 ;
        RECT 214.680 90.020 214.850 90.210 ;
        RECT 217.900 90.020 218.070 90.210 ;
        RECT 220.660 90.000 220.830 90.190 ;
        RECT 222.500 90.000 222.670 90.210 ;
        RECT 223.760 90.170 224.650 91.120 ;
        RECT 224.660 90.210 226.490 91.020 ;
        RECT 226.510 90.295 226.940 91.080 ;
        RECT 226.960 90.920 227.910 91.120 ;
        RECT 229.240 90.920 230.170 91.120 ;
        RECT 226.960 90.440 230.170 90.920 ;
        RECT 226.960 90.240 230.025 90.440 ;
        RECT 226.960 90.210 227.895 90.240 ;
        RECT 222.970 90.055 223.130 90.165 ;
        RECT 223.880 90.020 224.050 90.170 ;
        RECT 224.800 90.020 224.970 90.210 ;
        RECT 227.100 90.000 227.270 90.190 ;
        RECT 227.560 90.000 227.730 90.190 ;
        RECT 229.855 90.020 230.025 90.240 ;
        RECT 230.180 90.210 235.690 91.020 ;
        RECT 235.700 90.210 237.530 91.020 ;
        RECT 240.740 90.890 241.670 91.120 ;
        RECT 243.015 90.920 243.970 91.120 ;
        RECT 238.000 90.210 241.670 90.890 ;
        RECT 241.690 90.240 243.970 90.920 ;
        RECT 230.320 90.020 230.490 90.210 ;
        RECT 233.080 90.000 233.250 90.190 ;
        RECT 235.840 90.160 236.010 90.210 ;
        RECT 235.835 90.050 236.010 90.160 ;
        RECT 237.675 90.050 237.795 90.160 ;
        RECT 235.840 90.020 236.010 90.050 ;
        RECT 238.140 90.020 238.310 90.210 ;
        RECT 239.070 90.000 239.240 90.190 ;
        RECT 239.980 90.020 240.150 90.190 ;
        RECT 241.815 90.020 241.985 90.240 ;
        RECT 243.015 90.210 243.970 90.240 ;
        RECT 243.980 90.210 249.490 91.020 ;
        RECT 249.500 90.210 252.250 91.020 ;
        RECT 252.270 90.295 252.700 91.080 ;
        RECT 252.720 90.210 258.230 91.020 ;
        RECT 258.700 90.210 261.910 91.120 ;
        RECT 261.920 90.210 267.430 91.020 ;
        RECT 267.440 90.210 272.950 91.020 ;
        RECT 272.960 90.210 276.630 91.020 ;
        RECT 276.640 90.210 278.010 90.990 ;
        RECT 278.030 90.295 278.460 91.080 ;
        RECT 278.480 90.890 279.410 91.120 ;
        RECT 278.480 90.210 282.380 90.890 ;
        RECT 282.620 90.210 283.990 90.990 ;
        RECT 284.000 90.210 289.510 91.020 ;
        RECT 289.980 90.890 290.910 91.120 ;
        RECT 289.980 90.210 293.880 90.890 ;
        RECT 294.120 90.210 295.950 91.020 ;
        RECT 299.160 90.890 300.090 91.120 ;
        RECT 296.190 90.210 300.090 90.890 ;
        RECT 300.100 90.210 301.470 90.990 ;
        RECT 301.480 90.210 303.310 91.020 ;
        RECT 303.790 90.295 304.220 91.080 ;
        RECT 304.240 90.210 309.750 91.020 ;
        RECT 309.760 90.210 311.130 91.020 ;
        RECT 239.990 90.000 240.150 90.020 ;
        RECT 244.120 90.000 244.290 90.210 ;
        RECT 249.640 90.000 249.810 90.210 ;
        RECT 252.860 90.020 253.030 90.210 ;
        RECT 253.315 90.050 253.435 90.160 ;
        RECT 256.550 90.000 256.720 90.190 ;
        RECT 257.005 90.000 257.175 90.190 ;
        RECT 258.375 90.050 258.495 90.160 ;
        RECT 258.830 90.020 259.000 90.210 ;
        RECT 260.685 90.000 260.855 90.190 ;
        RECT 262.060 90.020 262.230 90.210 ;
        RECT 264.370 90.045 264.530 90.155 ;
        RECT 265.740 90.020 265.910 90.190 ;
        RECT 267.580 90.020 267.750 90.210 ;
        RECT 265.745 90.000 265.910 90.020 ;
        RECT 268.040 90.000 268.210 90.190 ;
        RECT 273.100 90.020 273.270 90.210 ;
        RECT 274.480 90.000 274.650 90.190 ;
        RECT 274.940 90.000 275.110 90.190 ;
        RECT 277.700 90.020 277.870 90.210 ;
        RECT 278.895 90.020 279.065 90.210 ;
        RECT 282.760 90.020 282.930 90.210 ;
        RECT 284.140 90.020 284.310 90.210 ;
        RECT 284.415 90.000 284.585 90.190 ;
        RECT 288.280 90.000 288.450 90.190 ;
        RECT 289.660 90.160 289.830 90.190 ;
        RECT 289.655 90.050 289.830 90.160 ;
        RECT 289.660 90.000 289.830 90.050 ;
        RECT 290.395 90.020 290.565 90.210 ;
        RECT 291.500 90.000 291.670 90.190 ;
        RECT 294.260 90.020 294.430 90.210 ;
        RECT 299.505 90.020 299.675 90.210 ;
        RECT 300.240 90.020 300.410 90.210 ;
        RECT 300.700 90.000 300.870 90.190 ;
        RECT 301.620 90.020 301.790 90.210 ;
        RECT 303.455 90.050 303.575 90.160 ;
        RECT 304.380 90.020 304.550 90.210 ;
        RECT 310.820 90.000 310.990 90.210 ;
        RECT 162.100 89.190 163.470 90.000 ;
        RECT 163.480 89.190 164.850 90.000 ;
        RECT 164.860 89.220 166.230 90.000 ;
        RECT 166.240 89.320 175.850 90.000 ;
        RECT 175.900 89.320 185.510 90.000 ;
        RECT 170.750 89.100 171.680 89.320 ;
        RECT 174.510 89.090 175.850 89.320 ;
        RECT 180.410 89.100 181.340 89.320 ;
        RECT 184.170 89.090 185.510 89.320 ;
        RECT 186.480 89.220 187.850 90.000 ;
        RECT 187.870 89.130 188.300 89.915 ;
        RECT 188.320 89.220 189.690 90.000 ;
        RECT 189.700 89.320 198.890 90.000 ;
        RECT 194.210 89.100 195.140 89.320 ;
        RECT 197.970 89.090 198.890 89.320 ;
        RECT 199.820 89.220 201.190 90.000 ;
        RECT 201.200 89.320 210.810 90.000 ;
        RECT 210.860 89.320 212.690 90.000 ;
        RECT 205.710 89.100 206.640 89.320 ;
        RECT 209.470 89.090 210.810 89.320 ;
        RECT 211.345 89.090 212.690 89.320 ;
        RECT 213.630 89.130 214.060 89.915 ;
        RECT 214.080 89.190 217.750 90.000 ;
        RECT 218.690 89.090 222.810 90.000 ;
        RECT 222.830 89.960 223.750 90.000 ;
        RECT 222.820 89.770 223.750 89.960 ;
        RECT 225.840 89.770 227.410 90.000 ;
        RECT 222.820 89.410 227.410 89.770 ;
        RECT 222.830 89.320 227.410 89.410 ;
        RECT 222.830 89.090 225.830 89.320 ;
        RECT 227.420 89.190 232.930 90.000 ;
        RECT 232.940 89.190 235.690 90.000 ;
        RECT 236.160 89.090 239.370 90.000 ;
        RECT 239.390 89.130 239.820 89.915 ;
        RECT 239.990 89.090 243.645 90.000 ;
        RECT 243.980 89.190 249.490 90.000 ;
        RECT 249.500 89.190 253.170 90.000 ;
        RECT 253.640 89.090 256.850 90.000 ;
        RECT 256.860 89.090 260.530 90.000 ;
        RECT 260.540 89.090 264.210 90.000 ;
        RECT 265.150 89.130 265.580 89.915 ;
        RECT 265.745 89.320 267.580 90.000 ;
        RECT 266.650 89.090 267.580 89.320 ;
        RECT 267.900 89.190 269.730 90.000 ;
        RECT 269.975 89.320 274.790 90.000 ;
        RECT 274.800 89.320 283.990 90.000 ;
        RECT 279.310 89.100 280.240 89.320 ;
        RECT 283.070 89.090 283.990 89.320 ;
        RECT 284.000 89.320 287.900 90.000 ;
        RECT 284.000 89.090 284.930 89.320 ;
        RECT 288.140 89.190 289.510 90.000 ;
        RECT 289.520 89.220 290.890 90.000 ;
        RECT 290.910 89.130 291.340 89.915 ;
        RECT 291.360 89.320 300.550 90.000 ;
        RECT 300.560 89.320 309.750 90.000 ;
        RECT 295.870 89.100 296.800 89.320 ;
        RECT 299.630 89.090 300.550 89.320 ;
        RECT 305.070 89.100 306.000 89.320 ;
        RECT 308.830 89.090 309.750 89.320 ;
        RECT 309.760 89.190 311.130 90.000 ;
      LAYER nwell ;
        RECT 161.905 85.970 311.325 88.800 ;
      LAYER pwell ;
        RECT 162.100 84.770 163.470 85.580 ;
        RECT 163.480 84.770 168.990 85.580 ;
        RECT 169.460 84.770 170.830 85.550 ;
        RECT 170.840 85.450 171.770 85.680 ;
        RECT 170.840 84.770 174.740 85.450 ;
        RECT 174.990 84.855 175.420 85.640 ;
        RECT 175.440 85.450 176.370 85.680 ;
        RECT 175.440 84.770 179.340 85.450 ;
        RECT 179.580 84.770 183.250 85.580 ;
        RECT 188.690 85.450 189.620 85.670 ;
        RECT 192.450 85.450 193.790 85.680 ;
        RECT 184.180 84.770 193.790 85.450 ;
        RECT 193.840 84.770 199.350 85.580 ;
        RECT 199.360 84.770 200.730 85.580 ;
        RECT 200.750 84.855 201.180 85.640 ;
        RECT 201.200 84.770 203.950 85.680 ;
        RECT 204.420 84.770 206.250 85.450 ;
        RECT 206.260 84.770 208.030 85.680 ;
        RECT 208.110 85.590 209.700 85.680 ;
        RECT 208.110 84.770 210.680 85.590 ;
        RECT 210.860 84.770 212.690 85.450 ;
        RECT 212.700 84.770 218.210 85.580 ;
        RECT 218.220 84.770 220.050 85.580 ;
        RECT 220.520 84.770 226.090 85.680 ;
        RECT 226.510 84.855 226.940 85.640 ;
        RECT 226.960 84.770 232.470 85.580 ;
        RECT 232.940 84.770 236.830 85.680 ;
        RECT 237.080 84.770 238.450 85.580 ;
        RECT 238.460 84.770 242.130 85.680 ;
        RECT 243.190 85.450 244.120 85.680 ;
        RECT 242.285 84.770 244.120 85.450 ;
        RECT 244.440 84.770 249.950 85.580 ;
        RECT 249.960 84.770 251.790 85.580 ;
        RECT 252.270 84.855 252.700 85.640 ;
        RECT 252.720 84.770 255.470 85.580 ;
        RECT 255.940 84.770 259.150 85.680 ;
        RECT 259.770 84.770 263.425 85.680 ;
        RECT 263.910 84.770 267.565 85.680 ;
        RECT 268.095 84.770 271.570 85.680 ;
        RECT 271.580 84.770 277.090 85.580 ;
        RECT 278.030 84.855 278.460 85.640 ;
        RECT 278.480 84.770 281.230 85.680 ;
        RECT 281.240 84.770 283.070 85.580 ;
        RECT 287.590 85.450 288.520 85.670 ;
        RECT 291.350 85.450 292.690 85.680 ;
        RECT 283.080 84.770 292.690 85.450 ;
        RECT 293.200 84.770 294.570 85.550 ;
        RECT 298.240 85.450 299.170 85.680 ;
        RECT 295.270 84.770 299.170 85.450 ;
        RECT 299.180 84.770 300.550 85.550 ;
        RECT 300.560 84.770 303.310 85.580 ;
        RECT 303.790 84.855 304.220 85.640 ;
        RECT 304.240 84.770 307.910 85.580 ;
        RECT 308.380 84.770 309.750 85.550 ;
        RECT 309.760 84.770 311.130 85.580 ;
        RECT 162.240 84.560 162.410 84.770 ;
        RECT 163.620 84.560 163.790 84.770 ;
        RECT 169.140 84.720 169.310 84.750 ;
        RECT 169.135 84.610 169.310 84.720 ;
        RECT 169.140 84.560 169.310 84.610 ;
        RECT 169.600 84.580 169.770 84.770 ;
        RECT 171.255 84.580 171.425 84.770 ;
        RECT 174.660 84.560 174.830 84.750 ;
        RECT 175.855 84.580 176.025 84.770 ;
        RECT 179.720 84.580 179.890 84.770 ;
        RECT 183.410 84.615 183.570 84.725 ;
        RECT 184.320 84.580 184.490 84.770 ;
        RECT 187.540 84.560 187.710 84.750 ;
        RECT 188.470 84.605 188.630 84.715 ;
        RECT 190.300 84.560 190.470 84.750 ;
        RECT 190.770 84.605 190.930 84.715 ;
        RECT 193.980 84.580 194.150 84.770 ;
        RECT 196.280 84.560 196.450 84.750 ;
        RECT 196.740 84.560 196.910 84.750 ;
        RECT 199.500 84.580 199.670 84.770 ;
        RECT 200.420 84.560 200.590 84.750 ;
        RECT 201.340 84.580 201.510 84.770 ;
        RECT 201.800 84.560 201.970 84.750 ;
        RECT 204.095 84.610 204.215 84.720 ;
        RECT 204.560 84.580 204.730 84.770 ;
        RECT 206.405 84.580 206.575 84.770 ;
        RECT 210.540 84.750 210.680 84.770 ;
        RECT 206.855 84.610 206.975 84.720 ;
        RECT 209.620 84.580 209.790 84.750 ;
        RECT 210.075 84.610 210.195 84.720 ;
        RECT 210.540 84.580 210.710 84.750 ;
        RECT 211.000 84.580 211.170 84.770 ;
        RECT 212.840 84.580 213.010 84.770 ;
        RECT 213.295 84.610 213.415 84.720 ;
        RECT 209.620 84.560 209.760 84.580 ;
        RECT 212.840 84.560 212.980 84.580 ;
        RECT 214.220 84.560 214.390 84.750 ;
        RECT 218.360 84.580 218.530 84.770 ;
        RECT 220.205 84.720 220.375 84.750 ;
        RECT 219.735 84.610 219.855 84.720 ;
        RECT 220.195 84.610 220.375 84.720 ;
        RECT 220.205 84.560 220.375 84.610 ;
        RECT 220.665 84.580 220.835 84.770 ;
        RECT 162.100 83.750 163.470 84.560 ;
        RECT 163.480 83.750 168.990 84.560 ;
        RECT 169.000 83.750 174.510 84.560 ;
        RECT 174.520 83.750 178.190 84.560 ;
        RECT 178.240 83.880 187.850 84.560 ;
        RECT 178.240 83.650 179.580 83.880 ;
        RECT 182.410 83.660 183.340 83.880 ;
        RECT 187.870 83.690 188.300 84.475 ;
        RECT 189.240 83.780 190.610 84.560 ;
        RECT 191.775 83.880 196.590 84.560 ;
        RECT 196.600 83.750 200.270 84.560 ;
        RECT 200.280 83.750 201.650 84.560 ;
        RECT 201.660 83.880 206.475 84.560 ;
        RECT 207.190 83.740 209.760 84.560 ;
        RECT 210.410 83.740 212.980 84.560 ;
        RECT 207.190 83.650 208.780 83.740 ;
        RECT 210.410 83.650 212.000 83.740 ;
        RECT 213.630 83.690 214.060 84.475 ;
        RECT 214.080 83.750 219.590 84.560 ;
        RECT 220.060 83.650 226.570 84.560 ;
        RECT 227.100 84.530 227.270 84.770 ;
        RECT 229.860 84.560 230.030 84.750 ;
        RECT 232.620 84.720 232.790 84.750 ;
        RECT 232.615 84.610 232.790 84.720 ;
        RECT 232.620 84.560 232.790 84.610 ;
        RECT 233.085 84.580 233.255 84.770 ;
        RECT 237.220 84.580 237.390 84.770 ;
        RECT 238.140 84.560 238.310 84.750 ;
        RECT 238.605 84.580 238.775 84.770 ;
        RECT 242.285 84.750 242.450 84.770 ;
        RECT 239.980 84.560 240.150 84.750 ;
        RECT 241.815 84.610 241.935 84.720 ;
        RECT 242.280 84.580 242.455 84.750 ;
        RECT 244.580 84.580 244.750 84.770 ;
        RECT 242.285 84.560 242.455 84.580 ;
        RECT 245.965 84.560 246.135 84.750 ;
        RECT 249.180 84.560 249.350 84.750 ;
        RECT 250.100 84.580 250.270 84.770 ;
        RECT 251.935 84.610 252.055 84.720 ;
        RECT 252.860 84.580 253.030 84.770 ;
        RECT 254.700 84.560 254.870 84.750 ;
        RECT 255.615 84.610 255.735 84.720 ;
        RECT 258.850 84.580 259.020 84.770 ;
        RECT 259.770 84.750 259.930 84.770 ;
        RECT 263.910 84.750 264.070 84.770 ;
        RECT 259.295 84.610 259.415 84.720 ;
        RECT 259.760 84.580 259.930 84.750 ;
        RECT 260.220 84.560 260.390 84.750 ;
        RECT 263.900 84.580 264.070 84.750 ;
        RECT 264.815 84.560 264.985 84.750 ;
        RECT 265.740 84.580 265.910 84.750 ;
        RECT 265.745 84.560 265.910 84.580 ;
        RECT 268.040 84.560 268.210 84.750 ;
        RECT 271.255 84.580 271.425 84.770 ;
        RECT 271.720 84.560 271.890 84.770 ;
        RECT 273.100 84.560 273.270 84.750 ;
        RECT 277.250 84.615 277.410 84.725 ;
        RECT 280.920 84.580 281.090 84.770 ;
        RECT 281.380 84.580 281.550 84.770 ;
        RECT 282.300 84.560 282.470 84.750 ;
        RECT 283.220 84.580 283.390 84.770 ;
        RECT 288.280 84.560 288.450 84.750 ;
        RECT 288.740 84.560 288.910 84.750 ;
        RECT 290.575 84.610 290.695 84.720 ;
        RECT 291.510 84.605 291.670 84.715 ;
        RECT 292.875 84.610 292.995 84.720 ;
        RECT 293.340 84.580 293.510 84.770 ;
        RECT 294.720 84.720 294.890 84.750 ;
        RECT 294.715 84.610 294.890 84.720 ;
        RECT 295.175 84.610 295.295 84.720 ;
        RECT 294.720 84.560 294.890 84.610 ;
        RECT 295.915 84.560 296.085 84.750 ;
        RECT 298.585 84.580 298.755 84.770 ;
        RECT 299.320 84.580 299.490 84.770 ;
        RECT 299.780 84.560 299.950 84.750 ;
        RECT 300.700 84.580 300.870 84.770 ;
        RECT 303.455 84.610 303.575 84.720 ;
        RECT 304.380 84.580 304.550 84.770 ;
        RECT 309.440 84.720 309.610 84.770 ;
        RECT 308.055 84.610 308.175 84.720 ;
        RECT 309.435 84.610 309.610 84.720 ;
        RECT 309.440 84.580 309.610 84.610 ;
        RECT 310.820 84.560 310.990 84.770 ;
        RECT 228.315 84.530 229.710 84.560 ;
        RECT 226.975 83.850 229.710 84.530 ;
        RECT 229.720 83.880 232.460 84.560 ;
        RECT 228.300 83.650 229.710 83.850 ;
        RECT 232.480 83.750 237.990 84.560 ;
        RECT 238.000 83.750 239.370 84.560 ;
        RECT 239.390 83.690 239.820 84.475 ;
        RECT 239.840 83.750 241.670 84.560 ;
        RECT 242.140 83.650 245.795 84.560 ;
        RECT 245.820 83.650 248.740 84.560 ;
        RECT 249.040 83.750 254.550 84.560 ;
        RECT 254.560 83.750 260.070 84.560 ;
        RECT 260.080 83.750 261.910 84.560 ;
        RECT 262.210 83.650 265.130 84.560 ;
        RECT 265.150 83.690 265.580 84.475 ;
        RECT 265.745 83.880 267.580 84.560 ;
        RECT 266.650 83.650 267.580 83.880 ;
        RECT 267.900 83.750 271.570 84.560 ;
        RECT 271.580 83.750 272.950 84.560 ;
        RECT 272.960 83.880 282.150 84.560 ;
        RECT 282.160 83.880 286.975 84.560 ;
        RECT 277.470 83.660 278.400 83.880 ;
        RECT 281.230 83.650 282.150 83.880 ;
        RECT 287.220 83.780 288.590 84.560 ;
        RECT 288.600 83.750 290.430 84.560 ;
        RECT 290.910 83.690 291.340 84.475 ;
        RECT 292.290 83.880 295.030 84.560 ;
        RECT 295.500 83.880 299.400 84.560 ;
        RECT 299.640 83.880 309.250 84.560 ;
        RECT 295.500 83.650 296.430 83.880 ;
        RECT 304.150 83.660 305.080 83.880 ;
        RECT 307.910 83.650 309.250 83.880 ;
        RECT 309.760 83.750 311.130 84.560 ;
      LAYER nwell ;
        RECT 161.905 80.530 311.325 83.360 ;
      LAYER pwell ;
        RECT 162.100 79.330 163.470 80.140 ;
        RECT 163.480 79.330 168.990 80.140 ;
        RECT 169.460 79.330 170.830 80.110 ;
        RECT 170.840 79.330 172.210 80.110 ;
        RECT 173.140 79.330 174.510 80.110 ;
        RECT 174.990 79.415 175.420 80.200 ;
        RECT 175.440 80.010 176.370 80.240 ;
        RECT 175.440 79.330 179.340 80.010 ;
        RECT 179.580 79.330 185.090 80.140 ;
        RECT 185.560 79.330 186.930 80.110 ;
        RECT 191.450 80.010 192.380 80.230 ;
        RECT 195.210 80.010 196.130 80.240 ;
        RECT 186.940 79.330 196.130 80.010 ;
        RECT 196.140 79.330 199.810 80.140 ;
        RECT 200.750 79.415 201.180 80.200 ;
        RECT 207.650 80.150 209.240 80.240 ;
        RECT 201.200 79.330 206.710 80.140 ;
        RECT 207.650 79.330 210.220 80.150 ;
        RECT 210.400 79.330 215.910 80.140 ;
        RECT 215.920 79.330 218.670 80.140 ;
        RECT 219.210 79.560 223.560 80.240 ;
        RECT 219.790 79.330 223.560 79.560 ;
        RECT 223.740 79.330 226.490 80.140 ;
        RECT 226.510 79.415 226.940 80.200 ;
        RECT 226.960 79.330 230.170 80.240 ;
        RECT 230.180 79.330 235.690 80.140 ;
        RECT 236.620 79.330 239.830 80.240 ;
        RECT 239.840 79.330 243.495 80.240 ;
        RECT 243.520 79.330 247.175 80.240 ;
        RECT 247.200 79.330 250.870 80.140 ;
        RECT 250.880 79.330 252.250 80.140 ;
        RECT 252.270 79.415 252.700 80.200 ;
        RECT 252.720 79.330 258.230 80.140 ;
        RECT 258.240 79.330 261.450 80.240 ;
        RECT 261.460 79.330 266.970 80.140 ;
        RECT 266.980 79.330 272.490 80.140 ;
        RECT 272.500 79.330 273.870 80.140 ;
        RECT 273.880 79.330 275.250 80.110 ;
        RECT 275.260 79.330 276.630 80.110 ;
        RECT 276.640 79.330 278.010 80.140 ;
        RECT 278.030 79.415 278.460 80.200 ;
        RECT 278.480 79.330 283.990 80.140 ;
        RECT 289.430 80.010 290.360 80.230 ;
        RECT 293.190 80.010 294.530 80.240 ;
        RECT 284.920 79.330 294.530 80.010 ;
        RECT 294.580 80.010 295.510 80.240 ;
        RECT 298.720 80.010 299.650 80.240 ;
        RECT 294.580 79.330 298.480 80.010 ;
        RECT 298.720 79.330 302.620 80.010 ;
        RECT 303.790 79.415 304.220 80.200 ;
        RECT 304.240 79.330 305.610 80.110 ;
        RECT 305.620 79.330 309.290 80.140 ;
        RECT 309.760 79.330 311.130 80.140 ;
        RECT 162.240 79.120 162.410 79.330 ;
        RECT 163.620 79.120 163.790 79.330 ;
        RECT 167.310 79.165 167.470 79.275 ;
        RECT 168.220 79.120 168.390 79.310 ;
        RECT 169.135 79.170 169.255 79.280 ;
        RECT 170.520 79.140 170.690 79.330 ;
        RECT 171.900 79.140 172.070 79.330 ;
        RECT 172.370 79.175 172.530 79.285 ;
        RECT 173.280 79.140 173.450 79.330 ;
        RECT 174.655 79.170 174.775 79.280 ;
        RECT 175.855 79.140 176.025 79.330 ;
        RECT 177.880 79.120 178.050 79.310 ;
        RECT 179.720 79.140 179.890 79.330 ;
        RECT 185.235 79.170 185.355 79.280 ;
        RECT 185.700 79.140 185.870 79.330 ;
        RECT 187.080 79.140 187.250 79.330 ;
        RECT 187.535 79.170 187.655 79.280 ;
        RECT 188.460 79.120 188.630 79.310 ;
        RECT 196.280 79.140 196.450 79.330 ;
        RECT 198.395 79.120 198.565 79.310 ;
        RECT 199.970 79.175 200.130 79.285 ;
        RECT 201.340 79.140 201.510 79.330 ;
        RECT 210.080 79.310 210.220 79.330 ;
        RECT 202.260 79.120 202.430 79.310 ;
        RECT 205.940 79.120 206.110 79.310 ;
        RECT 206.870 79.175 207.030 79.285 ;
        RECT 209.160 79.120 209.330 79.310 ;
        RECT 210.080 79.140 210.250 79.310 ;
        RECT 210.540 79.140 210.710 79.330 ;
        RECT 211.000 79.120 211.170 79.310 ;
        RECT 214.220 79.120 214.390 79.310 ;
        RECT 216.060 79.140 216.230 79.330 ;
        RECT 223.420 79.310 223.560 79.330 ;
        RECT 223.880 79.310 224.050 79.330 ;
        RECT 218.825 79.280 218.995 79.310 ;
        RECT 217.910 79.165 218.070 79.275 ;
        RECT 218.815 79.170 218.995 79.280 ;
        RECT 218.825 79.120 218.995 79.170 ;
        RECT 222.500 79.120 222.670 79.310 ;
        RECT 223.420 79.140 223.590 79.310 ;
        RECT 223.880 79.140 224.055 79.310 ;
        RECT 223.885 79.120 224.055 79.140 ;
        RECT 227.565 79.120 227.735 79.310 ;
        RECT 229.860 79.120 230.030 79.330 ;
        RECT 230.320 79.140 230.490 79.330 ;
        RECT 235.375 79.170 235.495 79.280 ;
        RECT 235.840 79.120 236.010 79.310 ;
        RECT 236.760 79.140 236.930 79.330 ;
        RECT 239.985 79.120 240.155 79.330 ;
        RECT 243.665 79.310 243.835 79.330 ;
        RECT 243.660 79.140 243.835 79.310 ;
        RECT 243.660 79.120 243.830 79.140 ;
        RECT 162.100 78.310 163.470 79.120 ;
        RECT 163.480 78.310 167.150 79.120 ;
        RECT 168.080 78.440 177.690 79.120 ;
        RECT 177.740 78.440 187.350 79.120 ;
        RECT 172.590 78.220 173.520 78.440 ;
        RECT 176.350 78.210 177.690 78.440 ;
        RECT 182.250 78.220 183.180 78.440 ;
        RECT 186.010 78.210 187.350 78.440 ;
        RECT 187.870 78.250 188.300 79.035 ;
        RECT 188.320 78.440 197.930 79.120 ;
        RECT 192.830 78.220 193.760 78.440 ;
        RECT 196.590 78.210 197.930 78.440 ;
        RECT 197.980 78.440 201.880 79.120 ;
        RECT 197.980 78.210 198.910 78.440 ;
        RECT 202.120 78.310 205.790 79.120 ;
        RECT 205.800 78.440 209.010 79.120 ;
        RECT 209.020 78.440 210.850 79.120 ;
        RECT 207.875 78.210 209.010 78.440 ;
        RECT 210.860 78.310 213.610 79.120 ;
        RECT 213.630 78.250 214.060 79.035 ;
        RECT 214.080 78.310 217.750 79.120 ;
        RECT 218.680 78.210 222.335 79.120 ;
        RECT 222.360 78.310 223.730 79.120 ;
        RECT 223.740 78.210 227.395 79.120 ;
        RECT 227.420 78.210 229.630 79.120 ;
        RECT 229.720 78.310 235.230 79.120 ;
        RECT 235.700 78.440 239.370 79.120 ;
        RECT 238.440 78.210 239.370 78.440 ;
        RECT 239.390 78.250 239.820 79.035 ;
        RECT 239.840 78.210 243.495 79.120 ;
        RECT 243.520 78.210 246.730 79.120 ;
        RECT 246.875 79.090 247.045 79.310 ;
        RECT 247.340 79.140 247.510 79.330 ;
        RECT 249.180 79.120 249.350 79.310 ;
        RECT 251.020 79.140 251.190 79.330 ;
        RECT 252.860 79.140 253.030 79.330 ;
        RECT 254.700 79.120 254.870 79.310 ;
        RECT 256.545 79.120 256.715 79.310 ;
        RECT 260.225 79.120 260.395 79.310 ;
        RECT 261.140 79.140 261.310 79.330 ;
        RECT 261.600 79.140 261.770 79.330 ;
        RECT 263.900 79.120 264.070 79.310 ;
        RECT 265.740 79.120 265.910 79.310 ;
        RECT 267.120 79.140 267.290 79.330 ;
        RECT 271.260 79.120 271.430 79.310 ;
        RECT 272.640 79.120 272.810 79.330 ;
        RECT 274.940 79.140 275.110 79.330 ;
        RECT 276.320 79.140 276.490 79.330 ;
        RECT 276.780 79.140 276.950 79.330 ;
        RECT 278.620 79.140 278.790 79.330 ;
        RECT 282.300 79.120 282.470 79.310 ;
        RECT 284.150 79.175 284.310 79.285 ;
        RECT 285.060 79.140 285.230 79.330 ;
        RECT 285.980 79.120 286.150 79.310 ;
        RECT 291.500 79.120 291.670 79.310 ;
        RECT 294.255 79.170 294.375 79.280 ;
        RECT 294.720 79.120 294.890 79.310 ;
        RECT 294.995 79.140 295.165 79.330 ;
        RECT 299.135 79.140 299.305 79.330 ;
        RECT 303.010 79.175 303.170 79.285 ;
        RECT 304.380 79.120 304.550 79.310 ;
        RECT 305.300 79.140 305.470 79.330 ;
        RECT 305.760 79.140 305.930 79.330 ;
        RECT 309.435 79.170 309.555 79.280 ;
        RECT 310.820 79.120 310.990 79.330 ;
        RECT 248.075 79.090 249.030 79.120 ;
        RECT 246.750 78.410 249.030 79.090 ;
        RECT 248.075 78.210 249.030 78.410 ;
        RECT 249.040 78.310 254.550 79.120 ;
        RECT 254.560 78.310 256.390 79.120 ;
        RECT 256.400 78.210 260.055 79.120 ;
        RECT 260.080 78.210 263.735 79.120 ;
        RECT 263.760 78.310 265.130 79.120 ;
        RECT 265.150 78.250 265.580 79.035 ;
        RECT 265.600 78.310 271.110 79.120 ;
        RECT 271.120 78.310 272.490 79.120 ;
        RECT 272.500 78.440 282.110 79.120 ;
        RECT 277.010 78.220 277.940 78.440 ;
        RECT 280.770 78.210 282.110 78.440 ;
        RECT 282.160 78.310 285.830 79.120 ;
        RECT 285.840 78.440 290.655 79.120 ;
        RECT 290.910 78.250 291.340 79.035 ;
        RECT 291.360 78.310 294.110 79.120 ;
        RECT 294.580 78.440 304.190 79.120 ;
        RECT 299.090 78.220 300.020 78.440 ;
        RECT 302.850 78.210 304.190 78.440 ;
        RECT 304.240 78.310 309.750 79.120 ;
        RECT 309.760 78.310 311.130 79.120 ;
      LAYER nwell ;
        RECT 161.905 75.090 311.325 77.920 ;
      LAYER pwell ;
        RECT 162.100 73.890 163.470 74.700 ;
        RECT 163.480 73.890 165.310 74.700 ;
        RECT 169.830 74.570 170.760 74.790 ;
        RECT 173.590 74.570 174.930 74.800 ;
        RECT 165.320 73.890 174.930 74.570 ;
        RECT 174.990 73.975 175.420 74.760 ;
        RECT 175.900 74.570 176.830 74.800 ;
        RECT 190.070 74.570 191.000 74.790 ;
        RECT 193.830 74.570 195.170 74.800 ;
        RECT 175.900 73.890 179.800 74.570 ;
        RECT 180.735 73.890 185.550 74.570 ;
        RECT 185.560 73.890 195.170 74.570 ;
        RECT 195.220 74.570 196.150 74.800 ;
        RECT 195.220 73.890 199.120 74.570 ;
        RECT 199.360 73.890 200.730 74.670 ;
        RECT 200.750 73.975 201.180 74.760 ;
        RECT 201.200 73.890 203.940 74.570 ;
        RECT 203.960 73.890 206.710 74.700 ;
        RECT 206.720 73.890 210.375 74.800 ;
        RECT 210.400 73.890 214.070 74.700 ;
        RECT 162.240 73.680 162.410 73.890 ;
        RECT 163.620 73.680 163.790 73.890 ;
        RECT 165.460 73.700 165.630 73.890 ;
        RECT 169.150 73.725 169.310 73.835 ;
        RECT 170.980 73.680 171.150 73.870 ;
        RECT 171.440 73.680 171.610 73.870 ;
        RECT 173.555 73.680 173.725 73.870 ;
        RECT 175.575 73.730 175.695 73.840 ;
        RECT 176.315 73.700 176.485 73.890 ;
        RECT 177.695 73.680 177.865 73.870 ;
        RECT 180.175 73.730 180.295 73.840 ;
        RECT 181.560 73.680 181.730 73.870 ;
        RECT 183.395 73.730 183.515 73.840 ;
        RECT 185.240 73.700 185.410 73.890 ;
        RECT 185.700 73.700 185.870 73.890 ;
        RECT 187.265 73.680 187.435 73.870 ;
        RECT 193.060 73.680 193.230 73.870 ;
        RECT 193.515 73.730 193.635 73.840 ;
        RECT 193.980 73.680 194.150 73.870 ;
        RECT 195.635 73.700 195.805 73.890 ;
        RECT 200.420 73.700 200.590 73.890 ;
        RECT 201.340 73.700 201.510 73.890 ;
        RECT 203.640 73.680 203.810 73.870 ;
        RECT 204.100 73.700 204.270 73.890 ;
        RECT 206.400 73.680 206.570 73.870 ;
        RECT 206.865 73.700 207.035 73.890 ;
        RECT 210.540 73.700 210.710 73.890 ;
        RECT 211.920 73.680 212.090 73.870 ;
        RECT 214.080 73.850 214.970 74.800 ;
        RECT 218.660 74.570 219.590 74.800 ;
        RECT 215.920 73.890 219.590 74.570 ;
        RECT 219.600 73.890 226.110 74.800 ;
        RECT 226.510 73.975 226.940 74.760 ;
        RECT 228.295 74.600 229.250 74.800 ;
        RECT 226.970 73.920 229.250 74.600 ;
        RECT 214.220 73.680 214.390 73.850 ;
        RECT 214.680 73.700 214.850 73.850 ;
        RECT 215.150 73.735 215.310 73.845 ;
        RECT 216.060 73.700 216.230 73.890 ;
        RECT 219.745 73.700 219.915 73.890 ;
        RECT 162.100 72.870 163.470 73.680 ;
        RECT 163.480 72.870 168.990 73.680 ;
        RECT 169.920 72.900 171.290 73.680 ;
        RECT 171.300 72.870 173.130 73.680 ;
        RECT 173.140 73.000 177.040 73.680 ;
        RECT 177.280 73.000 181.180 73.680 ;
        RECT 173.140 72.770 174.070 73.000 ;
        RECT 177.280 72.770 178.210 73.000 ;
        RECT 181.420 72.870 183.250 73.680 ;
        RECT 183.950 73.000 187.850 73.680 ;
        RECT 186.920 72.770 187.850 73.000 ;
        RECT 187.870 72.810 188.300 73.595 ;
        RECT 188.555 73.000 193.370 73.680 ;
        RECT 193.840 73.000 203.450 73.680 ;
        RECT 198.350 72.780 199.280 73.000 ;
        RECT 202.110 72.770 203.450 73.000 ;
        RECT 203.500 72.770 206.250 73.680 ;
        RECT 206.260 72.870 211.770 73.680 ;
        RECT 211.780 72.870 213.610 73.680 ;
        RECT 213.630 72.810 214.060 73.595 ;
        RECT 214.080 72.870 219.590 73.680 ;
        RECT 220.660 73.650 220.830 73.870 ;
        RECT 224.340 73.680 224.510 73.870 ;
        RECT 227.095 73.700 227.265 73.920 ;
        RECT 228.295 73.890 229.250 73.920 ;
        RECT 229.260 73.890 232.930 74.700 ;
        RECT 236.600 74.570 237.530 74.800 ;
        RECT 233.860 73.890 237.530 74.570 ;
        RECT 237.540 73.890 241.210 74.700 ;
        RECT 243.475 74.600 244.430 74.800 ;
        RECT 242.150 73.920 244.430 74.600 ;
        RECT 229.400 73.700 229.570 73.890 ;
        RECT 229.860 73.680 230.030 73.870 ;
        RECT 233.090 73.735 233.250 73.845 ;
        RECT 234.000 73.700 234.170 73.890 ;
        RECT 235.380 73.680 235.550 73.870 ;
        RECT 237.680 73.700 237.850 73.890 ;
        RECT 239.055 73.730 239.175 73.840 ;
        RECT 239.985 73.680 240.155 73.870 ;
        RECT 241.370 73.735 241.530 73.845 ;
        RECT 242.275 73.700 242.445 73.920 ;
        RECT 243.475 73.890 244.430 73.920 ;
        RECT 244.440 73.890 249.950 74.700 ;
        RECT 249.960 73.890 251.790 74.700 ;
        RECT 252.270 73.975 252.700 74.760 ;
        RECT 252.720 73.890 256.390 74.700 ;
        RECT 257.320 73.890 260.530 74.800 ;
        RECT 261.875 74.600 262.830 74.800 ;
        RECT 264.175 74.600 265.130 74.800 ;
        RECT 260.550 73.920 262.830 74.600 ;
        RECT 262.850 73.920 265.130 74.600 ;
        RECT 243.660 73.680 243.830 73.870 ;
        RECT 244.580 73.700 244.750 73.890 ;
        RECT 249.180 73.680 249.350 73.870 ;
        RECT 250.100 73.700 250.270 73.890 ;
        RECT 251.935 73.730 252.055 73.840 ;
        RECT 252.860 73.700 253.030 73.890 ;
        RECT 254.695 73.730 254.815 73.840 ;
        RECT 255.165 73.680 255.335 73.870 ;
        RECT 256.550 73.735 256.710 73.845 ;
        RECT 257.460 73.700 257.630 73.890 ;
        RECT 258.840 73.680 259.010 73.870 ;
        RECT 260.675 73.700 260.845 73.920 ;
        RECT 261.875 73.890 262.830 73.920 ;
        RECT 262.975 73.700 263.145 73.920 ;
        RECT 264.175 73.890 265.130 73.920 ;
        RECT 265.140 73.890 270.650 74.700 ;
        RECT 270.660 73.890 273.410 74.700 ;
        RECT 273.880 74.570 274.810 74.800 ;
        RECT 273.880 73.890 277.780 74.570 ;
        RECT 278.030 73.975 278.460 74.760 ;
        RECT 278.480 74.570 279.410 74.800 ;
        RECT 278.480 73.890 282.380 74.570 ;
        RECT 282.620 73.890 284.450 74.700 ;
        RECT 284.920 73.890 286.290 74.670 ;
        RECT 286.300 74.570 287.220 74.800 ;
        RECT 290.050 74.570 290.980 74.790 ;
        RECT 299.160 74.570 300.090 74.800 ;
        RECT 286.300 73.890 295.490 74.570 ;
        RECT 296.190 73.890 300.090 74.570 ;
        RECT 300.100 73.890 301.470 74.670 ;
        RECT 301.480 73.890 303.310 74.700 ;
        RECT 303.790 73.975 304.220 74.760 ;
        RECT 304.240 74.570 305.170 74.800 ;
        RECT 304.240 73.890 308.140 74.570 ;
        RECT 308.380 73.890 309.750 74.700 ;
        RECT 309.760 73.890 311.130 74.700 ;
        RECT 264.370 73.725 264.530 73.835 ;
        RECT 265.280 73.700 265.450 73.890 ;
        RECT 265.740 73.680 265.910 73.870 ;
        RECT 270.800 73.700 270.970 73.890 ;
        RECT 271.260 73.680 271.430 73.870 ;
        RECT 273.555 73.730 273.675 73.840 ;
        RECT 274.295 73.700 274.465 73.890 ;
        RECT 276.780 73.680 276.950 73.870 ;
        RECT 278.895 73.700 279.065 73.890 ;
        RECT 280.920 73.680 281.090 73.870 ;
        RECT 281.380 73.680 281.550 73.870 ;
        RECT 282.760 73.700 282.930 73.890 ;
        RECT 284.595 73.730 284.715 73.840 ;
        RECT 285.060 73.700 285.230 73.890 ;
        RECT 285.980 73.680 286.150 73.870 ;
        RECT 291.500 73.680 291.670 73.870 ;
        RECT 293.335 73.730 293.455 73.840 ;
        RECT 293.800 73.680 293.970 73.870 ;
        RECT 295.180 73.680 295.350 73.890 ;
        RECT 295.635 73.730 295.755 73.840 ;
        RECT 299.505 73.700 299.675 73.890 ;
        RECT 301.160 73.700 301.330 73.890 ;
        RECT 301.620 73.700 301.790 73.890 ;
        RECT 303.455 73.730 303.575 73.840 ;
        RECT 304.655 73.700 304.825 73.890 ;
        RECT 304.840 73.680 305.010 73.870 ;
        RECT 308.520 73.680 308.690 73.890 ;
        RECT 310.820 73.680 310.990 73.890 ;
        RECT 222.820 73.650 224.190 73.680 ;
        RECT 220.520 72.970 224.190 73.650 ;
        RECT 222.805 72.770 224.190 72.970 ;
        RECT 224.200 72.870 229.710 73.680 ;
        RECT 229.720 72.870 235.230 73.680 ;
        RECT 235.240 72.870 238.910 73.680 ;
        RECT 239.390 72.810 239.820 73.595 ;
        RECT 239.840 72.770 243.495 73.680 ;
        RECT 243.520 72.870 249.030 73.680 ;
        RECT 249.040 72.870 254.550 73.680 ;
        RECT 255.020 72.770 258.675 73.680 ;
        RECT 258.700 72.870 264.210 73.680 ;
        RECT 265.150 72.810 265.580 73.595 ;
        RECT 265.600 72.870 271.110 73.680 ;
        RECT 271.120 72.870 276.630 73.680 ;
        RECT 276.640 72.870 278.470 73.680 ;
        RECT 278.480 72.770 281.230 73.680 ;
        RECT 281.240 72.870 284.910 73.680 ;
        RECT 285.840 73.000 290.655 73.680 ;
        RECT 290.910 72.810 291.340 73.595 ;
        RECT 291.360 72.870 293.190 73.680 ;
        RECT 293.660 72.900 295.030 73.680 ;
        RECT 295.040 73.000 304.650 73.680 ;
        RECT 299.550 72.780 300.480 73.000 ;
        RECT 303.310 72.770 304.650 73.000 ;
        RECT 304.700 72.870 308.370 73.680 ;
        RECT 308.380 72.870 309.750 73.680 ;
        RECT 309.760 72.870 311.130 73.680 ;
      LAYER nwell ;
        RECT 161.905 69.650 311.325 72.480 ;
      LAYER pwell ;
        RECT 162.100 68.450 163.470 69.260 ;
        RECT 163.480 68.450 165.310 69.260 ;
        RECT 169.830 69.130 170.760 69.350 ;
        RECT 173.590 69.130 174.930 69.360 ;
        RECT 165.320 68.450 174.930 69.130 ;
        RECT 174.990 68.535 175.420 69.320 ;
        RECT 176.360 69.130 177.290 69.360 ;
        RECT 176.360 68.450 180.260 69.130 ;
        RECT 180.500 68.450 186.010 69.260 ;
        RECT 186.020 68.450 187.850 69.260 ;
        RECT 188.320 68.450 189.690 69.230 ;
        RECT 189.700 69.130 190.630 69.360 ;
        RECT 193.840 69.130 195.185 69.360 ;
        RECT 199.340 69.130 200.270 69.360 ;
        RECT 189.700 68.450 193.600 69.130 ;
        RECT 193.840 68.450 195.670 69.130 ;
        RECT 196.370 68.450 200.270 69.130 ;
        RECT 200.750 68.535 201.180 69.320 ;
        RECT 201.200 68.450 203.030 69.260 ;
        RECT 203.040 68.450 206.240 69.360 ;
        RECT 206.260 68.450 209.460 69.360 ;
        RECT 209.480 68.450 212.220 69.130 ;
        RECT 212.240 68.450 214.070 69.130 ;
        RECT 214.080 68.450 219.590 69.260 ;
        RECT 219.600 68.450 225.110 69.260 ;
        RECT 225.120 68.450 226.490 69.260 ;
        RECT 226.510 68.535 226.940 69.320 ;
        RECT 226.960 68.450 230.615 69.360 ;
        RECT 230.640 68.450 232.010 69.260 ;
        RECT 162.240 68.240 162.410 68.450 ;
        RECT 163.620 68.240 163.790 68.450 ;
        RECT 165.460 68.260 165.630 68.450 ;
        RECT 170.060 68.240 170.230 68.430 ;
        RECT 170.520 68.240 170.690 68.430 ;
        RECT 171.900 68.240 172.070 68.430 ;
        RECT 175.590 68.295 175.750 68.405 ;
        RECT 176.775 68.260 176.945 68.450 ;
        RECT 180.640 68.260 180.810 68.450 ;
        RECT 181.560 68.240 181.730 68.430 ;
        RECT 185.240 68.240 185.410 68.430 ;
        RECT 186.160 68.260 186.330 68.450 ;
        RECT 186.620 68.240 186.790 68.430 ;
        RECT 187.995 68.290 188.115 68.400 ;
        RECT 188.460 68.240 188.630 68.430 ;
        RECT 189.380 68.260 189.550 68.450 ;
        RECT 190.115 68.260 190.285 68.450 ;
        RECT 195.360 68.260 195.530 68.450 ;
        RECT 195.815 68.290 195.935 68.400 ;
        RECT 198.395 68.240 198.565 68.430 ;
        RECT 199.685 68.260 199.855 68.450 ;
        RECT 200.415 68.290 200.535 68.400 ;
        RECT 201.340 68.260 201.510 68.450 ;
        RECT 202.260 68.240 202.430 68.430 ;
        RECT 204.095 68.290 204.215 68.400 ;
        RECT 205.945 68.260 206.115 68.450 ;
        RECT 208.695 68.240 208.865 68.430 ;
        RECT 209.165 68.260 209.335 68.450 ;
        RECT 209.620 68.260 209.790 68.450 ;
        RECT 212.380 68.260 212.550 68.450 ;
        RECT 213.295 68.240 213.465 68.430 ;
        RECT 214.220 68.240 214.390 68.450 ;
        RECT 216.980 68.240 217.150 68.430 ;
        RECT 219.740 68.260 219.910 68.450 ;
        RECT 220.670 68.285 220.830 68.395 ;
        RECT 221.580 68.260 221.750 68.430 ;
        RECT 225.260 68.240 225.430 68.450 ;
        RECT 227.105 68.260 227.275 68.450 ;
        RECT 162.100 67.430 163.470 68.240 ;
        RECT 163.480 67.430 168.990 68.240 ;
        RECT 169.000 67.460 170.370 68.240 ;
        RECT 170.380 67.460 171.750 68.240 ;
        RECT 171.760 67.560 181.370 68.240 ;
        RECT 176.270 67.340 177.200 67.560 ;
        RECT 180.030 67.330 181.370 67.560 ;
        RECT 181.420 67.430 185.090 68.240 ;
        RECT 185.100 67.460 186.470 68.240 ;
        RECT 186.480 67.460 187.850 68.240 ;
        RECT 187.870 67.370 188.300 68.155 ;
        RECT 188.320 67.560 197.930 68.240 ;
        RECT 192.830 67.340 193.760 67.560 ;
        RECT 196.590 67.330 197.930 67.560 ;
        RECT 197.980 67.560 201.880 68.240 ;
        RECT 197.980 67.330 198.910 67.560 ;
        RECT 202.120 67.430 203.950 68.240 ;
        RECT 205.380 68.010 209.010 68.240 ;
        RECT 209.980 68.010 213.610 68.240 ;
        RECT 204.420 67.330 209.010 68.010 ;
        RECT 209.020 67.330 213.610 68.010 ;
        RECT 213.630 67.370 214.060 68.155 ;
        RECT 214.080 67.560 216.820 68.240 ;
        RECT 216.840 67.430 220.510 68.240 ;
        RECT 221.780 67.560 225.110 68.240 ;
        RECT 222.285 67.330 225.110 67.560 ;
        RECT 225.120 67.330 228.330 68.240 ;
        RECT 228.340 68.210 229.295 68.240 ;
        RECT 230.325 68.210 230.495 68.430 ;
        RECT 230.780 68.240 230.950 68.450 ;
        RECT 232.020 68.410 232.910 69.360 ;
        RECT 236.600 69.130 237.530 69.360 ;
        RECT 233.860 68.450 237.530 69.130 ;
        RECT 237.540 68.450 243.050 69.260 ;
        RECT 245.135 69.130 246.270 69.360 ;
        RECT 243.060 68.450 246.270 69.130 ;
        RECT 246.280 68.450 251.790 69.260 ;
        RECT 252.270 68.535 252.700 69.320 ;
        RECT 252.720 68.450 256.375 69.360 ;
        RECT 258.460 69.270 259.410 69.360 ;
        RECT 257.480 68.450 259.410 69.270 ;
        RECT 259.620 68.450 265.130 69.260 ;
        RECT 265.140 68.450 270.650 69.260 ;
        RECT 270.660 68.450 272.490 69.260 ;
        RECT 272.500 69.130 273.430 69.360 ;
        RECT 272.500 68.450 276.400 69.130 ;
        RECT 276.640 68.450 278.010 69.260 ;
        RECT 278.030 68.535 278.460 69.320 ;
        RECT 278.480 68.450 281.230 69.360 ;
        RECT 281.240 68.450 282.610 69.230 ;
        RECT 282.620 69.130 283.550 69.360 ;
        RECT 286.760 69.130 287.690 69.360 ;
        RECT 282.620 68.450 286.520 69.130 ;
        RECT 286.760 68.450 290.660 69.130 ;
        RECT 290.900 68.450 293.650 69.260 ;
        RECT 298.630 69.130 299.560 69.350 ;
        RECT 302.390 69.130 303.730 69.360 ;
        RECT 294.120 68.450 303.730 69.130 ;
        RECT 303.790 68.535 304.220 69.320 ;
        RECT 304.725 69.130 306.070 69.360 ;
        RECT 304.240 68.450 306.070 69.130 ;
        RECT 306.080 68.450 307.910 69.260 ;
        RECT 308.380 68.450 309.750 69.230 ;
        RECT 309.760 68.450 311.130 69.260 ;
        RECT 232.620 68.260 232.790 68.410 ;
        RECT 233.090 68.295 233.250 68.405 ;
        RECT 234.000 68.260 234.170 68.450 ;
        RECT 236.300 68.240 236.470 68.430 ;
        RECT 237.680 68.260 237.850 68.450 ;
        RECT 243.200 68.260 243.370 68.450 ;
        RECT 246.420 68.260 246.590 68.450 ;
        RECT 248.720 68.240 248.890 68.430 ;
        RECT 249.180 68.240 249.350 68.430 ;
        RECT 251.935 68.290 252.055 68.400 ;
        RECT 252.865 68.260 253.035 68.450 ;
        RECT 257.480 68.430 257.630 68.450 ;
        RECT 254.700 68.240 254.870 68.430 ;
        RECT 256.550 68.295 256.710 68.405 ;
        RECT 257.460 68.260 257.630 68.430 ;
        RECT 257.915 68.290 258.035 68.400 ;
        RECT 259.760 68.260 259.930 68.450 ;
        RECT 261.595 68.240 261.765 68.430 ;
        RECT 264.820 68.240 264.990 68.430 ;
        RECT 265.280 68.260 265.450 68.450 ;
        RECT 265.740 68.240 265.910 68.430 ;
        RECT 268.495 68.290 268.615 68.400 ;
        RECT 268.960 68.240 269.130 68.430 ;
        RECT 270.340 68.240 270.510 68.430 ;
        RECT 270.800 68.260 270.970 68.450 ;
        RECT 272.915 68.260 273.085 68.450 ;
        RECT 276.780 68.260 276.950 68.450 ;
        RECT 279.995 68.290 280.115 68.400 ;
        RECT 280.460 68.240 280.630 68.430 ;
        RECT 280.920 68.260 281.090 68.450 ;
        RECT 282.300 68.260 282.470 68.450 ;
        RECT 283.035 68.260 283.205 68.450 ;
        RECT 287.175 68.260 287.345 68.450 ;
        RECT 289.660 68.240 289.830 68.430 ;
        RECT 291.040 68.260 291.210 68.450 ;
        RECT 291.500 68.240 291.670 68.430 ;
        RECT 293.800 68.400 293.970 68.430 ;
        RECT 293.335 68.290 293.455 68.400 ;
        RECT 293.795 68.290 293.970 68.400 ;
        RECT 293.800 68.240 293.970 68.290 ;
        RECT 294.260 68.260 294.430 68.450 ;
        RECT 295.180 68.240 295.350 68.430 ;
        RECT 304.380 68.260 304.550 68.450 ;
        RECT 306.220 68.260 306.390 68.450 ;
        RECT 307.140 68.240 307.310 68.430 ;
        RECT 307.600 68.240 307.770 68.430 ;
        RECT 309.440 68.400 309.610 68.450 ;
        RECT 308.055 68.290 308.175 68.400 ;
        RECT 309.435 68.290 309.610 68.400 ;
        RECT 309.440 68.260 309.610 68.290 ;
        RECT 310.820 68.240 310.990 68.450 ;
        RECT 228.340 67.530 230.620 68.210 ;
        RECT 228.340 67.330 229.295 67.530 ;
        RECT 230.640 67.430 236.150 68.240 ;
        RECT 236.160 67.330 239.370 68.240 ;
        RECT 239.390 67.370 239.820 68.155 ;
        RECT 239.925 67.560 249.030 68.240 ;
        RECT 249.040 67.430 254.550 68.240 ;
        RECT 254.560 67.330 257.770 68.240 ;
        RECT 258.255 67.330 261.910 68.240 ;
        RECT 261.920 67.330 265.130 68.240 ;
        RECT 265.150 67.370 265.580 68.155 ;
        RECT 265.600 67.430 268.350 68.240 ;
        RECT 268.820 67.460 270.190 68.240 ;
        RECT 270.200 67.560 279.810 68.240 ;
        RECT 280.320 67.560 289.510 68.240 ;
        RECT 274.710 67.340 275.640 67.560 ;
        RECT 278.470 67.330 279.810 67.560 ;
        RECT 284.830 67.340 285.760 67.560 ;
        RECT 288.590 67.330 289.510 67.560 ;
        RECT 289.520 67.430 290.890 68.240 ;
        RECT 290.910 67.370 291.340 68.155 ;
        RECT 291.360 67.430 293.190 68.240 ;
        RECT 293.660 67.460 295.030 68.240 ;
        RECT 295.040 67.560 304.650 68.240 ;
        RECT 304.710 67.560 307.450 68.240 ;
        RECT 299.550 67.340 300.480 67.560 ;
        RECT 303.310 67.330 304.650 67.560 ;
        RECT 307.460 67.430 309.290 68.240 ;
        RECT 309.760 67.430 311.130 68.240 ;
      LAYER nwell ;
        RECT 161.905 64.210 311.325 67.040 ;
      LAYER pwell ;
        RECT 162.100 63.010 163.470 63.820 ;
        RECT 163.480 63.010 165.310 63.820 ;
        RECT 169.830 63.690 170.760 63.910 ;
        RECT 173.590 63.690 174.930 63.920 ;
        RECT 165.320 63.010 174.930 63.690 ;
        RECT 174.990 63.095 175.420 63.880 ;
        RECT 175.440 63.690 176.370 63.920 ;
        RECT 175.440 63.010 179.340 63.690 ;
        RECT 179.580 63.010 185.090 63.820 ;
        RECT 190.530 63.690 191.460 63.910 ;
        RECT 194.290 63.690 195.630 63.920 ;
        RECT 186.020 63.010 195.630 63.690 ;
        RECT 195.680 63.010 199.350 63.820 ;
        RECT 199.360 63.010 200.730 63.820 ;
        RECT 200.750 63.095 201.180 63.880 ;
        RECT 201.200 63.010 203.030 63.820 ;
        RECT 203.500 63.720 204.430 63.920 ;
        RECT 205.760 63.720 206.710 63.920 ;
        RECT 203.500 63.240 206.710 63.720 ;
        RECT 203.645 63.040 206.710 63.240 ;
        RECT 162.240 62.800 162.410 63.010 ;
        RECT 163.620 62.820 163.790 63.010 ;
        RECT 165.000 62.800 165.170 62.990 ;
        RECT 165.460 62.800 165.630 63.010 ;
        RECT 168.215 62.850 168.335 62.960 ;
        RECT 169.600 62.800 169.770 62.990 ;
        RECT 170.060 62.800 170.230 62.990 ;
        RECT 171.895 62.850 172.015 62.960 ;
        RECT 172.635 62.800 172.805 62.990 ;
        RECT 175.855 62.820 176.025 63.010 ;
        RECT 176.775 62.800 176.945 62.990 ;
        RECT 179.720 62.820 179.890 63.010 ;
        RECT 180.640 62.800 180.810 62.990 ;
        RECT 185.250 62.855 185.410 62.965 ;
        RECT 186.160 62.800 186.330 63.010 ;
        RECT 188.460 62.800 188.630 62.990 ;
        RECT 193.060 62.800 193.230 62.990 ;
        RECT 193.520 62.800 193.690 62.990 ;
        RECT 195.820 62.820 195.990 63.010 ;
        RECT 199.040 62.800 199.210 62.990 ;
        RECT 199.500 62.820 199.670 63.010 ;
        RECT 201.340 62.820 201.510 63.010 ;
        RECT 203.175 62.850 203.295 62.960 ;
        RECT 203.645 62.820 203.815 63.040 ;
        RECT 205.775 63.010 206.710 63.040 ;
        RECT 206.890 63.240 211.240 63.920 ;
        RECT 211.320 63.720 212.250 63.920 ;
        RECT 213.580 63.720 214.530 63.920 ;
        RECT 211.320 63.240 214.530 63.720 ;
        RECT 206.890 63.010 210.660 63.240 ;
        RECT 211.465 63.040 214.530 63.240 ;
        RECT 206.890 62.990 207.030 63.010 ;
        RECT 205.485 62.800 205.655 62.990 ;
        RECT 205.940 62.800 206.110 62.990 ;
        RECT 206.860 62.820 207.030 62.990 ;
        RECT 162.100 61.990 163.470 62.800 ;
        RECT 163.480 62.120 165.310 62.800 ;
        RECT 163.480 61.890 164.825 62.120 ;
        RECT 165.320 61.990 168.070 62.800 ;
        RECT 168.540 62.020 169.910 62.800 ;
        RECT 169.920 61.990 171.750 62.800 ;
        RECT 172.220 62.120 176.120 62.800 ;
        RECT 176.360 62.120 180.260 62.800 ;
        RECT 172.220 61.890 173.150 62.120 ;
        RECT 176.360 61.890 177.290 62.120 ;
        RECT 180.500 61.990 186.010 62.800 ;
        RECT 186.020 61.990 187.850 62.800 ;
        RECT 187.870 61.930 188.300 62.715 ;
        RECT 188.320 61.990 191.990 62.800 ;
        RECT 192.000 62.020 193.370 62.800 ;
        RECT 193.380 61.990 198.890 62.800 ;
        RECT 198.900 61.990 202.570 62.800 ;
        RECT 202.580 61.890 205.780 62.800 ;
        RECT 205.800 61.990 207.630 62.800 ;
        RECT 207.780 62.770 207.950 62.990 ;
        RECT 210.540 62.800 210.710 62.990 ;
        RECT 211.465 62.820 211.635 63.040 ;
        RECT 213.595 63.010 214.530 63.040 ;
        RECT 214.540 63.010 220.050 63.820 ;
        RECT 221.000 63.010 224.650 63.920 ;
        RECT 224.660 63.010 226.010 63.920 ;
        RECT 226.510 63.095 226.940 63.880 ;
        RECT 226.960 63.010 232.470 63.820 ;
        RECT 232.480 63.010 237.990 63.820 ;
        RECT 238.000 63.010 239.830 63.820 ;
        RECT 242.580 63.690 243.510 63.920 ;
        RECT 239.840 63.010 243.510 63.690 ;
        RECT 243.520 63.010 249.030 63.820 ;
        RECT 251.295 63.720 252.250 63.920 ;
        RECT 249.970 63.040 252.250 63.720 ;
        RECT 252.270 63.095 252.700 63.880 ;
        RECT 213.295 62.850 213.415 62.960 ;
        RECT 214.220 62.820 214.390 62.990 ;
        RECT 214.680 62.820 214.850 63.010 ;
        RECT 216.980 62.820 217.150 62.990 ;
        RECT 219.740 62.820 219.910 62.990 ;
        RECT 220.210 62.855 220.370 62.965 ;
        RECT 214.250 62.800 214.390 62.820 ;
        RECT 217.010 62.800 217.150 62.820 ;
        RECT 219.770 62.800 219.910 62.820 ;
        RECT 222.500 62.800 222.670 62.990 ;
        RECT 224.335 62.820 224.505 63.010 ;
        RECT 225.725 62.820 225.895 63.010 ;
        RECT 226.175 62.850 226.295 62.960 ;
        RECT 227.100 62.820 227.270 63.010 ;
        RECT 228.030 62.845 228.190 62.955 ;
        RECT 228.940 62.820 229.110 62.990 ;
        RECT 232.620 62.820 232.790 63.010 ;
        RECT 228.945 62.800 229.110 62.820 ;
        RECT 234.455 62.800 234.625 62.990 ;
        RECT 234.925 62.800 235.095 62.990 ;
        RECT 238.140 62.800 238.310 63.010 ;
        RECT 239.980 62.800 240.150 63.010 ;
        RECT 243.660 62.820 243.830 63.010 ;
        RECT 245.500 62.800 245.670 62.990 ;
        RECT 249.190 62.855 249.350 62.965 ;
        RECT 250.095 62.820 250.265 63.040 ;
        RECT 251.295 63.010 252.250 63.040 ;
        RECT 252.735 63.010 256.390 63.920 ;
        RECT 257.320 63.010 259.610 63.920 ;
        RECT 259.620 63.010 265.130 63.820 ;
        RECT 265.140 63.010 266.970 63.820 ;
        RECT 266.980 63.010 268.350 63.790 ;
        RECT 268.400 63.690 269.740 63.920 ;
        RECT 272.570 63.690 273.500 63.910 ;
        RECT 268.400 63.010 278.010 63.690 ;
        RECT 278.030 63.095 278.460 63.880 ;
        RECT 278.480 63.010 283.990 63.820 ;
        RECT 284.000 63.010 289.510 63.820 ;
        RECT 293.640 63.690 294.570 63.920 ;
        RECT 298.700 63.690 299.630 63.920 ;
        RECT 290.670 63.010 294.570 63.690 ;
        RECT 295.730 63.010 299.630 63.690 ;
        RECT 299.640 63.010 303.310 63.820 ;
        RECT 303.790 63.095 304.220 63.880 ;
        RECT 304.240 63.010 309.750 63.820 ;
        RECT 309.760 63.010 311.130 63.820 ;
        RECT 251.020 62.800 251.190 62.990 ;
        RECT 254.700 62.800 254.870 62.990 ;
        RECT 255.160 62.800 255.330 62.990 ;
        RECT 256.075 62.820 256.245 63.010 ;
        RECT 256.550 62.855 256.710 62.965 ;
        RECT 257.460 62.820 257.630 63.010 ;
        RECT 258.380 62.800 258.550 62.990 ;
        RECT 258.840 62.800 259.010 62.990 ;
        RECT 259.760 62.820 259.930 63.010 ;
        RECT 264.370 62.845 264.530 62.955 ;
        RECT 265.280 62.820 265.450 63.010 ;
        RECT 265.740 62.800 265.910 62.990 ;
        RECT 267.120 62.820 267.290 63.010 ;
        RECT 270.800 62.800 270.970 62.990 ;
        RECT 271.260 62.800 271.430 62.990 ;
        RECT 272.915 62.800 273.085 62.990 ;
        RECT 276.780 62.800 276.950 62.990 ;
        RECT 277.700 62.820 277.870 63.010 ;
        RECT 278.620 62.820 278.790 63.010 ;
        RECT 280.920 62.800 281.090 62.990 ;
        RECT 281.390 62.845 281.550 62.955 ;
        RECT 282.575 62.800 282.745 62.990 ;
        RECT 284.140 62.820 284.310 63.010 ;
        RECT 289.670 62.855 289.830 62.965 ;
        RECT 289.845 62.800 290.015 62.990 ;
        RECT 290.575 62.850 290.695 62.960 ;
        RECT 291.500 62.800 291.670 62.990 ;
        RECT 292.880 62.800 293.050 62.990 ;
        RECT 293.985 62.820 294.155 63.010 ;
        RECT 294.260 62.800 294.430 62.990 ;
        RECT 294.730 62.855 294.890 62.965 ;
        RECT 299.045 62.820 299.215 63.010 ;
        RECT 299.780 62.820 299.950 63.010 ;
        RECT 303.455 62.850 303.575 62.960 ;
        RECT 303.920 62.800 304.090 62.990 ;
        RECT 304.380 62.820 304.550 63.010 ;
        RECT 309.435 62.850 309.555 62.960 ;
        RECT 310.820 62.800 310.990 63.010 ;
        RECT 208.995 62.770 210.390 62.800 ;
        RECT 207.655 62.090 210.390 62.770 ;
        RECT 210.400 62.120 213.140 62.800 ;
        RECT 208.980 61.890 210.390 62.090 ;
        RECT 213.630 61.930 214.060 62.715 ;
        RECT 214.250 61.980 216.820 62.800 ;
        RECT 217.010 61.980 219.580 62.800 ;
        RECT 219.770 61.980 222.340 62.800 ;
        RECT 222.360 61.990 227.870 62.800 ;
        RECT 228.945 62.120 230.780 62.800 ;
        RECT 215.230 61.890 216.820 61.980 ;
        RECT 217.990 61.890 219.580 61.980 ;
        RECT 220.750 61.890 222.340 61.980 ;
        RECT 229.850 61.890 230.780 62.120 ;
        RECT 231.295 61.890 234.770 62.800 ;
        RECT 234.780 61.890 237.700 62.800 ;
        RECT 238.000 61.990 239.370 62.800 ;
        RECT 239.390 61.930 239.820 62.715 ;
        RECT 239.840 61.990 245.350 62.800 ;
        RECT 245.360 61.990 250.870 62.800 ;
        RECT 250.880 61.990 252.250 62.800 ;
        RECT 252.260 61.890 255.010 62.800 ;
        RECT 255.020 61.990 256.850 62.800 ;
        RECT 256.860 61.890 258.675 62.800 ;
        RECT 258.700 61.990 264.210 62.800 ;
        RECT 265.150 61.930 265.580 62.715 ;
        RECT 265.600 61.990 267.430 62.800 ;
        RECT 267.535 62.120 271.000 62.800 ;
        RECT 267.535 61.890 268.455 62.120 ;
        RECT 271.120 61.990 272.490 62.800 ;
        RECT 272.500 62.120 276.400 62.800 ;
        RECT 272.500 61.890 273.430 62.120 ;
        RECT 276.640 61.990 278.470 62.800 ;
        RECT 278.480 61.890 281.230 62.800 ;
        RECT 282.160 62.120 286.060 62.800 ;
        RECT 286.530 62.120 290.430 62.800 ;
        RECT 282.160 61.890 283.090 62.120 ;
        RECT 289.500 61.890 290.430 62.120 ;
        RECT 290.910 61.930 291.340 62.715 ;
        RECT 291.360 61.990 292.730 62.800 ;
        RECT 292.740 62.020 294.110 62.800 ;
        RECT 294.120 62.120 303.730 62.800 ;
        RECT 298.630 61.900 299.560 62.120 ;
        RECT 302.390 61.890 303.730 62.120 ;
        RECT 303.780 61.990 309.290 62.800 ;
        RECT 309.760 61.990 311.130 62.800 ;
      LAYER nwell ;
        RECT 161.905 58.770 311.325 61.600 ;
      LAYER pwell ;
        RECT 162.100 57.570 163.470 58.380 ;
        RECT 163.480 57.570 165.310 58.380 ;
        RECT 169.830 58.250 170.760 58.470 ;
        RECT 173.590 58.250 174.930 58.480 ;
        RECT 165.320 57.570 174.930 58.250 ;
        RECT 174.990 57.655 175.420 58.440 ;
        RECT 175.900 58.250 176.830 58.480 ;
        RECT 180.040 58.250 180.970 58.480 ;
        RECT 175.900 57.570 179.800 58.250 ;
        RECT 180.040 57.570 183.940 58.250 ;
        RECT 184.180 57.570 187.850 58.380 ;
        RECT 192.370 58.250 193.300 58.470 ;
        RECT 196.020 58.250 198.230 58.480 ;
        RECT 187.860 57.570 198.230 58.250 ;
        RECT 198.440 57.570 199.810 58.350 ;
        RECT 200.750 57.655 201.180 58.440 ;
        RECT 201.200 57.570 203.030 58.380 ;
        RECT 203.040 58.250 203.970 58.480 ;
        RECT 217.310 58.390 218.900 58.480 ;
        RECT 203.040 57.570 206.940 58.250 ;
        RECT 207.180 57.570 209.920 58.250 ;
        RECT 209.940 57.570 215.450 58.380 ;
        RECT 215.460 57.570 217.290 58.380 ;
        RECT 217.310 57.570 219.880 58.390 ;
        RECT 220.060 57.570 223.730 58.380 ;
        RECT 224.510 58.250 225.440 58.480 ;
        RECT 224.510 57.570 226.345 58.250 ;
        RECT 226.510 57.655 226.940 58.440 ;
        RECT 227.155 57.570 230.630 58.480 ;
        RECT 230.640 57.570 234.675 58.480 ;
        RECT 234.780 57.570 237.700 58.480 ;
        RECT 239.970 58.250 240.900 58.480 ;
        RECT 239.065 57.570 240.900 58.250 ;
        RECT 241.220 57.570 244.140 58.480 ;
        RECT 162.240 57.360 162.410 57.570 ;
        RECT 163.620 57.360 163.790 57.570 ;
        RECT 165.460 57.380 165.630 57.570 ;
        RECT 167.300 57.360 167.470 57.550 ;
        RECT 167.760 57.360 167.930 57.550 ;
        RECT 175.575 57.410 175.695 57.520 ;
        RECT 176.315 57.380 176.485 57.570 ;
        RECT 177.420 57.360 177.590 57.550 ;
        RECT 180.455 57.380 180.625 57.570 ;
        RECT 184.320 57.380 184.490 57.570 ;
        RECT 188.000 57.380 188.170 57.570 ;
        RECT 188.460 57.360 188.630 57.550 ;
        RECT 191.220 57.360 191.390 57.550 ;
        RECT 199.500 57.380 199.670 57.570 ;
        RECT 199.970 57.415 200.130 57.525 ;
        RECT 200.880 57.360 201.050 57.550 ;
        RECT 201.340 57.380 201.510 57.570 ;
        RECT 202.995 57.360 203.165 57.550 ;
        RECT 203.455 57.380 203.625 57.570 ;
        RECT 207.320 57.380 207.490 57.570 ;
        RECT 210.080 57.360 210.250 57.570 ;
        RECT 210.545 57.360 210.715 57.550 ;
        RECT 215.600 57.380 215.770 57.570 ;
        RECT 219.740 57.550 219.880 57.570 ;
        RECT 216.975 57.360 217.145 57.550 ;
        RECT 217.440 57.360 217.610 57.550 ;
        RECT 219.740 57.380 219.910 57.550 ;
        RECT 220.200 57.380 220.370 57.570 ;
        RECT 226.180 57.550 226.345 57.570 ;
        RECT 223.880 57.520 224.050 57.550 ;
        RECT 222.970 57.405 223.130 57.515 ;
        RECT 223.875 57.410 224.050 57.520 ;
        RECT 223.880 57.360 224.050 57.410 ;
        RECT 225.720 57.360 225.890 57.550 ;
        RECT 226.180 57.380 226.350 57.550 ;
        RECT 230.315 57.380 230.485 57.570 ;
        RECT 230.785 57.380 230.955 57.570 ;
        RECT 234.925 57.550 235.095 57.570 ;
        RECT 239.065 57.550 239.230 57.570 ;
        RECT 234.455 57.360 234.625 57.550 ;
        RECT 234.920 57.380 235.095 57.550 ;
        RECT 238.150 57.415 238.310 57.525 ;
        RECT 238.610 57.405 238.770 57.515 ;
        RECT 239.060 57.380 239.230 57.550 ;
        RECT 234.920 57.360 235.090 57.380 ;
        RECT 239.985 57.360 240.155 57.550 ;
        RECT 241.365 57.380 241.535 57.570 ;
        RECT 243.660 57.360 243.830 57.550 ;
        RECT 244.590 57.415 244.750 57.525 ;
        RECT 162.100 56.550 163.470 57.360 ;
        RECT 163.480 56.550 166.230 57.360 ;
        RECT 166.240 56.580 167.610 57.360 ;
        RECT 167.620 56.680 177.230 57.360 ;
        RECT 177.280 56.680 187.650 57.360 ;
        RECT 172.130 56.460 173.060 56.680 ;
        RECT 175.890 56.450 177.230 56.680 ;
        RECT 181.790 56.460 182.720 56.680 ;
        RECT 185.440 56.450 187.650 56.680 ;
        RECT 187.870 56.490 188.300 57.275 ;
        RECT 188.320 56.550 191.070 57.360 ;
        RECT 191.080 56.680 200.690 57.360 ;
        RECT 195.590 56.460 196.520 56.680 ;
        RECT 199.350 56.450 200.690 56.680 ;
        RECT 200.740 56.550 202.570 57.360 ;
        RECT 202.580 56.680 206.480 57.360 ;
        RECT 206.720 56.680 210.390 57.360 ;
        RECT 202.580 56.450 203.510 56.680 ;
        RECT 206.720 56.450 207.650 56.680 ;
        RECT 210.400 56.450 213.610 57.360 ;
        RECT 213.630 56.490 214.060 57.275 ;
        RECT 214.080 56.450 217.290 57.360 ;
        RECT 217.300 56.550 222.810 57.360 ;
        RECT 223.740 56.680 225.570 57.360 ;
        RECT 224.225 56.450 225.570 56.680 ;
        RECT 225.580 56.450 229.710 57.360 ;
        RECT 229.900 56.450 234.770 57.360 ;
        RECT 234.780 56.550 238.450 57.360 ;
        RECT 239.390 56.490 239.820 57.275 ;
        RECT 239.840 56.450 243.315 57.360 ;
        RECT 243.520 56.550 244.890 57.360 ;
        RECT 245.035 57.330 245.205 57.550 ;
        RECT 245.380 57.530 246.270 58.480 ;
        RECT 248.250 58.250 249.180 58.480 ;
        RECT 249.985 58.250 251.330 58.480 ;
        RECT 247.345 57.570 249.180 58.250 ;
        RECT 249.500 57.570 251.330 58.250 ;
        RECT 252.270 57.655 252.700 58.440 ;
        RECT 252.720 57.570 254.090 58.380 ;
        RECT 254.295 57.570 257.770 58.480 ;
        RECT 258.830 58.250 259.760 58.480 ;
        RECT 257.925 57.570 259.760 58.250 ;
        RECT 260.830 57.570 263.750 58.480 ;
        RECT 263.760 57.570 266.970 58.480 ;
        RECT 266.980 57.570 268.350 58.380 ;
        RECT 268.455 58.250 269.375 58.480 ;
        RECT 268.455 57.570 271.920 58.250 ;
        RECT 272.040 57.570 277.550 58.380 ;
        RECT 278.030 57.655 278.460 58.440 ;
        RECT 278.940 57.570 280.310 58.350 ;
        RECT 284.830 58.250 285.760 58.470 ;
        RECT 288.590 58.250 289.510 58.480 ;
        RECT 280.320 57.570 289.510 58.250 ;
        RECT 289.520 57.570 290.890 58.350 ;
        RECT 290.900 57.570 294.570 58.380 ;
        RECT 294.580 58.250 295.510 58.480 ;
        RECT 294.580 57.570 298.480 58.250 ;
        RECT 298.720 57.570 300.090 58.350 ;
        RECT 300.100 57.570 303.770 58.380 ;
        RECT 303.790 57.655 304.220 58.440 ;
        RECT 304.240 57.570 309.750 58.380 ;
        RECT 309.760 57.570 311.130 58.380 ;
        RECT 247.345 57.550 247.510 57.570 ;
        RECT 245.500 57.380 245.670 57.530 ;
        RECT 246.430 57.415 246.590 57.525 ;
        RECT 247.340 57.520 247.510 57.550 ;
        RECT 247.335 57.410 247.510 57.520 ;
        RECT 247.340 57.380 247.510 57.410 ;
        RECT 247.795 57.360 247.965 57.550 ;
        RECT 249.640 57.380 249.810 57.570 ;
        RECT 251.490 57.415 251.650 57.525 ;
        RECT 252.860 57.380 253.030 57.570 ;
        RECT 254.700 57.360 254.870 57.550 ;
        RECT 246.235 57.330 247.190 57.360 ;
        RECT 244.910 56.650 247.190 57.330 ;
        RECT 246.235 56.450 247.190 56.650 ;
        RECT 247.670 56.450 250.870 57.360 ;
        RECT 250.880 56.450 255.010 57.360 ;
        RECT 255.160 57.330 255.330 57.550 ;
        RECT 257.455 57.380 257.625 57.570 ;
        RECT 257.925 57.550 258.090 57.570 ;
        RECT 257.920 57.380 258.090 57.550 ;
        RECT 258.380 57.360 258.550 57.550 ;
        RECT 260.215 57.410 260.335 57.520 ;
        RECT 261.135 57.410 261.255 57.520 ;
        RECT 261.595 57.380 261.765 57.550 ;
        RECT 263.435 57.380 263.605 57.570 ;
        RECT 266.660 57.380 266.830 57.570 ;
        RECT 267.120 57.380 267.290 57.570 ;
        RECT 261.630 57.360 261.765 57.380 ;
        RECT 269.420 57.360 269.590 57.550 ;
        RECT 269.880 57.360 270.050 57.550 ;
        RECT 271.720 57.520 271.890 57.570 ;
        RECT 271.715 57.410 271.890 57.520 ;
        RECT 271.720 57.380 271.890 57.410 ;
        RECT 272.180 57.380 272.350 57.570 ;
        RECT 277.695 57.410 277.815 57.520 ;
        RECT 278.615 57.410 278.735 57.520 ;
        RECT 279.080 57.380 279.250 57.570 ;
        RECT 280.460 57.380 280.630 57.570 ;
        RECT 280.920 57.360 281.090 57.550 ;
        RECT 290.580 57.360 290.750 57.570 ;
        RECT 291.040 57.380 291.210 57.570 ;
        RECT 291.500 57.360 291.670 57.550 ;
        RECT 293.340 57.360 293.510 57.550 ;
        RECT 294.720 57.360 294.890 57.550 ;
        RECT 294.995 57.380 295.165 57.570 ;
        RECT 297.480 57.360 297.650 57.550 ;
        RECT 299.780 57.380 299.950 57.570 ;
        RECT 300.240 57.380 300.410 57.570 ;
        RECT 304.380 57.380 304.550 57.570 ;
        RECT 307.140 57.360 307.310 57.550 ;
        RECT 309.440 57.360 309.610 57.550 ;
        RECT 310.820 57.360 310.990 57.570 ;
        RECT 257.285 57.330 258.230 57.360 ;
        RECT 255.160 57.130 258.230 57.330 ;
        RECT 255.020 56.650 258.230 57.130 ;
        RECT 255.020 56.450 255.950 56.650 ;
        RECT 257.285 56.450 258.230 56.650 ;
        RECT 258.240 56.550 260.990 57.360 ;
        RECT 261.630 56.450 265.130 57.360 ;
        RECT 265.150 56.490 265.580 57.275 ;
        RECT 265.670 56.450 269.730 57.360 ;
        RECT 269.740 56.550 271.570 57.360 ;
        RECT 272.040 56.680 281.230 57.360 ;
        RECT 281.280 56.680 290.890 57.360 ;
        RECT 272.040 56.450 272.960 56.680 ;
        RECT 275.790 56.460 276.720 56.680 ;
        RECT 281.280 56.450 282.620 56.680 ;
        RECT 285.450 56.460 286.380 56.680 ;
        RECT 290.910 56.490 291.340 57.275 ;
        RECT 291.360 56.550 293.190 57.360 ;
        RECT 293.200 56.580 294.570 57.360 ;
        RECT 294.580 56.550 297.330 57.360 ;
        RECT 297.340 56.680 306.950 57.360 ;
        RECT 301.850 56.460 302.780 56.680 ;
        RECT 305.610 56.450 306.950 56.680 ;
        RECT 307.000 56.550 308.370 57.360 ;
        RECT 308.380 56.580 309.750 57.360 ;
        RECT 309.760 56.550 311.130 57.360 ;
      LAYER nwell ;
        RECT 161.905 53.330 311.325 56.160 ;
      LAYER pwell ;
        RECT 162.100 52.130 163.470 52.940 ;
        RECT 163.480 52.130 165.310 52.940 ;
        RECT 169.830 52.810 170.760 53.030 ;
        RECT 173.590 52.810 174.930 53.040 ;
        RECT 165.320 52.130 174.930 52.810 ;
        RECT 174.990 52.215 175.420 53.000 ;
        RECT 175.440 52.130 176.810 52.910 ;
        RECT 176.820 52.130 180.490 52.940 ;
        RECT 180.500 52.130 181.870 52.910 ;
        RECT 181.880 52.130 187.390 52.940 ;
        RECT 187.400 52.130 190.150 52.940 ;
        RECT 190.395 52.130 195.210 52.810 ;
        RECT 195.220 52.130 200.730 52.940 ;
        RECT 200.750 52.215 201.180 53.000 ;
        RECT 201.235 52.360 206.710 53.040 ;
        RECT 162.240 51.920 162.410 52.130 ;
        RECT 163.620 51.920 163.790 52.130 ;
        RECT 165.460 51.940 165.630 52.130 ;
        RECT 169.140 51.920 169.310 52.110 ;
        RECT 174.660 51.920 174.830 52.110 ;
        RECT 176.500 51.940 176.670 52.130 ;
        RECT 176.960 51.940 177.130 52.130 ;
        RECT 180.180 51.920 180.350 52.110 ;
        RECT 181.560 51.940 181.730 52.130 ;
        RECT 182.020 51.940 182.190 52.130 ;
        RECT 185.700 51.920 185.870 52.110 ;
        RECT 187.540 52.080 187.710 52.130 ;
        RECT 187.535 51.970 187.710 52.080 ;
        RECT 187.540 51.940 187.710 51.970 ;
        RECT 188.460 51.920 188.630 52.110 ;
        RECT 194.440 51.920 194.610 52.110 ;
        RECT 194.900 51.920 195.070 52.130 ;
        RECT 195.360 51.940 195.530 52.130 ;
        RECT 198.575 51.970 198.695 52.080 ;
        RECT 199.040 51.920 199.210 52.110 ;
        RECT 200.420 51.920 200.590 52.110 ;
        RECT 201.340 51.940 201.510 52.360 ;
        RECT 202.620 52.130 206.710 52.360 ;
        RECT 206.720 52.130 209.470 52.940 ;
        RECT 209.965 52.810 211.305 53.040 ;
        RECT 216.160 52.810 217.750 53.040 ;
        RECT 209.480 52.130 214.070 52.810 ;
        RECT 214.080 52.130 217.750 52.810 ;
        RECT 218.050 52.130 220.970 53.040 ;
        RECT 221.240 52.130 225.110 53.040 ;
        RECT 225.120 52.130 226.490 52.940 ;
        RECT 226.510 52.215 226.940 53.000 ;
        RECT 226.960 52.130 230.170 53.040 ;
        RECT 230.735 52.810 231.655 53.040 ;
        RECT 230.735 52.130 234.200 52.810 ;
        RECT 234.490 52.130 237.990 53.040 ;
        RECT 238.000 52.130 242.130 53.040 ;
        RECT 242.140 52.130 244.890 52.940 ;
        RECT 245.070 52.130 248.570 53.040 ;
        RECT 248.580 52.840 249.530 53.040 ;
        RECT 250.860 52.840 251.790 53.040 ;
        RECT 248.580 52.360 251.790 52.840 ;
        RECT 248.580 52.160 251.645 52.360 ;
        RECT 252.270 52.215 252.700 53.000 ;
        RECT 248.580 52.130 249.515 52.160 ;
        RECT 205.755 51.920 205.925 52.110 ;
        RECT 206.860 51.940 207.030 52.130 ;
        RECT 209.625 52.110 209.795 52.130 ;
        RECT 214.225 52.110 214.395 52.130 ;
        RECT 209.620 51.940 209.795 52.110 ;
        RECT 212.850 51.965 213.010 52.075 ;
        RECT 214.220 51.940 214.395 52.110 ;
        RECT 220.655 51.940 220.825 52.130 ;
        RECT 224.795 52.110 224.965 52.130 ;
        RECT 209.620 51.920 209.790 51.940 ;
        RECT 214.220 51.920 214.390 51.940 ;
        RECT 222.500 51.920 222.670 52.110 ;
        RECT 222.960 51.920 223.130 52.110 ;
        RECT 224.795 51.940 224.970 52.110 ;
        RECT 225.260 51.940 225.430 52.130 ;
        RECT 227.100 51.940 227.270 52.130 ;
        RECT 230.315 51.970 230.435 52.080 ;
        RECT 224.800 51.920 224.970 51.940 ;
        RECT 234.000 51.920 234.170 52.130 ;
        RECT 234.490 52.110 234.625 52.130 ;
        RECT 234.455 51.940 234.625 52.110 ;
        RECT 235.835 51.970 235.955 52.080 ;
        RECT 238.140 51.940 238.310 52.130 ;
        RECT 239.060 51.920 239.230 52.110 ;
        RECT 242.280 51.940 242.450 52.130 ;
        RECT 245.070 52.110 245.205 52.130 ;
        RECT 243.200 51.920 243.370 52.110 ;
        RECT 243.660 51.920 243.830 52.110 ;
        RECT 245.035 51.940 245.205 52.110 ;
        RECT 248.720 51.920 248.890 52.110 ;
        RECT 249.180 51.920 249.350 52.110 ;
        RECT 251.475 51.940 251.645 52.160 ;
        RECT 252.740 52.130 254.090 53.040 ;
        RECT 254.100 52.130 259.610 52.940 ;
        RECT 260.670 52.810 261.600 53.040 ;
        RECT 266.430 52.810 267.360 53.030 ;
        RECT 270.190 52.810 271.110 53.040 ;
        RECT 259.765 52.130 261.600 52.810 ;
        RECT 261.920 52.130 271.110 52.810 ;
        RECT 271.215 52.810 272.135 53.040 ;
        RECT 271.215 52.130 274.680 52.810 ;
        RECT 274.800 52.130 277.550 52.940 ;
        RECT 278.030 52.215 278.460 53.000 ;
        RECT 280.520 52.950 281.470 53.040 ;
        RECT 291.560 52.950 292.510 53.040 ;
        RECT 278.480 52.130 280.310 52.940 ;
        RECT 280.520 52.130 282.450 52.950 ;
        RECT 282.620 52.130 284.450 52.940 ;
        RECT 284.460 52.130 289.275 52.810 ;
        RECT 289.520 52.130 291.350 52.940 ;
        RECT 291.560 52.130 293.490 52.950 ;
        RECT 299.090 52.810 300.020 53.030 ;
        RECT 302.850 52.810 303.770 53.040 ;
        RECT 294.580 52.130 303.770 52.810 ;
        RECT 303.790 52.215 304.220 53.000 ;
        RECT 304.240 52.130 306.070 52.940 ;
        RECT 306.175 52.810 307.095 53.040 ;
        RECT 306.175 52.130 309.640 52.810 ;
        RECT 309.760 52.130 311.130 52.940 ;
        RECT 251.935 51.970 252.055 52.080 ;
        RECT 252.855 51.940 253.025 52.130 ;
        RECT 254.240 51.940 254.410 52.130 ;
        RECT 259.765 52.110 259.930 52.130 ;
        RECT 259.300 51.920 259.470 52.110 ;
        RECT 259.760 51.940 259.935 52.110 ;
        RECT 262.060 51.940 262.230 52.130 ;
        RECT 259.765 51.920 259.935 51.940 ;
        RECT 263.440 51.920 263.610 52.110 ;
        RECT 265.740 51.920 265.910 52.110 ;
        RECT 274.480 51.940 274.650 52.130 ;
        RECT 274.940 51.940 275.110 52.130 ;
        RECT 274.960 51.920 275.110 51.940 ;
        RECT 277.240 51.920 277.410 52.110 ;
        RECT 277.695 51.970 277.815 52.080 ;
        RECT 278.620 51.940 278.790 52.130 ;
        RECT 282.300 52.110 282.450 52.130 ;
        RECT 280.925 51.920 281.095 52.110 ;
        RECT 282.300 51.940 282.470 52.110 ;
        RECT 282.760 51.940 282.930 52.130 ;
        RECT 284.600 51.920 284.770 52.130 ;
        RECT 289.660 51.920 289.830 52.130 ;
        RECT 293.340 52.110 293.490 52.130 ;
        RECT 291.500 51.920 291.670 52.110 ;
        RECT 293.340 51.940 293.510 52.110 ;
        RECT 293.810 51.975 293.970 52.085 ;
        RECT 294.720 51.940 294.890 52.130 ;
        RECT 295.175 51.970 295.295 52.080 ;
        RECT 295.915 51.920 296.085 52.110 ;
        RECT 299.780 51.920 299.950 52.110 ;
        RECT 304.380 51.940 304.550 52.130 ;
        RECT 309.440 52.080 309.610 52.130 ;
        RECT 309.435 51.970 309.610 52.080 ;
        RECT 309.440 51.940 309.610 51.970 ;
        RECT 310.820 51.920 310.990 52.130 ;
        RECT 162.100 51.110 163.470 51.920 ;
        RECT 163.480 51.110 168.990 51.920 ;
        RECT 169.000 51.110 174.510 51.920 ;
        RECT 174.520 51.110 180.030 51.920 ;
        RECT 180.040 51.110 185.550 51.920 ;
        RECT 185.560 51.110 187.390 51.920 ;
        RECT 187.870 51.050 188.300 51.835 ;
        RECT 188.320 51.110 189.690 51.920 ;
        RECT 189.935 51.240 194.750 51.920 ;
        RECT 194.760 51.110 198.430 51.920 ;
        RECT 198.900 51.140 200.270 51.920 ;
        RECT 200.420 51.690 205.325 51.920 ;
        RECT 200.280 51.010 205.325 51.690 ;
        RECT 205.340 51.240 209.240 51.920 ;
        RECT 209.480 51.240 212.690 51.920 ;
        RECT 205.340 51.010 206.270 51.240 ;
        RECT 211.555 51.010 212.690 51.240 ;
        RECT 213.630 51.050 214.060 51.835 ;
        RECT 214.080 51.240 217.750 51.920 ;
        RECT 217.995 51.240 222.810 51.920 ;
        RECT 216.820 51.010 217.750 51.240 ;
        RECT 222.820 51.110 224.650 51.920 ;
        RECT 224.660 51.240 233.850 51.920 ;
        RECT 229.170 51.020 230.100 51.240 ;
        RECT 232.930 51.010 233.850 51.240 ;
        RECT 233.860 51.110 235.690 51.920 ;
        RECT 236.160 51.010 239.370 51.920 ;
        RECT 239.390 51.050 239.820 51.835 ;
        RECT 239.935 51.240 243.400 51.920 ;
        RECT 239.935 51.010 240.855 51.240 ;
        RECT 243.520 51.110 245.350 51.920 ;
        RECT 245.455 51.240 248.920 51.920 ;
        RECT 245.455 51.010 246.375 51.240 ;
        RECT 249.040 51.110 254.550 51.920 ;
        RECT 254.795 51.240 259.610 51.920 ;
        RECT 259.620 51.240 263.290 51.920 ;
        RECT 259.620 51.010 260.545 51.240 ;
        RECT 263.300 51.110 265.130 51.920 ;
        RECT 265.150 51.050 265.580 51.835 ;
        RECT 265.600 51.240 274.790 51.920 ;
        RECT 270.110 51.020 271.040 51.240 ;
        RECT 273.870 51.010 274.790 51.240 ;
        RECT 274.960 51.100 276.890 51.920 ;
        RECT 277.210 51.240 280.675 51.920 ;
        RECT 275.940 51.010 276.890 51.100 ;
        RECT 279.755 51.010 280.675 51.240 ;
        RECT 280.780 51.010 284.435 51.920 ;
        RECT 284.460 51.240 289.275 51.920 ;
        RECT 289.520 51.110 290.890 51.920 ;
        RECT 290.910 51.050 291.340 51.835 ;
        RECT 291.470 51.240 294.935 51.920 ;
        RECT 294.015 51.010 294.935 51.240 ;
        RECT 295.500 51.240 299.400 51.920 ;
        RECT 299.640 51.240 308.920 51.920 ;
        RECT 295.500 51.010 296.430 51.240 ;
        RECT 301.000 51.020 301.920 51.240 ;
        RECT 306.585 51.120 308.920 51.240 ;
        RECT 308.000 51.010 308.920 51.120 ;
        RECT 309.760 51.110 311.130 51.920 ;
      LAYER nwell ;
        RECT 161.905 47.890 311.325 50.720 ;
      LAYER pwell ;
        RECT 162.100 46.690 163.470 47.500 ;
        RECT 163.480 46.690 168.990 47.500 ;
        RECT 169.000 46.690 174.510 47.500 ;
        RECT 174.990 46.775 175.420 47.560 ;
        RECT 175.440 46.690 176.810 47.500 ;
        RECT 176.820 46.690 178.190 47.470 ;
        RECT 178.200 46.690 179.570 47.500 ;
        RECT 184.090 47.370 185.020 47.590 ;
        RECT 187.740 47.370 189.950 47.600 ;
        RECT 179.580 46.690 189.950 47.370 ;
        RECT 190.160 46.690 191.530 47.470 ;
        RECT 196.050 47.370 196.980 47.590 ;
        RECT 199.810 47.370 200.730 47.600 ;
        RECT 191.540 46.690 200.730 47.370 ;
        RECT 200.750 46.775 201.180 47.560 ;
        RECT 201.210 46.690 203.950 47.370 ;
        RECT 204.440 46.690 205.790 47.600 ;
        RECT 205.800 46.690 208.550 47.500 ;
        RECT 213.620 47.400 214.550 47.600 ;
        RECT 215.880 47.400 216.830 47.600 ;
        RECT 218.900 47.510 219.850 47.600 ;
        RECT 208.795 46.690 213.610 47.370 ;
        RECT 213.620 46.920 216.830 47.400 ;
        RECT 213.765 46.720 216.830 46.920 ;
        RECT 162.240 46.480 162.410 46.690 ;
        RECT 163.620 46.480 163.790 46.690 ;
        RECT 169.140 46.480 169.310 46.690 ;
        RECT 172.830 46.525 172.990 46.635 ;
        RECT 174.655 46.530 174.775 46.640 ;
        RECT 175.580 46.500 175.750 46.690 ;
        RECT 176.960 46.480 177.130 46.690 ;
        RECT 177.420 46.480 177.590 46.670 ;
        RECT 178.340 46.500 178.510 46.690 ;
        RECT 179.720 46.500 179.890 46.690 ;
        RECT 188.735 46.480 188.905 46.670 ;
        RECT 190.300 46.500 190.470 46.690 ;
        RECT 191.680 46.500 191.850 46.690 ;
        RECT 192.610 46.525 192.770 46.635 ;
        RECT 193.795 46.480 193.965 46.670 ;
        RECT 197.660 46.480 197.830 46.670 ;
        RECT 199.495 46.530 199.615 46.640 ;
        RECT 199.960 46.480 200.130 46.670 ;
        RECT 203.640 46.500 203.810 46.690 ;
        RECT 204.095 46.530 204.215 46.640 ;
        RECT 205.475 46.500 205.645 46.690 ;
        RECT 205.940 46.500 206.110 46.690 ;
        RECT 210.540 46.480 210.710 46.670 ;
        RECT 213.300 46.640 213.470 46.690 ;
        RECT 213.295 46.530 213.470 46.640 ;
        RECT 213.300 46.500 213.470 46.530 ;
        RECT 213.765 46.500 213.935 46.720 ;
        RECT 215.895 46.690 216.830 46.720 ;
        RECT 217.920 46.690 219.850 47.510 ;
        RECT 220.060 46.690 221.890 47.500 ;
        RECT 222.845 47.370 224.190 47.600 ;
        RECT 222.360 46.690 224.190 47.370 ;
        RECT 224.660 46.690 226.030 47.470 ;
        RECT 226.510 46.775 226.940 47.560 ;
        RECT 227.445 47.370 228.790 47.600 ;
        RECT 234.230 47.370 235.160 47.590 ;
        RECT 237.990 47.370 238.910 47.600 ;
        RECT 243.430 47.370 244.360 47.590 ;
        RECT 247.190 47.370 248.110 47.600 ;
        RECT 226.960 46.690 228.790 47.370 ;
        RECT 229.720 46.690 238.910 47.370 ;
        RECT 238.920 46.690 248.110 47.370 ;
        RECT 248.120 46.690 251.790 47.500 ;
        RECT 252.270 46.775 252.700 47.560 ;
        RECT 252.720 46.690 255.470 47.500 ;
        RECT 259.990 47.370 260.920 47.590 ;
        RECT 263.750 47.370 264.670 47.600 ;
        RECT 267.335 47.370 268.255 47.600 ;
        RECT 255.480 46.690 264.670 47.370 ;
        RECT 264.790 46.690 268.255 47.370 ;
        RECT 268.375 46.690 272.030 47.600 ;
        RECT 272.055 46.690 275.710 47.600 ;
        RECT 275.920 47.510 276.870 47.600 ;
        RECT 275.920 46.690 277.850 47.510 ;
        RECT 278.030 46.775 278.460 47.560 ;
        RECT 278.575 47.370 279.495 47.600 ;
        RECT 282.360 47.510 283.310 47.600 ;
        RECT 278.575 46.690 282.040 47.370 ;
        RECT 282.360 46.690 284.290 47.510 ;
        RECT 285.380 47.370 286.300 47.600 ;
        RECT 289.130 47.370 290.060 47.590 ;
        RECT 299.090 47.370 300.020 47.590 ;
        RECT 302.850 47.370 303.770 47.600 ;
        RECT 285.380 46.690 294.570 47.370 ;
        RECT 294.580 46.690 303.770 47.370 ;
        RECT 303.790 46.775 304.220 47.560 ;
        RECT 304.335 47.370 305.255 47.600 ;
        RECT 304.335 46.690 307.800 47.370 ;
        RECT 307.920 46.690 309.750 47.500 ;
        RECT 309.760 46.690 311.130 47.500 ;
        RECT 217.920 46.670 218.070 46.690 ;
        RECT 214.230 46.525 214.390 46.635 ;
        RECT 215.140 46.480 215.310 46.670 ;
        RECT 216.980 46.480 217.150 46.670 ;
        RECT 217.900 46.500 218.070 46.670 ;
        RECT 218.360 46.480 218.530 46.670 ;
        RECT 219.740 46.480 219.910 46.670 ;
        RECT 220.200 46.500 220.370 46.690 ;
        RECT 222.035 46.530 222.155 46.640 ;
        RECT 222.500 46.500 222.670 46.690 ;
        RECT 224.335 46.530 224.455 46.640 ;
        RECT 225.720 46.500 225.890 46.690 ;
        RECT 226.175 46.530 226.295 46.640 ;
        RECT 227.100 46.500 227.270 46.690 ;
        RECT 228.950 46.535 229.110 46.645 ;
        RECT 229.860 46.500 230.030 46.690 ;
        RECT 230.320 46.480 230.490 46.670 ;
        RECT 233.080 46.480 233.250 46.670 ;
        RECT 238.610 46.525 238.770 46.635 ;
        RECT 239.060 46.500 239.230 46.690 ;
        RECT 239.980 46.480 240.150 46.670 ;
        RECT 243.660 46.480 243.830 46.670 ;
        RECT 248.260 46.500 248.430 46.690 ;
        RECT 252.860 46.640 253.030 46.690 ;
        RECT 251.935 46.530 252.055 46.640 ;
        RECT 252.855 46.530 253.030 46.640 ;
        RECT 252.860 46.500 253.030 46.530 ;
        RECT 255.620 46.500 255.790 46.690 ;
        RECT 256.540 46.480 256.710 46.670 ;
        RECT 258.840 46.500 259.010 46.670 ;
        RECT 259.310 46.525 259.470 46.635 ;
        RECT 258.840 46.480 258.990 46.500 ;
        RECT 264.820 46.480 264.990 46.690 ;
        RECT 268.960 46.480 269.130 46.670 ;
        RECT 269.420 46.500 269.590 46.670 ;
        RECT 271.715 46.635 271.885 46.690 ;
        RECT 271.715 46.525 271.890 46.635 ;
        RECT 271.715 46.500 271.885 46.525 ;
        RECT 269.440 46.480 269.590 46.500 ;
        RECT 272.640 46.480 272.810 46.670 ;
        RECT 275.395 46.500 275.565 46.690 ;
        RECT 277.700 46.670 277.850 46.690 ;
        RECT 277.700 46.500 277.870 46.670 ;
        RECT 281.840 46.500 282.010 46.690 ;
        RECT 284.140 46.670 284.290 46.690 ;
        RECT 284.140 46.500 284.310 46.670 ;
        RECT 284.610 46.535 284.770 46.645 ;
        RECT 290.580 46.480 290.750 46.670 ;
        RECT 291.505 46.480 291.675 46.670 ;
        RECT 294.260 46.500 294.430 46.690 ;
        RECT 294.720 46.500 294.890 46.690 ;
        RECT 295.175 46.530 295.295 46.640 ;
        RECT 295.640 46.480 295.810 46.670 ;
        RECT 299.315 46.530 299.435 46.640 ;
        RECT 307.600 46.500 307.770 46.690 ;
        RECT 308.060 46.500 308.230 46.690 ;
        RECT 308.980 46.480 309.150 46.670 ;
        RECT 309.435 46.530 309.555 46.640 ;
        RECT 310.820 46.480 310.990 46.690 ;
        RECT 162.100 45.670 163.470 46.480 ;
        RECT 163.480 45.670 168.990 46.480 ;
        RECT 169.000 45.670 172.670 46.480 ;
        RECT 173.695 45.800 177.160 46.480 ;
        RECT 177.280 45.800 187.650 46.480 ;
        RECT 173.695 45.570 174.615 45.800 ;
        RECT 181.790 45.580 182.720 45.800 ;
        RECT 185.440 45.570 187.650 45.800 ;
        RECT 187.870 45.610 188.300 46.395 ;
        RECT 188.320 45.800 192.220 46.480 ;
        RECT 193.380 45.800 197.280 46.480 ;
        RECT 188.320 45.570 189.250 45.800 ;
        RECT 193.380 45.570 194.310 45.800 ;
        RECT 197.520 45.670 199.350 46.480 ;
        RECT 199.820 45.800 210.190 46.480 ;
        RECT 204.330 45.580 205.260 45.800 ;
        RECT 207.980 45.570 210.190 45.800 ;
        RECT 210.400 45.670 213.150 46.480 ;
        RECT 213.630 45.610 214.060 46.395 ;
        RECT 215.000 45.800 216.830 46.480 ;
        RECT 216.850 45.570 218.200 46.480 ;
        RECT 218.220 45.670 219.590 46.480 ;
        RECT 219.600 45.800 229.970 46.480 ;
        RECT 230.180 45.800 232.920 46.480 ;
        RECT 224.110 45.580 225.040 45.800 ;
        RECT 227.760 45.570 229.970 45.800 ;
        RECT 232.940 45.670 238.450 46.480 ;
        RECT 239.390 45.610 239.820 46.395 ;
        RECT 239.840 45.670 243.510 46.480 ;
        RECT 243.520 45.800 252.710 46.480 ;
        RECT 248.030 45.580 248.960 45.800 ;
        RECT 251.790 45.570 252.710 45.800 ;
        RECT 253.275 45.800 256.740 46.480 ;
        RECT 253.275 45.570 254.195 45.800 ;
        RECT 257.060 45.660 258.990 46.480 ;
        RECT 260.315 45.800 265.130 46.480 ;
        RECT 257.060 45.570 258.010 45.660 ;
        RECT 265.150 45.610 265.580 46.395 ;
        RECT 265.695 45.800 269.160 46.480 ;
        RECT 265.695 45.570 266.615 45.800 ;
        RECT 269.440 45.660 271.370 46.480 ;
        RECT 272.500 45.800 281.690 46.480 ;
        RECT 270.420 45.570 271.370 45.660 ;
        RECT 277.010 45.580 277.940 45.800 ;
        RECT 280.770 45.570 281.690 45.800 ;
        RECT 281.700 45.800 290.890 46.480 ;
        RECT 281.700 45.570 282.620 45.800 ;
        RECT 285.450 45.580 286.380 45.800 ;
        RECT 290.910 45.610 291.340 46.395 ;
        RECT 291.360 45.570 295.015 46.480 ;
        RECT 295.610 45.800 299.075 46.480 ;
        RECT 298.155 45.570 299.075 45.800 ;
        RECT 300.010 45.800 309.290 46.480 ;
        RECT 300.010 45.680 302.345 45.800 ;
        RECT 300.010 45.570 300.930 45.680 ;
        RECT 307.010 45.580 307.930 45.800 ;
        RECT 309.760 45.670 311.130 46.480 ;
      LAYER nwell ;
        RECT 161.905 42.450 311.325 45.280 ;
      LAYER pwell ;
        RECT 162.100 41.250 163.470 42.060 ;
        RECT 163.480 41.250 168.990 42.060 ;
        RECT 169.920 41.250 171.290 42.030 ;
        RECT 173.955 41.930 174.875 42.160 ;
        RECT 171.410 41.250 174.875 41.930 ;
        RECT 174.990 41.335 175.420 42.120 ;
        RECT 175.440 41.930 176.370 42.160 ;
        RECT 175.440 41.250 179.340 41.930 ;
        RECT 180.040 41.250 181.410 42.030 ;
        RECT 181.880 41.930 182.810 42.160 ;
        RECT 188.675 41.930 189.595 42.160 ;
        RECT 194.670 41.930 195.600 42.150 ;
        RECT 198.320 41.930 200.530 42.160 ;
        RECT 181.880 41.250 185.780 41.930 ;
        RECT 186.130 41.250 189.595 41.930 ;
        RECT 190.160 41.250 200.530 41.930 ;
        RECT 200.750 41.335 201.180 42.120 ;
        RECT 205.710 41.930 206.640 42.150 ;
        RECT 209.360 41.930 211.570 42.160 ;
        RECT 213.600 41.930 214.530 42.160 ;
        RECT 221.810 41.930 222.740 42.150 ;
        RECT 225.570 41.930 226.490 42.160 ;
        RECT 201.200 41.250 211.570 41.930 ;
        RECT 211.780 41.250 214.530 41.930 ;
        RECT 214.540 41.250 217.280 41.930 ;
        RECT 217.300 41.250 226.490 41.930 ;
        RECT 226.510 41.335 226.940 42.120 ;
        RECT 227.160 41.930 229.370 42.160 ;
        RECT 232.090 41.930 233.020 42.150 ;
        RECT 237.635 41.930 238.555 42.160 ;
        RECT 227.160 41.250 237.530 41.930 ;
        RECT 237.635 41.250 241.100 41.930 ;
        RECT 241.220 41.250 243.050 42.060 ;
        RECT 243.615 41.930 244.535 42.160 ;
        RECT 243.615 41.250 247.080 41.930 ;
        RECT 247.200 41.250 250.870 42.060 ;
        RECT 250.880 41.250 252.250 42.060 ;
        RECT 252.270 41.335 252.700 42.120 ;
        RECT 252.720 41.250 255.930 42.160 ;
        RECT 256.400 41.250 260.055 42.160 ;
        RECT 265.510 41.930 266.440 42.150 ;
        RECT 269.270 41.930 270.190 42.160 ;
        RECT 261.000 41.250 270.190 41.930 ;
        RECT 270.295 41.930 271.215 42.160 ;
        RECT 276.535 41.930 277.455 42.160 ;
        RECT 270.295 41.250 273.760 41.930 ;
        RECT 273.990 41.250 277.455 41.930 ;
        RECT 278.030 41.335 278.460 42.120 ;
        RECT 278.480 41.250 282.135 42.160 ;
        RECT 282.255 41.930 283.175 42.160 ;
        RECT 288.495 41.930 289.415 42.160 ;
        RECT 282.255 41.250 285.720 41.930 ;
        RECT 285.950 41.250 289.415 41.930 ;
        RECT 290.450 41.250 293.190 41.930 ;
        RECT 293.200 41.250 295.030 42.060 ;
        RECT 297.895 41.930 298.815 42.160 ;
        RECT 295.050 41.250 297.790 41.930 ;
        RECT 297.895 41.250 301.360 41.930 ;
        RECT 301.940 41.250 303.770 41.930 ;
        RECT 303.790 41.335 304.220 42.120 ;
        RECT 305.160 41.250 307.900 41.930 ;
        RECT 307.920 41.250 309.750 42.060 ;
        RECT 309.760 41.250 311.130 42.060 ;
        RECT 162.240 41.040 162.410 41.250 ;
        RECT 163.620 41.060 163.790 41.250 ;
        RECT 164.540 41.040 164.710 41.230 ;
        RECT 169.150 41.095 169.310 41.205 ;
        RECT 170.980 41.060 171.150 41.250 ;
        RECT 171.440 41.060 171.610 41.250 ;
        RECT 175.855 41.060 176.025 41.250 ;
        RECT 179.715 41.090 179.835 41.200 ;
        RECT 181.100 41.060 181.270 41.250 ;
        RECT 181.555 41.090 181.675 41.200 ;
        RECT 182.295 41.060 182.465 41.250 ;
        RECT 182.480 41.040 182.650 41.230 ;
        RECT 186.160 41.040 186.330 41.250 ;
        RECT 187.540 41.040 187.710 41.230 ;
        RECT 188.460 41.040 188.630 41.230 ;
        RECT 189.840 41.200 190.010 41.230 ;
        RECT 189.835 41.090 190.010 41.200 ;
        RECT 189.840 41.040 190.010 41.090 ;
        RECT 190.300 41.060 190.470 41.250 ;
        RECT 192.140 41.040 192.310 41.230 ;
        RECT 192.600 41.040 192.770 41.230 ;
        RECT 194.255 41.040 194.425 41.230 ;
        RECT 201.340 41.040 201.510 41.250 ;
        RECT 201.800 41.040 201.970 41.230 ;
        RECT 203.180 41.040 203.350 41.230 ;
        RECT 204.560 41.040 204.730 41.230 ;
        RECT 211.920 41.060 212.090 41.250 ;
        RECT 214.220 41.040 214.390 41.230 ;
        RECT 214.680 41.060 214.850 41.250 ;
        RECT 217.440 41.060 217.610 41.250 ;
        RECT 220.660 41.040 220.830 41.230 ;
        RECT 221.120 41.040 221.290 41.230 ;
        RECT 222.775 41.040 222.945 41.230 ;
        RECT 226.635 41.090 226.755 41.200 ;
        RECT 227.100 41.040 227.270 41.230 ;
        RECT 228.755 41.040 228.925 41.230 ;
        RECT 232.895 41.040 233.065 41.230 ;
        RECT 236.760 41.040 236.930 41.230 ;
        RECT 237.220 41.060 237.390 41.250 ;
        RECT 239.975 41.090 240.095 41.200 ;
        RECT 240.440 41.040 240.610 41.230 ;
        RECT 240.900 41.060 241.070 41.250 ;
        RECT 241.360 41.060 241.530 41.250 ;
        RECT 243.195 41.090 243.315 41.200 ;
        RECT 244.115 41.090 244.235 41.200 ;
        RECT 244.855 41.040 245.025 41.230 ;
        RECT 246.880 41.060 247.050 41.250 ;
        RECT 247.340 41.060 247.510 41.250 ;
        RECT 248.720 41.040 248.890 41.230 ;
        RECT 251.020 41.060 251.190 41.250 ;
        RECT 255.620 41.060 255.790 41.250 ;
        RECT 256.075 41.090 256.195 41.200 ;
        RECT 256.545 41.060 256.715 41.250 ;
        RECT 260.230 41.095 260.390 41.205 ;
        RECT 261.140 41.040 261.310 41.250 ;
        RECT 264.820 41.040 264.990 41.230 ;
        RECT 265.740 41.040 265.910 41.230 ;
        RECT 267.580 41.040 267.750 41.230 ;
        RECT 273.560 41.060 273.730 41.250 ;
        RECT 274.020 41.060 274.190 41.250 ;
        RECT 276.780 41.040 276.950 41.230 ;
        RECT 277.695 41.090 277.815 41.200 ;
        RECT 278.625 41.040 278.795 41.250 ;
        RECT 282.300 41.040 282.470 41.230 ;
        RECT 285.520 41.060 285.690 41.250 ;
        RECT 285.980 41.060 286.150 41.250 ;
        RECT 287.820 41.040 287.990 41.230 ;
        RECT 289.670 41.095 289.830 41.205 ;
        RECT 290.580 41.040 290.750 41.230 ;
        RECT 291.505 41.040 291.675 41.230 ;
        RECT 292.880 41.060 293.050 41.250 ;
        RECT 293.340 41.060 293.510 41.250 ;
        RECT 297.480 41.040 297.650 41.250 ;
        RECT 299.315 41.090 299.435 41.200 ;
        RECT 301.160 41.060 301.330 41.250 ;
        RECT 301.615 41.090 301.735 41.200 ;
        RECT 302.080 41.060 302.250 41.250 ;
        RECT 304.390 41.095 304.550 41.205 ;
        RECT 305.300 41.060 305.470 41.250 ;
        RECT 308.060 41.060 308.230 41.250 ;
        RECT 308.520 41.040 308.690 41.230 ;
        RECT 308.990 41.085 309.150 41.195 ;
        RECT 310.820 41.040 310.990 41.250 ;
        RECT 162.100 40.230 163.470 41.040 ;
        RECT 164.400 40.360 173.590 41.040 ;
        RECT 168.910 40.140 169.840 40.360 ;
        RECT 172.670 40.130 173.590 40.360 ;
        RECT 173.600 40.360 182.790 41.040 ;
        RECT 182.895 40.360 186.360 41.040 ;
        RECT 173.600 40.130 174.520 40.360 ;
        RECT 177.350 40.140 178.280 40.360 ;
        RECT 182.895 40.130 183.815 40.360 ;
        RECT 186.480 40.260 187.850 41.040 ;
        RECT 187.870 40.170 188.300 40.955 ;
        RECT 188.320 40.230 189.690 41.040 ;
        RECT 189.700 40.260 191.070 41.040 ;
        RECT 191.080 40.260 192.450 41.040 ;
        RECT 192.460 40.230 193.830 41.040 ;
        RECT 193.840 40.360 197.740 41.040 ;
        RECT 198.075 40.360 201.540 41.040 ;
        RECT 193.840 40.130 194.770 40.360 ;
        RECT 198.075 40.130 198.995 40.360 ;
        RECT 201.660 40.230 203.030 41.040 ;
        RECT 203.050 40.130 204.400 41.040 ;
        RECT 204.420 40.360 213.610 41.040 ;
        RECT 208.930 40.140 209.860 40.360 ;
        RECT 212.690 40.130 213.610 40.360 ;
        RECT 213.630 40.170 214.060 40.955 ;
        RECT 214.080 40.230 219.590 41.040 ;
        RECT 219.600 40.260 220.970 41.040 ;
        RECT 220.980 40.260 222.350 41.040 ;
        RECT 222.360 40.360 226.260 41.040 ;
        RECT 222.360 40.130 223.290 40.360 ;
        RECT 226.960 40.260 228.330 41.040 ;
        RECT 228.340 40.360 232.240 41.040 ;
        RECT 232.480 40.360 236.380 41.040 ;
        RECT 228.340 40.130 229.270 40.360 ;
        RECT 232.480 40.130 233.410 40.360 ;
        RECT 236.620 40.230 239.370 41.040 ;
        RECT 239.390 40.170 239.820 40.955 ;
        RECT 240.410 40.360 243.875 41.040 ;
        RECT 242.955 40.130 243.875 40.360 ;
        RECT 244.440 40.360 248.340 41.040 ;
        RECT 248.580 40.360 257.770 41.040 ;
        RECT 244.440 40.130 245.370 40.360 ;
        RECT 253.090 40.140 254.020 40.360 ;
        RECT 256.850 40.130 257.770 40.360 ;
        RECT 257.875 40.360 261.340 41.040 ;
        RECT 261.555 40.360 265.020 41.040 ;
        RECT 257.875 40.130 258.795 40.360 ;
        RECT 261.555 40.130 262.475 40.360 ;
        RECT 265.150 40.170 265.580 40.955 ;
        RECT 265.600 40.230 267.430 41.040 ;
        RECT 267.440 40.360 276.630 41.040 ;
        RECT 271.950 40.140 272.880 40.360 ;
        RECT 275.710 40.130 276.630 40.360 ;
        RECT 276.640 40.230 278.470 41.040 ;
        RECT 278.480 40.130 282.135 41.040 ;
        RECT 282.160 40.230 287.670 41.040 ;
        RECT 287.680 40.230 289.050 41.040 ;
        RECT 289.060 40.360 290.890 41.040 ;
        RECT 289.060 40.130 290.405 40.360 ;
        RECT 290.910 40.170 291.340 40.955 ;
        RECT 291.360 40.130 297.070 41.040 ;
        RECT 297.340 40.230 299.170 41.040 ;
        RECT 299.640 40.360 308.830 41.040 ;
        RECT 299.640 40.130 300.560 40.360 ;
        RECT 303.390 40.140 304.320 40.360 ;
        RECT 309.760 40.230 311.130 41.040 ;
      LAYER nwell ;
        RECT 161.905 37.010 311.325 39.840 ;
      LAYER pwell ;
        RECT 162.100 35.810 163.470 36.620 ;
        RECT 163.480 35.810 165.310 36.620 ;
        RECT 170.290 36.490 171.220 36.710 ;
        RECT 174.050 36.490 174.970 36.720 ;
        RECT 165.780 35.810 174.970 36.490 ;
        RECT 174.990 35.895 175.420 36.680 ;
        RECT 179.560 36.490 180.490 36.720 ;
        RECT 176.590 35.810 180.490 36.490 ;
        RECT 180.595 36.490 181.515 36.720 ;
        RECT 180.595 35.810 184.060 36.490 ;
        RECT 184.180 35.810 186.930 36.620 ;
        RECT 191.450 36.490 192.380 36.710 ;
        RECT 195.210 36.490 196.130 36.720 ;
        RECT 186.940 35.810 196.130 36.490 ;
        RECT 197.155 36.490 198.075 36.720 ;
        RECT 197.155 35.810 200.620 36.490 ;
        RECT 200.750 35.895 201.180 36.680 ;
        RECT 201.200 35.810 204.870 36.620 ;
        RECT 210.310 36.490 211.240 36.710 ;
        RECT 214.070 36.490 214.990 36.720 ;
        RECT 205.800 35.810 214.990 36.490 ;
        RECT 215.000 35.810 220.510 36.620 ;
        RECT 220.520 35.810 221.890 36.590 ;
        RECT 221.995 36.490 222.915 36.720 ;
        RECT 221.995 35.810 225.460 36.490 ;
        RECT 226.510 35.895 226.940 36.680 ;
        RECT 227.055 36.490 227.975 36.720 ;
        RECT 230.640 36.490 231.570 36.720 ;
        RECT 227.055 35.810 230.520 36.490 ;
        RECT 230.640 35.810 234.540 36.490 ;
        RECT 162.240 35.600 162.410 35.810 ;
        RECT 163.620 35.600 163.790 35.810 ;
        RECT 165.455 35.650 165.575 35.760 ;
        RECT 165.920 35.620 166.090 35.810 ;
        RECT 167.300 35.600 167.470 35.790 ;
        RECT 175.590 35.655 175.750 35.765 ;
        RECT 176.775 35.600 176.945 35.790 ;
        RECT 179.905 35.620 180.075 35.810 ;
        RECT 180.640 35.600 180.810 35.790 ;
        RECT 183.860 35.620 184.030 35.810 ;
        RECT 184.320 35.620 184.490 35.810 ;
        RECT 186.160 35.600 186.330 35.790 ;
        RECT 187.080 35.620 187.250 35.810 ;
        RECT 188.460 35.600 188.630 35.790 ;
        RECT 193.245 35.600 193.415 35.790 ;
        RECT 194.900 35.600 195.070 35.790 ;
        RECT 195.360 35.600 195.530 35.790 ;
        RECT 196.290 35.655 196.450 35.765 ;
        RECT 199.040 35.600 199.210 35.790 ;
        RECT 200.420 35.600 200.590 35.810 ;
        RECT 201.340 35.620 201.510 35.810 ;
        RECT 204.375 35.600 204.545 35.790 ;
        RECT 205.030 35.655 205.190 35.765 ;
        RECT 205.940 35.620 206.110 35.810 ;
        RECT 209.160 35.600 209.330 35.790 ;
        RECT 209.895 35.600 210.065 35.790 ;
        RECT 214.215 35.650 214.335 35.760 ;
        RECT 215.140 35.620 215.310 35.810 ;
        RECT 217.900 35.600 218.070 35.790 ;
        RECT 218.635 35.600 218.805 35.790 ;
        RECT 221.580 35.620 221.750 35.810 ;
        RECT 222.775 35.600 222.945 35.790 ;
        RECT 225.260 35.620 225.430 35.810 ;
        RECT 225.730 35.655 225.890 35.765 ;
        RECT 226.640 35.600 226.810 35.790 ;
        RECT 230.320 35.600 230.490 35.810 ;
        RECT 231.055 35.620 231.225 35.810 ;
        RECT 235.700 35.770 236.590 36.720 ;
        RECT 237.540 35.810 239.370 36.490 ;
        RECT 234.930 35.655 235.090 35.765 ;
        RECT 236.300 35.620 236.470 35.770 ;
        RECT 236.770 35.655 236.930 35.765 ;
        RECT 239.060 35.620 239.230 35.810 ;
        RECT 240.320 35.770 241.210 36.720 ;
        RECT 241.220 36.490 242.140 36.720 ;
        RECT 244.970 36.490 245.900 36.710 ;
        RECT 241.220 35.810 250.410 36.490 ;
        RECT 250.420 35.810 252.250 36.620 ;
        RECT 252.270 35.895 252.700 36.680 ;
        RECT 252.720 35.810 254.090 36.620 ;
        RECT 254.100 36.490 255.020 36.720 ;
        RECT 257.850 36.490 258.780 36.710 ;
        RECT 254.100 35.810 263.290 36.490 ;
        RECT 263.300 35.810 266.050 36.620 ;
        RECT 266.060 35.810 267.430 36.590 ;
        RECT 267.535 36.490 268.455 36.720 ;
        RECT 271.215 36.490 272.135 36.720 ;
        RECT 267.535 35.810 271.000 36.490 ;
        RECT 271.215 35.810 274.680 36.490 ;
        RECT 274.810 35.810 277.540 36.720 ;
        RECT 278.030 35.895 278.460 36.680 ;
        RECT 280.450 36.490 281.380 36.720 ;
        RECT 279.545 35.810 281.380 36.490 ;
        RECT 282.175 35.810 283.990 36.720 ;
        RECT 284.000 36.490 284.920 36.720 ;
        RECT 290.810 36.490 291.740 36.710 ;
        RECT 294.570 36.490 295.490 36.720 ;
        RECT 284.000 35.810 286.290 36.490 ;
        RECT 286.300 35.810 295.490 36.490 ;
        RECT 295.500 36.490 296.420 36.720 ;
        RECT 298.850 36.490 299.780 36.720 ;
        RECT 302.755 36.490 303.675 36.720 ;
        RECT 295.500 35.810 297.790 36.490 ;
        RECT 297.945 35.810 299.780 36.490 ;
        RECT 300.210 35.810 303.675 36.490 ;
        RECT 303.790 35.895 304.220 36.680 ;
        RECT 305.160 35.810 306.990 36.490 ;
        RECT 307.000 35.810 309.750 36.620 ;
        RECT 309.760 35.810 311.130 36.620 ;
        RECT 239.530 35.655 239.690 35.765 ;
        RECT 239.990 35.645 240.150 35.755 ;
        RECT 240.440 35.620 240.610 35.770 ;
        RECT 240.900 35.600 241.070 35.770 ;
        RECT 242.280 35.600 242.450 35.790 ;
        RECT 250.100 35.620 250.270 35.810 ;
        RECT 250.560 35.620 250.730 35.810 ;
        RECT 252.860 35.620 253.030 35.810 ;
        RECT 254.700 35.600 254.870 35.790 ;
        RECT 255.160 35.600 255.330 35.790 ;
        RECT 260.680 35.600 260.850 35.790 ;
        RECT 262.980 35.620 263.150 35.810 ;
        RECT 263.440 35.620 263.610 35.810 ;
        RECT 264.370 35.645 264.530 35.755 ;
        RECT 265.740 35.600 265.910 35.790 ;
        RECT 266.200 35.620 266.370 35.810 ;
        RECT 269.875 35.600 270.045 35.790 ;
        RECT 270.800 35.620 270.970 35.810 ;
        RECT 274.480 35.620 274.650 35.810 ;
        RECT 277.240 35.620 277.410 35.810 ;
        RECT 279.545 35.790 279.710 35.810 ;
        RECT 277.695 35.650 277.815 35.760 ;
        RECT 278.630 35.655 278.790 35.765 ;
        RECT 279.080 35.600 279.250 35.790 ;
        RECT 279.540 35.600 279.710 35.790 ;
        RECT 281.835 35.650 281.955 35.760 ;
        RECT 282.300 35.620 282.470 35.810 ;
        RECT 283.220 35.600 283.390 35.790 ;
        RECT 285.980 35.620 286.150 35.810 ;
        RECT 286.440 35.620 286.610 35.810 ;
        RECT 287.360 35.600 287.530 35.790 ;
        RECT 162.100 34.790 163.470 35.600 ;
        RECT 163.480 34.790 167.150 35.600 ;
        RECT 167.160 34.920 176.350 35.600 ;
        RECT 171.670 34.700 172.600 34.920 ;
        RECT 175.430 34.690 176.350 34.920 ;
        RECT 176.360 34.920 180.260 35.600 ;
        RECT 176.360 34.690 177.290 34.920 ;
        RECT 180.500 34.790 186.010 35.600 ;
        RECT 186.020 34.790 187.850 35.600 ;
        RECT 187.870 34.730 188.300 35.515 ;
        RECT 188.320 34.790 189.690 35.600 ;
        RECT 189.930 34.920 193.830 35.600 ;
        RECT 192.900 34.690 193.830 34.920 ;
        RECT 193.840 34.820 195.210 35.600 ;
        RECT 195.220 34.790 198.890 35.600 ;
        RECT 198.900 34.790 200.270 35.600 ;
        RECT 200.390 34.920 203.855 35.600 ;
        RECT 202.935 34.690 203.855 34.920 ;
        RECT 203.960 34.920 207.860 35.600 ;
        RECT 203.960 34.690 204.890 34.920 ;
        RECT 208.100 34.820 209.470 35.600 ;
        RECT 209.480 34.920 213.380 35.600 ;
        RECT 209.480 34.690 210.410 34.920 ;
        RECT 213.630 34.730 214.060 35.515 ;
        RECT 214.635 34.920 218.100 35.600 ;
        RECT 218.220 34.920 222.120 35.600 ;
        RECT 222.360 34.920 226.260 35.600 ;
        RECT 226.610 34.920 230.075 35.600 ;
        RECT 230.180 34.920 239.370 35.600 ;
        RECT 214.635 34.690 215.555 34.920 ;
        RECT 218.220 34.690 219.150 34.920 ;
        RECT 222.360 34.690 223.290 34.920 ;
        RECT 229.155 34.690 230.075 34.920 ;
        RECT 234.690 34.700 235.620 34.920 ;
        RECT 238.450 34.690 239.370 34.920 ;
        RECT 239.390 34.730 239.820 35.515 ;
        RECT 240.760 34.820 242.130 35.600 ;
        RECT 242.140 34.920 251.330 35.600 ;
        RECT 246.650 34.700 247.580 34.920 ;
        RECT 250.410 34.690 251.330 34.920 ;
        RECT 251.435 34.920 254.900 35.600 ;
        RECT 251.435 34.690 252.355 34.920 ;
        RECT 255.020 34.790 260.530 35.600 ;
        RECT 260.540 34.790 264.210 35.600 ;
        RECT 265.150 34.730 265.580 35.515 ;
        RECT 265.600 34.790 268.350 35.600 ;
        RECT 268.360 34.690 270.190 35.600 ;
        RECT 270.200 34.920 279.390 35.600 ;
        RECT 279.510 34.920 282.975 35.600 ;
        RECT 270.200 34.690 271.120 34.920 ;
        RECT 273.950 34.700 274.880 34.920 ;
        RECT 282.055 34.690 282.975 34.920 ;
        RECT 283.080 34.790 284.910 35.600 ;
        RECT 284.930 34.920 287.670 35.600 ;
        RECT 287.680 35.570 288.625 35.600 ;
        RECT 290.580 35.570 290.750 35.790 ;
        RECT 292.420 35.600 292.590 35.790 ;
        RECT 292.875 35.650 292.995 35.760 ;
        RECT 296.560 35.600 296.730 35.790 ;
        RECT 297.030 35.645 297.190 35.755 ;
        RECT 297.480 35.620 297.650 35.810 ;
        RECT 297.945 35.790 298.110 35.810 ;
        RECT 297.940 35.620 298.110 35.790 ;
        RECT 299.320 35.600 299.490 35.790 ;
        RECT 300.240 35.620 300.410 35.810 ;
        RECT 304.390 35.655 304.550 35.765 ;
        RECT 306.680 35.620 306.850 35.810 ;
        RECT 307.140 35.620 307.310 35.810 ;
        RECT 308.520 35.600 308.690 35.790 ;
        RECT 308.990 35.645 309.150 35.755 ;
        RECT 310.820 35.600 310.990 35.810 ;
        RECT 287.680 35.370 290.750 35.570 ;
        RECT 287.680 34.890 290.890 35.370 ;
        RECT 287.680 34.690 288.625 34.890 ;
        RECT 289.960 34.690 290.890 34.890 ;
        RECT 290.910 34.730 291.340 35.515 ;
        RECT 291.370 34.690 292.720 35.600 ;
        RECT 293.295 34.920 296.760 35.600 ;
        RECT 297.800 34.920 299.630 35.600 ;
        RECT 299.640 34.920 308.830 35.600 ;
        RECT 293.295 34.690 294.215 34.920 ;
        RECT 299.640 34.690 300.560 34.920 ;
        RECT 303.390 34.700 304.320 34.920 ;
        RECT 309.760 34.790 311.130 35.600 ;
      LAYER nwell ;
        RECT 161.905 31.570 311.325 34.400 ;
      LAYER pwell ;
        RECT 162.100 30.370 163.470 31.180 ;
        RECT 163.480 30.370 168.990 31.180 ;
        RECT 169.000 30.370 170.370 31.150 ;
        RECT 170.840 30.370 172.210 31.150 ;
        RECT 172.220 30.370 174.970 31.180 ;
        RECT 174.990 30.455 175.420 31.240 ;
        RECT 175.440 31.050 176.370 31.280 ;
        RECT 179.580 31.050 180.500 31.280 ;
        RECT 183.330 31.050 184.260 31.270 ;
        RECT 193.290 31.050 194.220 31.270 ;
        RECT 197.050 31.050 197.970 31.280 ;
        RECT 175.440 30.370 179.340 31.050 ;
        RECT 179.580 30.370 188.770 31.050 ;
        RECT 188.780 30.370 197.970 31.050 ;
        RECT 197.980 30.370 200.730 31.180 ;
        RECT 200.750 30.455 201.180 31.240 ;
        RECT 201.200 30.370 202.570 31.180 ;
        RECT 205.340 31.050 206.260 31.280 ;
        RECT 209.090 31.050 210.020 31.270 ;
        RECT 202.590 30.370 205.330 31.050 ;
        RECT 205.340 30.370 214.530 31.050 ;
        RECT 214.540 30.370 215.910 31.150 ;
        RECT 215.920 30.370 217.290 31.150 ;
        RECT 221.810 31.050 222.740 31.270 ;
        RECT 225.570 31.050 226.490 31.280 ;
        RECT 217.300 30.370 226.490 31.050 ;
        RECT 226.510 30.455 226.940 31.240 ;
        RECT 226.960 31.050 227.880 31.280 ;
        RECT 230.710 31.050 231.640 31.270 ;
        RECT 226.960 30.370 236.150 31.050 ;
        RECT 236.170 30.370 238.910 31.050 ;
        RECT 238.920 30.370 242.590 31.180 ;
        RECT 242.600 30.370 243.970 31.180 ;
        RECT 243.980 30.370 245.350 31.150 ;
        RECT 245.360 31.050 246.290 31.280 ;
        RECT 245.360 30.370 249.260 31.050 ;
        RECT 249.500 30.370 252.250 31.180 ;
        RECT 252.270 30.455 252.700 31.240 ;
        RECT 252.720 30.370 255.470 31.180 ;
        RECT 259.010 31.050 259.940 31.280 ;
        RECT 255.950 30.370 258.690 31.050 ;
        RECT 259.010 30.370 260.845 31.050 ;
        RECT 261.000 30.370 264.670 31.180 ;
        RECT 265.140 31.050 266.060 31.280 ;
        RECT 268.890 31.050 269.820 31.270 ;
        RECT 276.995 31.050 277.915 31.280 ;
        RECT 265.140 30.370 274.330 31.050 ;
        RECT 274.450 30.370 277.915 31.050 ;
        RECT 278.030 30.455 278.460 31.240 ;
        RECT 278.480 31.050 279.410 31.280 ;
        RECT 278.480 30.370 282.380 31.050 ;
        RECT 282.620 30.370 283.970 31.280 ;
        RECT 284.000 30.370 285.370 31.180 ;
        RECT 285.380 31.050 286.300 31.280 ;
        RECT 289.130 31.050 290.060 31.270 ;
        RECT 294.580 31.050 295.500 31.280 ;
        RECT 298.330 31.050 299.260 31.270 ;
        RECT 285.380 30.370 294.570 31.050 ;
        RECT 294.580 30.370 303.770 31.050 ;
        RECT 303.790 30.455 304.220 31.240 ;
        RECT 304.335 31.050 305.255 31.280 ;
        RECT 304.335 30.370 307.800 31.050 ;
        RECT 307.920 30.370 309.750 31.180 ;
        RECT 309.760 30.370 311.130 31.180 ;
        RECT 162.240 30.160 162.410 30.370 ;
        RECT 163.620 30.180 163.790 30.370 ;
        RECT 165.000 30.160 165.170 30.350 ;
        RECT 165.460 30.160 165.630 30.350 ;
        RECT 170.060 30.180 170.230 30.370 ;
        RECT 170.515 30.210 170.635 30.320 ;
        RECT 170.980 30.160 171.150 30.350 ;
        RECT 171.900 30.180 172.070 30.370 ;
        RECT 172.360 30.180 172.530 30.370 ;
        RECT 175.855 30.180 176.025 30.370 ;
        RECT 176.500 30.160 176.670 30.350 ;
        RECT 182.020 30.160 182.190 30.350 ;
        RECT 185.695 30.210 185.815 30.320 ;
        RECT 186.160 30.160 186.330 30.350 ;
        RECT 187.535 30.210 187.655 30.320 ;
        RECT 188.460 30.160 188.630 30.370 ;
        RECT 188.920 30.180 189.090 30.370 ;
        RECT 195.545 30.160 195.715 30.350 ;
        RECT 196.280 30.160 196.450 30.350 ;
        RECT 198.120 30.180 198.290 30.370 ;
        RECT 199.040 30.160 199.210 30.350 ;
        RECT 201.340 30.180 201.510 30.370 ;
        RECT 205.020 30.180 205.190 30.370 ;
        RECT 208.250 30.205 208.410 30.315 ;
        RECT 212.565 30.160 212.735 30.350 ;
        RECT 213.295 30.210 213.415 30.320 ;
        RECT 214.220 30.160 214.390 30.370 ;
        RECT 215.600 30.180 215.770 30.370 ;
        RECT 216.980 30.180 217.150 30.370 ;
        RECT 217.440 30.180 217.610 30.370 ;
        RECT 223.420 30.160 223.590 30.350 ;
        RECT 228.950 30.205 229.110 30.315 ;
        RECT 229.860 30.160 230.030 30.350 ;
        RECT 231.235 30.210 231.355 30.320 ;
        RECT 231.975 30.160 232.145 30.350 ;
        RECT 235.840 30.160 236.010 30.370 ;
        RECT 238.600 30.180 238.770 30.370 ;
        RECT 239.060 30.180 239.230 30.370 ;
        RECT 239.980 30.160 240.150 30.350 ;
        RECT 242.740 30.180 242.910 30.370 ;
        RECT 245.040 30.180 245.210 30.370 ;
        RECT 245.500 30.160 245.670 30.350 ;
        RECT 245.775 30.180 245.945 30.370 ;
        RECT 249.640 30.180 249.810 30.370 ;
        RECT 251.020 30.160 251.190 30.350 ;
        RECT 252.860 30.180 253.030 30.370 ;
        RECT 255.615 30.210 255.735 30.320 ;
        RECT 256.540 30.160 256.710 30.350 ;
        RECT 258.380 30.180 258.550 30.370 ;
        RECT 260.680 30.350 260.845 30.370 ;
        RECT 260.680 30.180 260.850 30.350 ;
        RECT 261.140 30.180 261.310 30.370 ;
        RECT 262.060 30.160 262.230 30.350 ;
        RECT 264.815 30.210 264.935 30.320 ;
        RECT 265.740 30.160 265.910 30.350 ;
        RECT 267.575 30.210 267.695 30.320 ;
        RECT 268.040 30.160 268.210 30.350 ;
        RECT 274.020 30.180 274.190 30.370 ;
        RECT 274.480 30.180 274.650 30.370 ;
        RECT 277.245 30.160 277.415 30.350 ;
        RECT 278.895 30.180 279.065 30.370 ;
        RECT 280.925 30.160 281.095 30.350 ;
        RECT 283.685 30.180 283.855 30.370 ;
        RECT 284.140 30.180 284.310 30.370 ;
        RECT 284.600 30.160 284.770 30.350 ;
        RECT 290.130 30.205 290.290 30.315 ;
        RECT 291.500 30.160 291.670 30.350 ;
        RECT 294.260 30.320 294.430 30.370 ;
        RECT 294.255 30.210 294.430 30.320 ;
        RECT 294.260 30.180 294.430 30.210 ;
        RECT 295.640 30.160 295.810 30.350 ;
        RECT 296.100 30.160 296.270 30.350 ;
        RECT 303.460 30.180 303.630 30.370 ;
        RECT 307.600 30.180 307.770 30.370 ;
        RECT 308.060 30.180 308.230 30.370 ;
        RECT 308.520 30.160 308.690 30.350 ;
        RECT 308.990 30.205 309.150 30.315 ;
        RECT 310.820 30.160 310.990 30.370 ;
        RECT 162.100 29.350 163.470 30.160 ;
        RECT 163.480 29.480 165.310 30.160 ;
        RECT 163.480 29.250 164.825 29.480 ;
        RECT 165.320 29.350 170.830 30.160 ;
        RECT 170.840 29.350 176.350 30.160 ;
        RECT 176.360 29.350 181.870 30.160 ;
        RECT 181.880 29.350 185.550 30.160 ;
        RECT 186.020 29.380 187.390 30.160 ;
        RECT 187.870 29.290 188.300 30.075 ;
        RECT 188.320 29.350 191.990 30.160 ;
        RECT 192.230 29.480 196.130 30.160 ;
        RECT 195.200 29.250 196.130 29.480 ;
        RECT 196.140 29.350 198.890 30.160 ;
        RECT 198.900 29.480 208.090 30.160 ;
        RECT 209.250 29.480 213.150 30.160 ;
        RECT 203.410 29.260 204.340 29.480 ;
        RECT 207.170 29.250 208.090 29.480 ;
        RECT 212.220 29.250 213.150 29.480 ;
        RECT 213.630 29.290 214.060 30.075 ;
        RECT 214.080 29.480 223.270 30.160 ;
        RECT 218.590 29.260 219.520 29.480 ;
        RECT 222.350 29.250 223.270 29.480 ;
        RECT 223.280 29.350 228.790 30.160 ;
        RECT 229.720 29.380 231.090 30.160 ;
        RECT 231.560 29.480 235.460 30.160 ;
        RECT 231.560 29.250 232.490 29.480 ;
        RECT 235.700 29.350 239.370 30.160 ;
        RECT 239.390 29.290 239.820 30.075 ;
        RECT 239.840 29.350 245.350 30.160 ;
        RECT 245.360 29.350 250.870 30.160 ;
        RECT 250.880 29.350 256.390 30.160 ;
        RECT 256.400 29.350 261.910 30.160 ;
        RECT 261.920 29.350 264.670 30.160 ;
        RECT 265.150 29.290 265.580 30.075 ;
        RECT 265.600 29.350 267.430 30.160 ;
        RECT 267.900 29.480 277.090 30.160 ;
        RECT 272.410 29.260 273.340 29.480 ;
        RECT 276.170 29.250 277.090 29.480 ;
        RECT 277.100 29.250 280.770 30.160 ;
        RECT 280.780 29.250 284.450 30.160 ;
        RECT 284.460 29.350 289.970 30.160 ;
        RECT 290.910 29.290 291.340 30.075 ;
        RECT 291.360 29.350 294.110 30.160 ;
        RECT 294.590 29.250 295.940 30.160 ;
        RECT 295.960 29.350 299.630 30.160 ;
        RECT 299.640 29.480 308.830 30.160 ;
        RECT 299.640 29.250 300.560 29.480 ;
        RECT 303.390 29.260 304.320 29.480 ;
        RECT 309.760 29.350 311.130 30.160 ;
      LAYER nwell ;
        RECT 161.905 26.130 311.325 28.960 ;
      LAYER pwell ;
        RECT 162.100 24.930 163.470 25.740 ;
        RECT 163.480 24.930 168.990 25.740 ;
        RECT 169.000 24.930 174.510 25.740 ;
        RECT 174.990 25.015 175.420 25.800 ;
        RECT 175.440 24.930 180.950 25.740 ;
        RECT 180.960 24.930 186.470 25.740 ;
        RECT 186.480 24.930 188.310 25.740 ;
        RECT 188.320 25.610 189.250 25.840 ;
        RECT 188.320 24.930 192.220 25.610 ;
        RECT 192.460 24.930 197.970 25.740 ;
        RECT 197.980 24.930 200.730 25.740 ;
        RECT 200.750 25.015 201.180 25.800 ;
        RECT 201.660 24.930 203.030 25.710 ;
        RECT 203.040 24.930 204.410 25.740 ;
        RECT 204.420 24.930 207.160 25.610 ;
        RECT 207.180 24.930 212.690 25.740 ;
        RECT 212.700 24.930 218.210 25.740 ;
        RECT 218.220 24.930 223.730 25.740 ;
        RECT 223.740 24.930 226.490 25.740 ;
        RECT 226.510 25.015 226.940 25.800 ;
        RECT 226.960 24.930 232.470 25.740 ;
        RECT 232.480 24.930 237.990 25.740 ;
        RECT 238.000 24.930 243.510 25.740 ;
        RECT 243.520 24.930 249.030 25.740 ;
        RECT 249.040 24.930 251.790 25.740 ;
        RECT 252.270 25.015 252.700 25.800 ;
        RECT 252.720 24.930 258.230 25.740 ;
        RECT 258.240 24.930 263.750 25.740 ;
        RECT 263.760 24.930 269.270 25.740 ;
        RECT 269.280 24.930 271.110 25.740 ;
        RECT 271.130 24.930 273.870 25.610 ;
        RECT 273.880 24.930 277.550 25.740 ;
        RECT 278.030 25.015 278.460 25.800 ;
        RECT 278.480 24.930 283.990 25.740 ;
        RECT 284.000 24.930 289.510 25.740 ;
        RECT 289.520 24.930 295.030 25.740 ;
        RECT 295.040 24.930 300.550 25.740 ;
        RECT 300.560 24.930 303.310 25.740 ;
        RECT 303.790 25.015 304.220 25.800 ;
        RECT 304.240 24.930 309.750 25.740 ;
        RECT 309.760 24.930 311.130 25.740 ;
        RECT 162.240 24.720 162.410 24.930 ;
        RECT 163.620 24.720 163.790 24.930 ;
        RECT 169.140 24.720 169.310 24.930 ;
        RECT 174.660 24.880 174.830 24.910 ;
        RECT 174.655 24.770 174.830 24.880 ;
        RECT 174.660 24.720 174.830 24.770 ;
        RECT 175.580 24.740 175.750 24.930 ;
        RECT 180.180 24.720 180.350 24.910 ;
        RECT 181.100 24.740 181.270 24.930 ;
        RECT 185.700 24.720 185.870 24.910 ;
        RECT 186.620 24.740 186.790 24.930 ;
        RECT 187.535 24.770 187.655 24.880 ;
        RECT 188.460 24.720 188.630 24.910 ;
        RECT 188.735 24.740 188.905 24.930 ;
        RECT 192.600 24.740 192.770 24.930 ;
        RECT 193.980 24.720 194.150 24.910 ;
        RECT 198.120 24.740 198.290 24.930 ;
        RECT 199.500 24.720 199.670 24.910 ;
        RECT 201.335 24.770 201.455 24.880 ;
        RECT 202.720 24.740 202.890 24.930 ;
        RECT 203.180 24.740 203.350 24.930 ;
        RECT 204.560 24.740 204.730 24.930 ;
        RECT 205.020 24.720 205.190 24.910 ;
        RECT 207.320 24.740 207.490 24.930 ;
        RECT 210.540 24.720 210.710 24.910 ;
        RECT 212.840 24.740 213.010 24.930 ;
        RECT 213.295 24.770 213.415 24.880 ;
        RECT 214.220 24.720 214.390 24.910 ;
        RECT 218.360 24.740 218.530 24.930 ;
        RECT 219.740 24.720 219.910 24.910 ;
        RECT 223.880 24.740 224.050 24.930 ;
        RECT 225.260 24.720 225.430 24.910 ;
        RECT 227.100 24.740 227.270 24.930 ;
        RECT 230.780 24.720 230.950 24.910 ;
        RECT 232.620 24.740 232.790 24.930 ;
        RECT 236.300 24.720 236.470 24.910 ;
        RECT 238.140 24.740 238.310 24.930 ;
        RECT 239.055 24.770 239.175 24.880 ;
        RECT 239.980 24.720 240.150 24.910 ;
        RECT 243.660 24.740 243.830 24.930 ;
        RECT 245.500 24.720 245.670 24.910 ;
        RECT 249.180 24.740 249.350 24.930 ;
        RECT 251.020 24.720 251.190 24.910 ;
        RECT 251.935 24.770 252.055 24.880 ;
        RECT 252.860 24.740 253.030 24.930 ;
        RECT 256.540 24.720 256.710 24.910 ;
        RECT 258.380 24.740 258.550 24.930 ;
        RECT 262.060 24.720 262.230 24.910 ;
        RECT 263.900 24.740 264.070 24.930 ;
        RECT 264.815 24.770 264.935 24.880 ;
        RECT 265.740 24.720 265.910 24.910 ;
        RECT 269.420 24.740 269.590 24.930 ;
        RECT 271.260 24.720 271.430 24.910 ;
        RECT 273.560 24.740 273.730 24.930 ;
        RECT 274.020 24.740 274.190 24.930 ;
        RECT 276.780 24.720 276.950 24.910 ;
        RECT 277.695 24.770 277.815 24.880 ;
        RECT 278.620 24.740 278.790 24.930 ;
        RECT 282.300 24.720 282.470 24.910 ;
        RECT 284.140 24.740 284.310 24.930 ;
        RECT 287.820 24.720 287.990 24.910 ;
        RECT 289.660 24.740 289.830 24.930 ;
        RECT 290.575 24.770 290.695 24.880 ;
        RECT 291.500 24.720 291.670 24.910 ;
        RECT 295.180 24.740 295.350 24.930 ;
        RECT 297.020 24.720 297.190 24.910 ;
        RECT 300.700 24.740 300.870 24.930 ;
        RECT 302.540 24.720 302.710 24.910 ;
        RECT 303.455 24.770 303.575 24.880 ;
        RECT 304.380 24.740 304.550 24.930 ;
        RECT 308.060 24.720 308.230 24.910 ;
        RECT 310.820 24.720 310.990 24.930 ;
        RECT 162.100 23.910 163.470 24.720 ;
        RECT 163.480 23.910 168.990 24.720 ;
        RECT 169.000 23.910 174.510 24.720 ;
        RECT 174.520 23.910 180.030 24.720 ;
        RECT 180.040 23.910 185.550 24.720 ;
        RECT 185.560 23.910 187.390 24.720 ;
        RECT 187.870 23.850 188.300 24.635 ;
        RECT 188.320 23.910 193.830 24.720 ;
        RECT 193.840 23.910 199.350 24.720 ;
        RECT 199.360 23.910 204.870 24.720 ;
        RECT 204.880 23.910 210.390 24.720 ;
        RECT 210.400 23.910 213.150 24.720 ;
        RECT 213.630 23.850 214.060 24.635 ;
        RECT 214.080 23.910 219.590 24.720 ;
        RECT 219.600 23.910 225.110 24.720 ;
        RECT 225.120 23.910 230.630 24.720 ;
        RECT 230.640 23.910 236.150 24.720 ;
        RECT 236.160 23.910 238.910 24.720 ;
        RECT 239.390 23.850 239.820 24.635 ;
        RECT 239.840 23.910 245.350 24.720 ;
        RECT 245.360 23.910 250.870 24.720 ;
        RECT 250.880 23.910 256.390 24.720 ;
        RECT 256.400 23.910 261.910 24.720 ;
        RECT 261.920 23.910 264.670 24.720 ;
        RECT 265.150 23.850 265.580 24.635 ;
        RECT 265.600 23.910 271.110 24.720 ;
        RECT 271.120 23.910 276.630 24.720 ;
        RECT 276.640 23.910 282.150 24.720 ;
        RECT 282.160 23.910 287.670 24.720 ;
        RECT 287.680 23.910 290.430 24.720 ;
        RECT 290.910 23.850 291.340 24.635 ;
        RECT 291.360 23.910 296.870 24.720 ;
        RECT 296.880 23.910 302.390 24.720 ;
        RECT 302.400 23.910 307.910 24.720 ;
        RECT 307.920 23.910 309.750 24.720 ;
        RECT 309.760 23.910 311.130 24.720 ;
      LAYER nwell ;
        RECT 161.905 20.690 311.325 23.520 ;
      LAYER pwell ;
        RECT 162.100 19.490 163.470 20.300 ;
        RECT 163.480 19.490 168.990 20.300 ;
        RECT 169.000 19.490 174.510 20.300 ;
        RECT 174.990 19.575 175.420 20.360 ;
        RECT 175.440 19.490 180.950 20.300 ;
        RECT 180.960 19.490 186.470 20.300 ;
        RECT 186.480 19.490 191.990 20.300 ;
        RECT 192.000 19.490 197.510 20.300 ;
        RECT 197.520 19.490 200.270 20.300 ;
        RECT 200.750 19.575 201.180 20.360 ;
        RECT 201.200 19.490 206.710 20.300 ;
        RECT 206.720 19.490 212.230 20.300 ;
        RECT 212.240 19.490 217.750 20.300 ;
        RECT 217.760 19.490 223.270 20.300 ;
        RECT 223.280 19.490 226.030 20.300 ;
        RECT 226.510 19.575 226.940 20.360 ;
        RECT 226.960 19.490 232.470 20.300 ;
        RECT 232.480 19.490 237.990 20.300 ;
        RECT 238.000 19.490 243.510 20.300 ;
        RECT 243.520 19.490 249.030 20.300 ;
        RECT 249.040 19.490 251.790 20.300 ;
        RECT 252.270 19.575 252.700 20.360 ;
        RECT 252.720 19.490 258.230 20.300 ;
        RECT 258.240 19.490 263.750 20.300 ;
        RECT 263.760 19.490 269.270 20.300 ;
        RECT 269.280 19.490 274.790 20.300 ;
        RECT 274.800 19.490 277.550 20.300 ;
        RECT 278.030 19.575 278.460 20.360 ;
        RECT 278.480 19.490 283.990 20.300 ;
        RECT 284.000 19.490 289.510 20.300 ;
        RECT 289.520 19.490 295.030 20.300 ;
        RECT 295.040 19.490 300.550 20.300 ;
        RECT 300.560 19.490 303.310 20.300 ;
        RECT 303.790 19.575 304.220 20.360 ;
        RECT 304.240 19.490 309.750 20.300 ;
        RECT 309.760 19.490 311.130 20.300 ;
        RECT 162.240 19.280 162.410 19.490 ;
        RECT 163.620 19.280 163.790 19.490 ;
        RECT 169.140 19.280 169.310 19.490 ;
        RECT 174.660 19.440 174.830 19.470 ;
        RECT 174.655 19.330 174.830 19.440 ;
        RECT 174.660 19.280 174.830 19.330 ;
        RECT 175.580 19.300 175.750 19.490 ;
        RECT 180.180 19.280 180.350 19.470 ;
        RECT 181.100 19.300 181.270 19.490 ;
        RECT 185.700 19.280 185.870 19.470 ;
        RECT 186.620 19.300 186.790 19.490 ;
        RECT 187.535 19.330 187.655 19.440 ;
        RECT 188.460 19.280 188.630 19.470 ;
        RECT 192.140 19.300 192.310 19.490 ;
        RECT 193.980 19.280 194.150 19.470 ;
        RECT 197.660 19.300 197.830 19.490 ;
        RECT 199.500 19.280 199.670 19.470 ;
        RECT 200.415 19.330 200.535 19.440 ;
        RECT 201.340 19.300 201.510 19.490 ;
        RECT 205.020 19.280 205.190 19.470 ;
        RECT 206.860 19.300 207.030 19.490 ;
        RECT 210.540 19.280 210.710 19.470 ;
        RECT 212.380 19.300 212.550 19.490 ;
        RECT 213.295 19.330 213.415 19.440 ;
        RECT 214.220 19.280 214.390 19.470 ;
        RECT 217.900 19.300 218.070 19.490 ;
        RECT 219.740 19.280 219.910 19.470 ;
        RECT 223.420 19.300 223.590 19.490 ;
        RECT 225.260 19.280 225.430 19.470 ;
        RECT 226.175 19.330 226.295 19.440 ;
        RECT 227.100 19.300 227.270 19.490 ;
        RECT 230.780 19.280 230.950 19.470 ;
        RECT 232.620 19.300 232.790 19.490 ;
        RECT 236.300 19.280 236.470 19.470 ;
        RECT 238.140 19.300 238.310 19.490 ;
        RECT 239.055 19.330 239.175 19.440 ;
        RECT 239.980 19.280 240.150 19.470 ;
        RECT 243.660 19.300 243.830 19.490 ;
        RECT 245.500 19.280 245.670 19.470 ;
        RECT 249.180 19.300 249.350 19.490 ;
        RECT 251.020 19.280 251.190 19.470 ;
        RECT 251.935 19.330 252.055 19.440 ;
        RECT 252.860 19.300 253.030 19.490 ;
        RECT 256.540 19.280 256.710 19.470 ;
        RECT 258.380 19.300 258.550 19.490 ;
        RECT 262.060 19.280 262.230 19.470 ;
        RECT 263.900 19.300 264.070 19.490 ;
        RECT 264.815 19.330 264.935 19.440 ;
        RECT 265.740 19.280 265.910 19.470 ;
        RECT 269.420 19.300 269.590 19.490 ;
        RECT 271.260 19.280 271.430 19.470 ;
        RECT 274.940 19.300 275.110 19.490 ;
        RECT 276.780 19.280 276.950 19.470 ;
        RECT 277.695 19.330 277.815 19.440 ;
        RECT 278.620 19.300 278.790 19.490 ;
        RECT 282.300 19.280 282.470 19.470 ;
        RECT 284.140 19.300 284.310 19.490 ;
        RECT 287.820 19.280 287.990 19.470 ;
        RECT 289.660 19.300 289.830 19.490 ;
        RECT 290.575 19.330 290.695 19.440 ;
        RECT 291.500 19.280 291.670 19.470 ;
        RECT 295.180 19.300 295.350 19.490 ;
        RECT 297.020 19.280 297.190 19.470 ;
        RECT 300.700 19.300 300.870 19.490 ;
        RECT 302.540 19.280 302.710 19.470 ;
        RECT 303.455 19.330 303.575 19.440 ;
        RECT 304.380 19.300 304.550 19.490 ;
        RECT 308.060 19.280 308.230 19.470 ;
        RECT 310.820 19.280 310.990 19.490 ;
        RECT 162.100 18.470 163.470 19.280 ;
        RECT 163.480 18.470 168.990 19.280 ;
        RECT 169.000 18.470 174.510 19.280 ;
        RECT 174.520 18.470 180.030 19.280 ;
        RECT 180.040 18.470 185.550 19.280 ;
        RECT 185.560 18.470 187.390 19.280 ;
        RECT 187.870 18.410 188.300 19.195 ;
        RECT 188.320 18.470 193.830 19.280 ;
        RECT 193.840 18.470 199.350 19.280 ;
        RECT 199.360 18.470 204.870 19.280 ;
        RECT 204.880 18.470 210.390 19.280 ;
        RECT 210.400 18.470 213.150 19.280 ;
        RECT 213.630 18.410 214.060 19.195 ;
        RECT 214.080 18.470 219.590 19.280 ;
        RECT 219.600 18.470 225.110 19.280 ;
        RECT 225.120 18.470 230.630 19.280 ;
        RECT 230.640 18.470 236.150 19.280 ;
        RECT 236.160 18.470 238.910 19.280 ;
        RECT 239.390 18.410 239.820 19.195 ;
        RECT 239.840 18.470 245.350 19.280 ;
        RECT 245.360 18.470 250.870 19.280 ;
        RECT 250.880 18.470 256.390 19.280 ;
        RECT 256.400 18.470 261.910 19.280 ;
        RECT 261.920 18.470 264.670 19.280 ;
        RECT 265.150 18.410 265.580 19.195 ;
        RECT 265.600 18.470 271.110 19.280 ;
        RECT 271.120 18.470 276.630 19.280 ;
        RECT 276.640 18.470 282.150 19.280 ;
        RECT 282.160 18.470 287.670 19.280 ;
        RECT 287.680 18.470 290.430 19.280 ;
        RECT 290.910 18.410 291.340 19.195 ;
        RECT 291.360 18.470 296.870 19.280 ;
        RECT 296.880 18.470 302.390 19.280 ;
        RECT 302.400 18.470 307.910 19.280 ;
        RECT 307.920 18.470 309.750 19.280 ;
        RECT 309.760 18.470 311.130 19.280 ;
      LAYER nwell ;
        RECT 161.905 15.250 311.325 18.080 ;
      LAYER pwell ;
        RECT 162.100 14.050 163.470 14.860 ;
        RECT 163.480 14.050 168.990 14.860 ;
        RECT 169.000 14.050 174.510 14.860 ;
        RECT 174.990 14.135 175.420 14.920 ;
        RECT 175.440 14.050 180.950 14.860 ;
        RECT 180.960 14.050 186.470 14.860 ;
        RECT 186.480 14.050 187.850 14.860 ;
        RECT 187.870 14.135 188.300 14.920 ;
        RECT 188.320 14.050 193.830 14.860 ;
        RECT 193.840 14.050 199.350 14.860 ;
        RECT 199.360 14.050 200.730 14.860 ;
        RECT 200.750 14.135 201.180 14.920 ;
        RECT 201.200 14.050 206.710 14.860 ;
        RECT 206.720 14.050 212.230 14.860 ;
        RECT 212.240 14.050 213.610 14.860 ;
        RECT 213.630 14.135 214.060 14.920 ;
        RECT 214.080 14.050 219.590 14.860 ;
        RECT 219.600 14.050 225.110 14.860 ;
        RECT 225.120 14.050 226.490 14.860 ;
        RECT 226.510 14.135 226.940 14.920 ;
        RECT 226.960 14.050 232.470 14.860 ;
        RECT 232.480 14.050 237.990 14.860 ;
        RECT 238.000 14.050 239.370 14.860 ;
        RECT 239.390 14.135 239.820 14.920 ;
        RECT 239.840 14.050 245.350 14.860 ;
        RECT 245.360 14.050 250.870 14.860 ;
        RECT 250.880 14.050 252.250 14.860 ;
        RECT 252.270 14.135 252.700 14.920 ;
        RECT 252.720 14.050 258.230 14.860 ;
        RECT 258.240 14.050 263.750 14.860 ;
        RECT 263.760 14.050 265.130 14.860 ;
        RECT 265.150 14.135 265.580 14.920 ;
        RECT 265.600 14.050 271.110 14.860 ;
        RECT 271.120 14.050 276.630 14.860 ;
        RECT 276.640 14.050 278.010 14.860 ;
        RECT 278.030 14.135 278.460 14.920 ;
        RECT 278.480 14.050 283.990 14.860 ;
        RECT 284.000 14.050 289.510 14.860 ;
        RECT 289.520 14.050 290.890 14.860 ;
        RECT 290.910 14.135 291.340 14.920 ;
        RECT 291.360 14.050 296.870 14.860 ;
        RECT 296.880 14.050 302.390 14.860 ;
        RECT 302.400 14.050 303.770 14.860 ;
        RECT 303.790 14.135 304.220 14.920 ;
        RECT 304.240 14.050 309.750 14.860 ;
        RECT 309.760 14.050 311.130 14.860 ;
        RECT 162.240 13.860 162.410 14.050 ;
        RECT 163.620 13.860 163.790 14.050 ;
        RECT 169.140 13.860 169.310 14.050 ;
        RECT 174.655 13.890 174.775 14.000 ;
        RECT 175.580 13.860 175.750 14.050 ;
        RECT 181.100 13.860 181.270 14.050 ;
        RECT 186.620 13.860 186.790 14.050 ;
        RECT 188.460 13.860 188.630 14.050 ;
        RECT 193.980 13.860 194.150 14.050 ;
        RECT 199.500 13.860 199.670 14.050 ;
        RECT 201.340 13.860 201.510 14.050 ;
        RECT 206.860 13.860 207.030 14.050 ;
        RECT 212.380 13.860 212.550 14.050 ;
        RECT 214.220 13.860 214.390 14.050 ;
        RECT 219.740 13.860 219.910 14.050 ;
        RECT 225.260 13.860 225.430 14.050 ;
        RECT 227.100 13.860 227.270 14.050 ;
        RECT 232.620 13.860 232.790 14.050 ;
        RECT 238.140 13.860 238.310 14.050 ;
        RECT 239.980 13.860 240.150 14.050 ;
        RECT 245.500 13.860 245.670 14.050 ;
        RECT 251.020 13.860 251.190 14.050 ;
        RECT 252.860 13.860 253.030 14.050 ;
        RECT 258.380 13.860 258.550 14.050 ;
        RECT 263.900 13.860 264.070 14.050 ;
        RECT 265.740 13.860 265.910 14.050 ;
        RECT 271.260 13.860 271.430 14.050 ;
        RECT 276.780 13.860 276.950 14.050 ;
        RECT 278.620 13.860 278.790 14.050 ;
        RECT 284.140 13.860 284.310 14.050 ;
        RECT 289.660 13.860 289.830 14.050 ;
        RECT 291.500 13.860 291.670 14.050 ;
        RECT 297.020 13.860 297.190 14.050 ;
        RECT 302.540 13.860 302.710 14.050 ;
        RECT 304.380 13.860 304.550 14.050 ;
        RECT 310.820 13.860 310.990 14.050 ;
      LAYER nwell ;
        RECT 3.250 3.250 156.750 5.750 ;
      LAYER li1 ;
        RECT 4.300 222.030 102.625 222.430 ;
        RECT 4.300 4.700 4.700 222.030 ;
        RECT 62.895 216.545 99.045 217.075 ;
        RECT 62.895 213.695 63.425 216.545 ;
        RECT 63.925 215.855 80.385 216.025 ;
        RECT 63.925 214.385 64.155 215.855 ;
        RECT 80.155 214.385 80.385 215.855 ;
        RECT 63.925 214.215 80.385 214.385 ;
        RECT 80.885 213.695 81.055 216.545 ;
        RECT 81.555 215.855 98.015 216.025 ;
        RECT 81.555 214.385 81.785 215.855 ;
        RECT 97.785 214.385 98.015 215.855 ;
        RECT 81.555 214.215 98.015 214.385 ;
        RECT 98.515 213.695 99.045 216.545 ;
        RECT 62.895 213.525 99.045 213.695 ;
        RECT 9.325 211.690 45.335 211.860 ;
        RECT 9.325 201.840 9.495 211.690 ;
        RECT 10.225 211.000 18.225 211.170 ;
        RECT 18.515 211.000 26.515 211.170 ;
        RECT 9.995 202.745 10.165 210.785 ;
        RECT 18.285 202.745 18.455 210.785 ;
        RECT 26.575 202.745 26.745 210.785 ;
        RECT 10.225 202.360 18.225 202.530 ;
        RECT 18.515 202.360 26.515 202.530 ;
        RECT 27.245 201.840 27.415 211.690 ;
        RECT 28.145 211.000 36.145 211.170 ;
        RECT 36.435 211.000 44.435 211.170 ;
        RECT 27.915 202.745 28.085 210.785 ;
        RECT 36.205 202.745 36.375 210.785 ;
        RECT 44.495 202.745 44.665 210.785 ;
        RECT 28.145 202.360 36.145 202.530 ;
        RECT 36.435 202.360 44.435 202.530 ;
        RECT 45.165 201.840 45.335 211.690 ;
        RECT 62.895 210.675 63.425 213.525 ;
        RECT 64.155 212.835 80.155 213.005 ;
        RECT 63.925 211.580 64.095 212.620 ;
        RECT 80.215 211.580 80.385 212.620 ;
        RECT 64.155 211.195 80.155 211.365 ;
        RECT 80.885 210.675 81.055 213.525 ;
        RECT 81.785 212.835 97.785 213.005 ;
        RECT 81.555 211.580 81.725 212.620 ;
        RECT 97.845 211.580 98.015 212.620 ;
        RECT 81.785 211.195 97.785 211.365 ;
        RECT 98.515 210.675 99.045 213.525 ;
        RECT 62.895 210.505 99.045 210.675 ;
        RECT 9.325 201.670 45.335 201.840 ;
        RECT 9.325 191.820 9.495 201.670 ;
        RECT 10.225 200.980 18.225 201.150 ;
        RECT 18.515 200.980 26.515 201.150 ;
        RECT 9.995 192.725 10.165 200.765 ;
        RECT 18.285 192.725 18.455 200.765 ;
        RECT 26.575 192.725 26.745 200.765 ;
        RECT 10.225 192.340 18.225 192.510 ;
        RECT 18.515 192.340 26.515 192.510 ;
        RECT 27.245 191.820 27.415 201.670 ;
        RECT 28.145 200.980 36.145 201.150 ;
        RECT 36.435 200.980 44.435 201.150 ;
        RECT 27.915 192.725 28.085 200.765 ;
        RECT 36.205 192.725 36.375 200.765 ;
        RECT 44.495 192.725 44.665 200.765 ;
        RECT 28.145 192.340 36.145 192.510 ;
        RECT 36.435 192.340 44.435 192.510 ;
        RECT 45.165 191.820 45.335 201.670 ;
        RECT 9.325 191.650 45.335 191.820 ;
        RECT 49.250 210.180 56.310 210.350 ;
        RECT 9.325 190.700 15.415 190.870 ;
        RECT 9.325 180.850 9.495 190.700 ;
        RECT 10.225 190.010 12.225 190.180 ;
        RECT 12.515 190.010 14.515 190.180 ;
        RECT 9.995 181.755 10.165 189.795 ;
        RECT 12.285 181.755 12.455 189.795 ;
        RECT 14.575 181.755 14.745 189.795 ;
        RECT 10.225 181.370 12.225 181.540 ;
        RECT 12.515 181.370 14.515 181.540 ;
        RECT 15.245 180.850 15.415 190.700 ;
        RECT 9.325 180.680 15.415 180.850 ;
        RECT 16.345 190.700 45.335 190.870 ;
        RECT 16.345 180.850 16.515 190.700 ;
        RECT 17.245 190.010 19.245 190.180 ;
        RECT 19.535 190.010 21.535 190.180 ;
        RECT 21.825 190.010 23.825 190.180 ;
        RECT 24.115 190.010 26.115 190.180 ;
        RECT 26.405 190.010 28.405 190.180 ;
        RECT 28.695 190.010 30.695 190.180 ;
        RECT 30.985 190.010 32.985 190.180 ;
        RECT 33.275 190.010 35.275 190.180 ;
        RECT 35.565 190.010 37.565 190.180 ;
        RECT 37.855 190.010 39.855 190.180 ;
        RECT 40.145 190.010 42.145 190.180 ;
        RECT 42.435 190.010 44.435 190.180 ;
        RECT 17.015 181.755 17.185 189.795 ;
        RECT 19.305 181.755 19.475 189.795 ;
        RECT 21.595 181.755 21.765 189.795 ;
        RECT 23.885 181.755 24.055 189.795 ;
        RECT 26.175 181.755 26.345 189.795 ;
        RECT 28.465 181.755 28.635 189.795 ;
        RECT 30.755 181.755 30.925 189.795 ;
        RECT 33.045 181.755 33.215 189.795 ;
        RECT 35.335 181.755 35.505 189.795 ;
        RECT 37.625 181.755 37.795 189.795 ;
        RECT 39.915 181.755 40.085 189.795 ;
        RECT 42.205 181.755 42.375 189.795 ;
        RECT 44.495 181.755 44.665 189.795 ;
        RECT 17.245 181.370 19.245 181.540 ;
        RECT 19.535 181.370 21.535 181.540 ;
        RECT 21.825 181.370 23.825 181.540 ;
        RECT 24.115 181.370 26.115 181.540 ;
        RECT 26.405 181.370 28.405 181.540 ;
        RECT 28.695 181.370 30.695 181.540 ;
        RECT 30.985 181.370 32.985 181.540 ;
        RECT 33.275 181.370 35.275 181.540 ;
        RECT 35.565 181.370 37.565 181.540 ;
        RECT 37.855 181.370 39.855 181.540 ;
        RECT 40.145 181.370 42.145 181.540 ;
        RECT 42.435 181.370 44.435 181.540 ;
        RECT 45.165 180.850 45.335 190.700 ;
        RECT 49.250 187.850 49.420 210.180 ;
        RECT 50.095 207.435 50.785 209.595 ;
        RECT 51.265 207.435 51.955 209.595 ;
        RECT 52.435 207.435 53.125 209.595 ;
        RECT 53.605 207.435 54.295 209.595 ;
        RECT 54.775 207.435 55.465 209.595 ;
        RECT 50.095 188.435 50.785 190.595 ;
        RECT 51.265 188.435 51.955 190.595 ;
        RECT 52.435 188.435 53.125 190.595 ;
        RECT 53.605 188.435 54.295 190.595 ;
        RECT 54.775 188.435 55.465 190.595 ;
        RECT 56.140 187.850 56.310 210.180 ;
        RECT 49.250 187.680 56.310 187.850 ;
        RECT 62.895 207.655 63.425 210.505 ;
        RECT 64.155 209.815 80.155 209.985 ;
        RECT 63.925 208.560 64.095 209.600 ;
        RECT 80.215 208.560 80.385 209.600 ;
        RECT 64.155 208.175 80.155 208.345 ;
        RECT 80.885 207.655 81.055 210.505 ;
        RECT 81.785 209.815 97.785 209.985 ;
        RECT 81.555 208.560 81.725 209.600 ;
        RECT 97.845 208.560 98.015 209.600 ;
        RECT 81.785 208.175 97.785 208.345 ;
        RECT 98.515 207.655 99.045 210.505 ;
        RECT 62.895 207.485 99.045 207.655 ;
        RECT 62.895 204.635 63.425 207.485 ;
        RECT 64.155 206.795 80.155 206.965 ;
        RECT 63.925 205.540 64.095 206.580 ;
        RECT 80.215 205.540 80.385 206.580 ;
        RECT 64.155 205.155 80.155 205.325 ;
        RECT 80.885 204.635 81.055 207.485 ;
        RECT 81.785 206.795 97.785 206.965 ;
        RECT 81.555 205.540 81.725 206.580 ;
        RECT 97.845 205.540 98.015 206.580 ;
        RECT 81.785 205.155 97.785 205.325 ;
        RECT 98.515 204.635 99.045 207.485 ;
        RECT 62.895 204.465 99.045 204.635 ;
        RECT 62.895 201.615 63.425 204.465 ;
        RECT 64.155 203.775 80.155 203.945 ;
        RECT 63.925 202.520 64.095 203.560 ;
        RECT 80.215 202.520 80.385 203.560 ;
        RECT 64.155 202.135 80.155 202.305 ;
        RECT 80.885 201.615 81.055 204.465 ;
        RECT 81.785 203.775 97.785 203.945 ;
        RECT 81.555 202.520 81.725 203.560 ;
        RECT 97.845 202.520 98.015 203.560 ;
        RECT 81.785 202.135 97.785 202.305 ;
        RECT 98.515 201.615 99.045 204.465 ;
        RECT 62.895 201.445 99.045 201.615 ;
        RECT 62.895 198.595 63.425 201.445 ;
        RECT 64.155 200.755 80.155 200.925 ;
        RECT 63.925 199.500 64.095 200.540 ;
        RECT 80.215 199.500 80.385 200.540 ;
        RECT 64.155 199.115 80.155 199.285 ;
        RECT 80.885 198.595 81.055 201.445 ;
        RECT 81.785 200.755 97.785 200.925 ;
        RECT 81.555 199.500 81.725 200.540 ;
        RECT 97.845 199.500 98.015 200.540 ;
        RECT 81.785 199.115 97.785 199.285 ;
        RECT 98.515 198.595 99.045 201.445 ;
        RECT 62.895 198.425 99.045 198.595 ;
        RECT 62.895 195.575 63.425 198.425 ;
        RECT 64.155 197.735 80.155 197.905 ;
        RECT 63.925 196.480 64.095 197.520 ;
        RECT 80.215 196.480 80.385 197.520 ;
        RECT 64.155 196.095 80.155 196.265 ;
        RECT 80.885 195.575 81.055 198.425 ;
        RECT 81.785 197.735 97.785 197.905 ;
        RECT 81.555 196.480 81.725 197.520 ;
        RECT 97.845 196.480 98.015 197.520 ;
        RECT 81.785 196.095 97.785 196.265 ;
        RECT 98.515 195.575 99.045 198.425 ;
        RECT 62.895 195.405 99.045 195.575 ;
        RECT 62.895 192.555 63.425 195.405 ;
        RECT 64.155 194.715 80.155 194.885 ;
        RECT 63.925 193.460 64.095 194.500 ;
        RECT 80.215 193.460 80.385 194.500 ;
        RECT 64.155 193.075 80.155 193.245 ;
        RECT 80.885 192.555 81.055 195.405 ;
        RECT 81.785 194.715 97.785 194.885 ;
        RECT 81.555 193.460 81.725 194.500 ;
        RECT 97.845 193.460 98.015 194.500 ;
        RECT 81.785 193.075 97.785 193.245 ;
        RECT 98.515 192.555 99.045 195.405 ;
        RECT 62.895 192.385 99.045 192.555 ;
        RECT 62.895 189.535 63.425 192.385 ;
        RECT 64.155 191.695 80.155 191.865 ;
        RECT 63.925 190.440 64.095 191.480 ;
        RECT 80.215 190.440 80.385 191.480 ;
        RECT 64.155 190.055 80.155 190.225 ;
        RECT 80.885 189.535 81.055 192.385 ;
        RECT 81.785 191.695 97.785 191.865 ;
        RECT 81.555 190.440 81.725 191.480 ;
        RECT 97.845 190.440 98.015 191.480 ;
        RECT 81.785 190.055 97.785 190.225 ;
        RECT 98.515 189.535 99.045 192.385 ;
        RECT 62.895 189.365 99.045 189.535 ;
        RECT 16.345 180.680 45.335 180.850 ;
        RECT 62.895 186.515 63.425 189.365 ;
        RECT 64.155 188.675 80.155 188.845 ;
        RECT 63.925 187.420 64.095 188.460 ;
        RECT 80.215 187.420 80.385 188.460 ;
        RECT 64.155 187.035 80.155 187.205 ;
        RECT 80.885 186.515 81.055 189.365 ;
        RECT 81.785 188.675 97.785 188.845 ;
        RECT 81.555 187.420 81.725 188.460 ;
        RECT 97.845 187.420 98.015 188.460 ;
        RECT 81.785 187.035 97.785 187.205 ;
        RECT 98.515 186.515 99.045 189.365 ;
        RECT 62.895 186.345 99.045 186.515 ;
        RECT 62.895 183.495 63.425 186.345 ;
        RECT 64.155 185.655 80.155 185.825 ;
        RECT 63.925 184.400 64.095 185.440 ;
        RECT 80.215 184.400 80.385 185.440 ;
        RECT 64.155 184.015 80.155 184.185 ;
        RECT 80.885 183.495 81.055 186.345 ;
        RECT 81.785 185.655 97.785 185.825 ;
        RECT 81.555 184.400 81.725 185.440 ;
        RECT 97.845 184.400 98.015 185.440 ;
        RECT 81.785 184.015 97.785 184.185 ;
        RECT 98.515 183.495 99.045 186.345 ;
        RECT 62.895 183.325 99.045 183.495 ;
        RECT 62.895 180.475 63.425 183.325 ;
        RECT 64.155 182.635 80.155 182.805 ;
        RECT 63.925 181.380 64.095 182.420 ;
        RECT 80.215 181.380 80.385 182.420 ;
        RECT 64.155 180.995 80.155 181.165 ;
        RECT 80.885 180.475 81.055 183.325 ;
        RECT 81.785 182.635 97.785 182.805 ;
        RECT 81.555 181.380 81.725 182.420 ;
        RECT 97.845 181.380 98.015 182.420 ;
        RECT 81.785 180.995 97.785 181.165 ;
        RECT 98.515 180.475 99.045 183.325 ;
        RECT 102.225 181.020 102.625 222.030 ;
        RECT 108.630 220.425 153.130 220.595 ;
        RECT 108.630 216.575 108.800 220.425 ;
        RECT 109.585 219.735 110.585 219.905 ;
        RECT 110.875 219.735 111.875 219.905 ;
        RECT 109.355 217.480 109.525 219.520 ;
        RECT 110.645 217.480 110.815 219.520 ;
        RECT 111.935 217.480 112.105 219.520 ;
        RECT 109.585 217.095 110.585 217.265 ;
        RECT 110.875 217.095 111.875 217.265 ;
        RECT 112.660 216.575 112.830 220.425 ;
        RECT 113.615 219.735 114.615 219.905 ;
        RECT 114.905 219.735 115.905 219.905 ;
        RECT 113.385 217.480 113.555 219.520 ;
        RECT 114.675 217.480 114.845 219.520 ;
        RECT 115.965 217.480 116.135 219.520 ;
        RECT 113.615 217.095 114.615 217.265 ;
        RECT 114.905 217.095 115.905 217.265 ;
        RECT 116.690 216.575 116.860 220.425 ;
        RECT 117.645 219.735 118.645 219.905 ;
        RECT 118.935 219.735 119.935 219.905 ;
        RECT 117.415 217.480 117.585 219.520 ;
        RECT 118.705 217.480 118.875 219.520 ;
        RECT 119.995 217.480 120.165 219.520 ;
        RECT 117.645 217.095 118.645 217.265 ;
        RECT 118.935 217.095 119.935 217.265 ;
        RECT 120.720 216.575 120.890 220.425 ;
        RECT 121.675 219.735 122.675 219.905 ;
        RECT 122.965 219.735 123.965 219.905 ;
        RECT 121.445 217.480 121.615 219.520 ;
        RECT 122.735 217.480 122.905 219.520 ;
        RECT 124.025 217.480 124.195 219.520 ;
        RECT 121.675 217.095 122.675 217.265 ;
        RECT 122.965 217.095 123.965 217.265 ;
        RECT 124.750 216.575 124.920 220.425 ;
        RECT 125.705 219.735 126.705 219.905 ;
        RECT 126.995 219.735 127.995 219.905 ;
        RECT 125.475 217.480 125.645 219.520 ;
        RECT 126.765 217.480 126.935 219.520 ;
        RECT 128.055 217.480 128.225 219.520 ;
        RECT 125.705 217.095 126.705 217.265 ;
        RECT 126.995 217.095 127.995 217.265 ;
        RECT 128.780 216.575 128.950 220.425 ;
        RECT 129.735 219.735 130.735 219.905 ;
        RECT 131.025 219.735 132.025 219.905 ;
        RECT 129.505 217.480 129.675 219.520 ;
        RECT 130.795 217.480 130.965 219.520 ;
        RECT 132.085 217.480 132.255 219.520 ;
        RECT 129.735 217.095 130.735 217.265 ;
        RECT 131.025 217.095 132.025 217.265 ;
        RECT 132.810 216.575 132.980 220.425 ;
        RECT 133.765 219.735 134.765 219.905 ;
        RECT 135.055 219.735 136.055 219.905 ;
        RECT 133.535 217.480 133.705 219.520 ;
        RECT 134.825 217.480 134.995 219.520 ;
        RECT 136.115 217.480 136.285 219.520 ;
        RECT 133.765 217.095 134.765 217.265 ;
        RECT 135.055 217.095 136.055 217.265 ;
        RECT 136.840 216.575 137.010 220.425 ;
        RECT 137.795 219.735 138.795 219.905 ;
        RECT 139.085 219.735 140.085 219.905 ;
        RECT 137.565 217.480 137.735 219.520 ;
        RECT 138.855 217.480 139.025 219.520 ;
        RECT 140.145 217.480 140.315 219.520 ;
        RECT 137.795 217.095 138.795 217.265 ;
        RECT 139.085 217.095 140.085 217.265 ;
        RECT 140.870 216.575 141.040 220.425 ;
        RECT 141.825 219.735 142.825 219.905 ;
        RECT 143.115 219.735 144.115 219.905 ;
        RECT 141.595 217.480 141.765 219.520 ;
        RECT 142.885 217.480 143.055 219.520 ;
        RECT 144.175 217.480 144.345 219.520 ;
        RECT 141.825 217.095 142.825 217.265 ;
        RECT 143.115 217.095 144.115 217.265 ;
        RECT 144.900 216.575 145.070 220.425 ;
        RECT 145.855 219.735 146.855 219.905 ;
        RECT 147.145 219.735 148.145 219.905 ;
        RECT 145.625 217.480 145.795 219.520 ;
        RECT 146.915 217.480 147.085 219.520 ;
        RECT 148.205 217.480 148.375 219.520 ;
        RECT 145.855 217.095 146.855 217.265 ;
        RECT 147.145 217.095 148.145 217.265 ;
        RECT 148.930 216.575 149.100 220.425 ;
        RECT 149.885 219.735 150.885 219.905 ;
        RECT 151.175 219.735 152.175 219.905 ;
        RECT 149.655 217.480 149.825 219.520 ;
        RECT 150.945 217.480 151.115 219.520 ;
        RECT 152.235 217.480 152.405 219.520 ;
        RECT 149.885 217.095 150.885 217.265 ;
        RECT 151.175 217.095 152.175 217.265 ;
        RECT 152.960 216.575 153.130 220.425 ;
        RECT 108.630 216.405 153.130 216.575 ;
        RECT 108.630 213.455 153.130 213.625 ;
        RECT 108.630 203.605 108.800 213.455 ;
        RECT 109.585 212.765 110.585 212.935 ;
        RECT 110.875 212.765 111.875 212.935 ;
        RECT 109.355 204.510 109.525 212.550 ;
        RECT 110.645 204.510 110.815 212.550 ;
        RECT 111.935 204.510 112.105 212.550 ;
        RECT 109.585 204.125 110.585 204.295 ;
        RECT 110.875 204.125 111.875 204.295 ;
        RECT 112.660 203.605 112.830 213.455 ;
        RECT 113.615 212.765 114.615 212.935 ;
        RECT 114.905 212.765 115.905 212.935 ;
        RECT 113.385 204.510 113.555 212.550 ;
        RECT 114.675 204.510 114.845 212.550 ;
        RECT 115.965 204.510 116.135 212.550 ;
        RECT 113.615 204.125 114.615 204.295 ;
        RECT 114.905 204.125 115.905 204.295 ;
        RECT 116.690 203.605 116.860 213.455 ;
        RECT 117.645 212.765 118.645 212.935 ;
        RECT 118.935 212.765 119.935 212.935 ;
        RECT 117.415 204.510 117.585 212.550 ;
        RECT 118.705 204.510 118.875 212.550 ;
        RECT 119.995 204.510 120.165 212.550 ;
        RECT 117.645 204.125 118.645 204.295 ;
        RECT 118.935 204.125 119.935 204.295 ;
        RECT 120.720 203.605 120.890 213.455 ;
        RECT 121.675 212.765 122.675 212.935 ;
        RECT 122.965 212.765 123.965 212.935 ;
        RECT 121.445 204.510 121.615 212.550 ;
        RECT 122.735 204.510 122.905 212.550 ;
        RECT 124.025 204.510 124.195 212.550 ;
        RECT 121.675 204.125 122.675 204.295 ;
        RECT 122.965 204.125 123.965 204.295 ;
        RECT 124.750 203.605 124.920 213.455 ;
        RECT 125.705 212.765 126.705 212.935 ;
        RECT 126.995 212.765 127.995 212.935 ;
        RECT 125.475 204.510 125.645 212.550 ;
        RECT 126.765 204.510 126.935 212.550 ;
        RECT 128.055 204.510 128.225 212.550 ;
        RECT 125.705 204.125 126.705 204.295 ;
        RECT 126.995 204.125 127.995 204.295 ;
        RECT 128.780 203.605 128.950 213.455 ;
        RECT 129.735 212.765 130.735 212.935 ;
        RECT 131.025 212.765 132.025 212.935 ;
        RECT 129.505 204.510 129.675 212.550 ;
        RECT 130.795 204.510 130.965 212.550 ;
        RECT 132.085 204.510 132.255 212.550 ;
        RECT 129.735 204.125 130.735 204.295 ;
        RECT 131.025 204.125 132.025 204.295 ;
        RECT 132.810 203.605 132.980 213.455 ;
        RECT 133.765 212.765 134.765 212.935 ;
        RECT 135.055 212.765 136.055 212.935 ;
        RECT 133.535 204.510 133.705 212.550 ;
        RECT 134.825 204.510 134.995 212.550 ;
        RECT 136.115 204.510 136.285 212.550 ;
        RECT 133.765 204.125 134.765 204.295 ;
        RECT 135.055 204.125 136.055 204.295 ;
        RECT 136.840 203.605 137.010 213.455 ;
        RECT 137.795 212.765 138.795 212.935 ;
        RECT 139.085 212.765 140.085 212.935 ;
        RECT 137.565 204.510 137.735 212.550 ;
        RECT 138.855 204.510 139.025 212.550 ;
        RECT 140.145 204.510 140.315 212.550 ;
        RECT 137.795 204.125 138.795 204.295 ;
        RECT 139.085 204.125 140.085 204.295 ;
        RECT 140.870 203.605 141.040 213.455 ;
        RECT 141.825 212.765 142.825 212.935 ;
        RECT 143.115 212.765 144.115 212.935 ;
        RECT 141.595 204.510 141.765 212.550 ;
        RECT 142.885 204.510 143.055 212.550 ;
        RECT 144.175 204.510 144.345 212.550 ;
        RECT 141.825 204.125 142.825 204.295 ;
        RECT 143.115 204.125 144.115 204.295 ;
        RECT 144.900 203.605 145.070 213.455 ;
        RECT 145.855 212.765 146.855 212.935 ;
        RECT 147.145 212.765 148.145 212.935 ;
        RECT 145.625 204.510 145.795 212.550 ;
        RECT 146.915 204.510 147.085 212.550 ;
        RECT 148.205 204.510 148.375 212.550 ;
        RECT 145.855 204.125 146.855 204.295 ;
        RECT 147.145 204.125 148.145 204.295 ;
        RECT 148.930 203.605 149.100 213.455 ;
        RECT 149.885 212.765 150.885 212.935 ;
        RECT 151.175 212.765 152.175 212.935 ;
        RECT 149.655 204.510 149.825 212.550 ;
        RECT 150.945 204.510 151.115 212.550 ;
        RECT 152.235 204.510 152.405 212.550 ;
        RECT 149.885 204.125 150.885 204.295 ;
        RECT 151.175 204.125 152.175 204.295 ;
        RECT 152.960 203.605 153.130 213.455 ;
        RECT 108.630 203.435 153.130 203.605 ;
        RECT 165.150 201.405 239.210 201.575 ;
        RECT 108.630 200.740 153.130 200.910 ;
        RECT 108.630 194.980 108.800 200.740 ;
        RECT 109.585 200.050 110.585 200.220 ;
        RECT 110.875 200.050 111.875 200.220 ;
        RECT 109.355 195.840 109.525 199.880 ;
        RECT 110.645 195.840 110.815 199.880 ;
        RECT 111.935 195.840 112.105 199.880 ;
        RECT 109.585 195.500 110.585 195.670 ;
        RECT 110.875 195.500 111.875 195.670 ;
        RECT 112.660 194.980 112.830 200.740 ;
        RECT 113.615 200.050 114.615 200.220 ;
        RECT 114.905 200.050 115.905 200.220 ;
        RECT 113.385 195.840 113.555 199.880 ;
        RECT 114.675 195.840 114.845 199.880 ;
        RECT 115.965 195.840 116.135 199.880 ;
        RECT 113.615 195.500 114.615 195.670 ;
        RECT 114.905 195.500 115.905 195.670 ;
        RECT 116.690 194.980 116.860 200.740 ;
        RECT 117.645 200.050 118.645 200.220 ;
        RECT 118.935 200.050 119.935 200.220 ;
        RECT 117.415 195.840 117.585 199.880 ;
        RECT 118.705 195.840 118.875 199.880 ;
        RECT 119.995 195.840 120.165 199.880 ;
        RECT 117.645 195.500 118.645 195.670 ;
        RECT 118.935 195.500 119.935 195.670 ;
        RECT 120.720 194.980 120.890 200.740 ;
        RECT 121.675 200.050 122.675 200.220 ;
        RECT 122.965 200.050 123.965 200.220 ;
        RECT 121.445 195.840 121.615 199.880 ;
        RECT 122.735 195.840 122.905 199.880 ;
        RECT 124.025 195.840 124.195 199.880 ;
        RECT 121.675 195.500 122.675 195.670 ;
        RECT 122.965 195.500 123.965 195.670 ;
        RECT 124.750 194.980 124.920 200.740 ;
        RECT 125.705 200.050 126.705 200.220 ;
        RECT 126.995 200.050 127.995 200.220 ;
        RECT 125.475 195.840 125.645 199.880 ;
        RECT 126.765 195.840 126.935 199.880 ;
        RECT 128.055 195.840 128.225 199.880 ;
        RECT 125.705 195.500 126.705 195.670 ;
        RECT 126.995 195.500 127.995 195.670 ;
        RECT 128.780 194.980 128.950 200.740 ;
        RECT 129.735 200.050 130.735 200.220 ;
        RECT 131.025 200.050 132.025 200.220 ;
        RECT 129.505 195.840 129.675 199.880 ;
        RECT 130.795 195.840 130.965 199.880 ;
        RECT 132.085 195.840 132.255 199.880 ;
        RECT 129.735 195.500 130.735 195.670 ;
        RECT 131.025 195.500 132.025 195.670 ;
        RECT 132.810 194.980 132.980 200.740 ;
        RECT 133.765 200.050 134.765 200.220 ;
        RECT 135.055 200.050 136.055 200.220 ;
        RECT 133.535 195.840 133.705 199.880 ;
        RECT 134.825 195.840 134.995 199.880 ;
        RECT 136.115 195.840 136.285 199.880 ;
        RECT 133.765 195.500 134.765 195.670 ;
        RECT 135.055 195.500 136.055 195.670 ;
        RECT 136.840 194.980 137.010 200.740 ;
        RECT 137.795 200.050 138.795 200.220 ;
        RECT 139.085 200.050 140.085 200.220 ;
        RECT 137.565 195.840 137.735 199.880 ;
        RECT 138.855 195.840 139.025 199.880 ;
        RECT 140.145 195.840 140.315 199.880 ;
        RECT 137.795 195.500 138.795 195.670 ;
        RECT 139.085 195.500 140.085 195.670 ;
        RECT 140.870 194.980 141.040 200.740 ;
        RECT 141.825 200.050 142.825 200.220 ;
        RECT 143.115 200.050 144.115 200.220 ;
        RECT 141.595 195.840 141.765 199.880 ;
        RECT 142.885 195.840 143.055 199.880 ;
        RECT 144.175 195.840 144.345 199.880 ;
        RECT 141.825 195.500 142.825 195.670 ;
        RECT 143.115 195.500 144.115 195.670 ;
        RECT 144.900 194.980 145.070 200.740 ;
        RECT 145.855 200.050 146.855 200.220 ;
        RECT 147.145 200.050 148.145 200.220 ;
        RECT 145.625 195.840 145.795 199.880 ;
        RECT 146.915 195.840 147.085 199.880 ;
        RECT 148.205 195.840 148.375 199.880 ;
        RECT 145.855 195.500 146.855 195.670 ;
        RECT 147.145 195.500 148.145 195.670 ;
        RECT 148.930 194.980 149.100 200.740 ;
        RECT 149.885 200.050 150.885 200.220 ;
        RECT 151.175 200.050 152.175 200.220 ;
        RECT 149.655 195.840 149.825 199.880 ;
        RECT 150.945 195.840 151.115 199.880 ;
        RECT 152.235 195.840 152.405 199.880 ;
        RECT 149.885 195.500 150.885 195.670 ;
        RECT 151.175 195.500 152.175 195.670 ;
        RECT 152.960 194.980 153.130 200.740 ;
        RECT 165.235 200.315 166.445 201.405 ;
        RECT 166.615 200.315 167.825 201.405 ;
        RECT 168.050 200.535 168.335 201.405 ;
        RECT 168.505 200.775 168.765 201.235 ;
        RECT 168.940 200.945 169.195 201.405 ;
        RECT 169.365 200.775 169.625 201.235 ;
        RECT 168.505 200.605 169.625 200.775 ;
        RECT 169.795 200.605 170.105 201.405 ;
        RECT 168.505 200.355 168.765 200.605 ;
        RECT 170.275 200.435 170.585 201.235 ;
        RECT 165.235 199.605 165.755 200.145 ;
        RECT 165.925 199.775 166.445 200.315 ;
        RECT 166.615 199.605 167.135 200.145 ;
        RECT 167.305 199.775 167.825 200.315 ;
        RECT 168.010 200.185 168.765 200.355 ;
        RECT 169.555 200.265 170.585 200.435 ;
        RECT 170.845 200.475 171.015 201.235 ;
        RECT 171.230 200.645 171.560 201.405 ;
        RECT 170.845 200.305 171.560 200.475 ;
        RECT 171.730 200.330 171.985 201.235 ;
        RECT 168.010 199.675 168.415 200.185 ;
        RECT 169.555 200.015 169.725 200.265 ;
        RECT 168.585 199.845 169.725 200.015 ;
        RECT 165.235 198.855 166.445 199.605 ;
        RECT 166.615 198.855 167.825 199.605 ;
        RECT 168.010 199.505 169.660 199.675 ;
        RECT 169.895 199.525 170.245 200.095 ;
        RECT 168.055 198.855 168.335 199.335 ;
        RECT 168.505 199.115 168.765 199.505 ;
        RECT 168.940 198.855 169.195 199.335 ;
        RECT 169.365 199.115 169.660 199.505 ;
        RECT 170.415 199.355 170.585 200.265 ;
        RECT 170.755 199.755 171.110 200.125 ;
        RECT 171.390 200.095 171.560 200.305 ;
        RECT 171.390 199.765 171.645 200.095 ;
        RECT 171.390 199.575 171.560 199.765 ;
        RECT 171.815 199.600 171.985 200.330 ;
        RECT 172.160 200.255 172.420 201.405 ;
        RECT 172.595 200.970 177.940 201.405 ;
        RECT 169.840 198.855 170.115 199.335 ;
        RECT 170.285 199.025 170.585 199.355 ;
        RECT 170.845 199.405 171.560 199.575 ;
        RECT 170.845 199.025 171.015 199.405 ;
        RECT 171.230 198.855 171.560 199.235 ;
        RECT 171.730 199.025 171.985 199.600 ;
        RECT 172.160 198.855 172.420 199.695 ;
        RECT 174.180 199.400 174.520 200.230 ;
        RECT 176.000 199.720 176.350 200.970 ;
        RECT 178.115 200.240 178.405 201.405 ;
        RECT 178.665 200.475 178.835 201.235 ;
        RECT 179.050 200.645 179.380 201.405 ;
        RECT 178.665 200.305 179.380 200.475 ;
        RECT 179.550 200.330 179.805 201.235 ;
        RECT 178.575 199.755 178.930 200.125 ;
        RECT 179.210 200.095 179.380 200.305 ;
        RECT 179.210 199.765 179.465 200.095 ;
        RECT 172.595 198.855 177.940 199.400 ;
        RECT 178.115 198.855 178.405 199.580 ;
        RECT 179.210 199.575 179.380 199.765 ;
        RECT 179.635 199.600 179.805 200.330 ;
        RECT 179.980 200.255 180.240 201.405 ;
        RECT 180.415 200.970 185.760 201.405 ;
        RECT 178.665 199.405 179.380 199.575 ;
        RECT 178.665 199.025 178.835 199.405 ;
        RECT 179.050 198.855 179.380 199.235 ;
        RECT 179.550 199.025 179.805 199.600 ;
        RECT 179.980 198.855 180.240 199.695 ;
        RECT 182.000 199.400 182.340 200.230 ;
        RECT 183.820 199.720 184.170 200.970 ;
        RECT 185.935 200.315 187.605 201.405 ;
        RECT 185.935 199.625 186.685 200.145 ;
        RECT 186.855 199.795 187.605 200.315 ;
        RECT 188.240 200.255 188.500 201.405 ;
        RECT 188.675 200.330 188.930 201.235 ;
        RECT 189.100 200.645 189.430 201.405 ;
        RECT 189.645 200.475 189.815 201.235 ;
        RECT 180.415 198.855 185.760 199.400 ;
        RECT 185.935 198.855 187.605 199.625 ;
        RECT 188.240 198.855 188.500 199.695 ;
        RECT 188.675 199.600 188.845 200.330 ;
        RECT 189.100 200.305 189.815 200.475 ;
        RECT 189.100 200.095 189.270 200.305 ;
        RECT 190.995 200.240 191.285 201.405 ;
        RECT 191.455 200.970 196.800 201.405 ;
        RECT 189.015 199.765 189.270 200.095 ;
        RECT 188.675 199.025 188.930 199.600 ;
        RECT 189.100 199.575 189.270 199.765 ;
        RECT 189.550 199.755 189.905 200.125 ;
        RECT 189.100 199.405 189.815 199.575 ;
        RECT 189.100 198.855 189.430 199.235 ;
        RECT 189.645 199.025 189.815 199.405 ;
        RECT 190.995 198.855 191.285 199.580 ;
        RECT 193.040 199.400 193.380 200.230 ;
        RECT 194.860 199.720 195.210 200.970 ;
        RECT 197.900 200.255 198.160 201.405 ;
        RECT 198.335 200.330 198.590 201.235 ;
        RECT 198.760 200.645 199.090 201.405 ;
        RECT 199.305 200.475 199.475 201.235 ;
        RECT 191.455 198.855 196.800 199.400 ;
        RECT 197.900 198.855 198.160 199.695 ;
        RECT 198.335 199.600 198.505 200.330 ;
        RECT 198.760 200.305 199.475 200.475 ;
        RECT 199.735 200.315 203.245 201.405 ;
        RECT 198.760 200.095 198.930 200.305 ;
        RECT 198.675 199.765 198.930 200.095 ;
        RECT 198.335 199.025 198.590 199.600 ;
        RECT 198.760 199.575 198.930 199.765 ;
        RECT 199.210 199.755 199.565 200.125 ;
        RECT 199.735 199.625 201.385 200.145 ;
        RECT 201.555 199.795 203.245 200.315 ;
        RECT 203.875 200.240 204.165 201.405 ;
        RECT 204.335 200.315 206.925 201.405 ;
        RECT 204.335 199.625 205.545 200.145 ;
        RECT 205.715 199.795 206.925 200.315 ;
        RECT 207.560 200.255 207.820 201.405 ;
        RECT 207.995 200.330 208.250 201.235 ;
        RECT 208.420 200.645 208.750 201.405 ;
        RECT 208.965 200.475 209.135 201.235 ;
        RECT 209.395 200.970 214.740 201.405 ;
        RECT 198.760 199.405 199.475 199.575 ;
        RECT 198.760 198.855 199.090 199.235 ;
        RECT 199.305 199.025 199.475 199.405 ;
        RECT 199.735 198.855 203.245 199.625 ;
        RECT 203.875 198.855 204.165 199.580 ;
        RECT 204.335 198.855 206.925 199.625 ;
        RECT 207.560 198.855 207.820 199.695 ;
        RECT 207.995 199.600 208.165 200.330 ;
        RECT 208.420 200.305 209.135 200.475 ;
        RECT 208.420 200.095 208.590 200.305 ;
        RECT 208.335 199.765 208.590 200.095 ;
        RECT 207.995 199.025 208.250 199.600 ;
        RECT 208.420 199.575 208.590 199.765 ;
        RECT 208.870 199.755 209.225 200.125 ;
        RECT 208.420 199.405 209.135 199.575 ;
        RECT 208.420 198.855 208.750 199.235 ;
        RECT 208.965 199.025 209.135 199.405 ;
        RECT 210.980 199.400 211.320 200.230 ;
        RECT 212.800 199.720 213.150 200.970 ;
        RECT 214.915 200.315 216.585 201.405 ;
        RECT 214.915 199.625 215.665 200.145 ;
        RECT 215.835 199.795 216.585 200.315 ;
        RECT 216.755 200.240 217.045 201.405 ;
        RECT 217.215 200.435 217.525 201.235 ;
        RECT 217.695 200.605 218.005 201.405 ;
        RECT 218.175 200.775 218.435 201.235 ;
        RECT 218.605 200.945 218.860 201.405 ;
        RECT 219.035 200.775 219.295 201.235 ;
        RECT 218.175 200.605 219.295 200.775 ;
        RECT 217.215 200.265 218.245 200.435 ;
        RECT 209.395 198.855 214.740 199.400 ;
        RECT 214.915 198.855 216.585 199.625 ;
        RECT 216.755 198.855 217.045 199.580 ;
        RECT 217.215 199.355 217.385 200.265 ;
        RECT 217.555 199.525 217.905 200.095 ;
        RECT 218.075 200.015 218.245 200.265 ;
        RECT 219.035 200.355 219.295 200.605 ;
        RECT 219.465 200.535 219.750 201.405 ;
        RECT 219.975 200.970 225.320 201.405 ;
        RECT 219.035 200.185 219.790 200.355 ;
        RECT 218.075 199.845 219.215 200.015 ;
        RECT 219.385 199.675 219.790 200.185 ;
        RECT 218.140 199.505 219.790 199.675 ;
        RECT 217.215 199.025 217.515 199.355 ;
        RECT 217.685 198.855 217.960 199.335 ;
        RECT 218.140 199.115 218.435 199.505 ;
        RECT 218.605 198.855 218.860 199.335 ;
        RECT 219.035 199.115 219.295 199.505 ;
        RECT 221.560 199.400 221.900 200.230 ;
        RECT 223.380 199.720 223.730 200.970 ;
        RECT 225.495 200.315 226.705 201.405 ;
        RECT 225.495 199.605 226.015 200.145 ;
        RECT 226.185 199.775 226.705 200.315 ;
        RECT 226.965 200.475 227.135 201.235 ;
        RECT 227.350 200.645 227.680 201.405 ;
        RECT 226.965 200.305 227.680 200.475 ;
        RECT 227.850 200.330 228.105 201.235 ;
        RECT 226.875 199.755 227.230 200.125 ;
        RECT 227.510 200.095 227.680 200.305 ;
        RECT 227.510 199.765 227.765 200.095 ;
        RECT 219.465 198.855 219.745 199.335 ;
        RECT 219.975 198.855 225.320 199.400 ;
        RECT 225.495 198.855 226.705 199.605 ;
        RECT 227.510 199.575 227.680 199.765 ;
        RECT 227.935 199.600 228.105 200.330 ;
        RECT 228.280 200.255 228.540 201.405 ;
        RECT 229.635 200.240 229.925 201.405 ;
        RECT 230.095 200.970 235.440 201.405 ;
        RECT 226.965 199.405 227.680 199.575 ;
        RECT 226.965 199.025 227.135 199.405 ;
        RECT 227.350 198.855 227.680 199.235 ;
        RECT 227.850 199.025 228.105 199.600 ;
        RECT 228.280 198.855 228.540 199.695 ;
        RECT 229.635 198.855 229.925 199.580 ;
        RECT 231.680 199.400 232.020 200.230 ;
        RECT 233.500 199.720 233.850 200.970 ;
        RECT 236.165 200.475 236.335 201.235 ;
        RECT 236.550 200.645 236.880 201.405 ;
        RECT 236.165 200.305 236.880 200.475 ;
        RECT 237.050 200.330 237.305 201.235 ;
        RECT 236.075 199.755 236.430 200.125 ;
        RECT 236.710 200.095 236.880 200.305 ;
        RECT 236.710 199.765 236.965 200.095 ;
        RECT 236.710 199.575 236.880 199.765 ;
        RECT 237.135 199.600 237.305 200.330 ;
        RECT 237.480 200.255 237.740 201.405 ;
        RECT 237.915 200.315 239.125 201.405 ;
        RECT 237.915 199.775 238.435 200.315 ;
        RECT 236.165 199.405 236.880 199.575 ;
        RECT 230.095 198.855 235.440 199.400 ;
        RECT 236.165 199.025 236.335 199.405 ;
        RECT 236.550 198.855 236.880 199.235 ;
        RECT 237.050 199.025 237.305 199.600 ;
        RECT 237.480 198.855 237.740 199.695 ;
        RECT 238.605 199.605 239.125 200.145 ;
        RECT 237.915 198.855 239.125 199.605 ;
        RECT 165.150 198.685 239.210 198.855 ;
        RECT 165.235 197.935 166.445 198.685 ;
        RECT 166.615 198.140 171.960 198.685 ;
        RECT 172.135 198.140 177.480 198.685 ;
        RECT 177.655 198.140 183.000 198.685 ;
        RECT 183.175 198.140 188.520 198.685 ;
        RECT 165.235 197.395 165.755 197.935 ;
        RECT 165.925 197.225 166.445 197.765 ;
        RECT 168.200 197.310 168.540 198.140 ;
        RECT 165.235 196.135 166.445 197.225 ;
        RECT 170.020 196.570 170.370 197.820 ;
        RECT 173.720 197.310 174.060 198.140 ;
        RECT 175.540 196.570 175.890 197.820 ;
        RECT 179.240 197.310 179.580 198.140 ;
        RECT 181.060 196.570 181.410 197.820 ;
        RECT 184.760 197.310 185.100 198.140 ;
        RECT 188.695 197.915 190.365 198.685 ;
        RECT 190.995 197.960 191.285 198.685 ;
        RECT 191.455 198.140 196.800 198.685 ;
        RECT 196.975 198.140 202.320 198.685 ;
        RECT 202.495 198.140 207.840 198.685 ;
        RECT 208.015 198.140 213.360 198.685 ;
        RECT 186.580 196.570 186.930 197.820 ;
        RECT 188.695 197.395 189.445 197.915 ;
        RECT 189.615 197.225 190.365 197.745 ;
        RECT 193.040 197.310 193.380 198.140 ;
        RECT 166.615 196.135 171.960 196.570 ;
        RECT 172.135 196.135 177.480 196.570 ;
        RECT 177.655 196.135 183.000 196.570 ;
        RECT 183.175 196.135 188.520 196.570 ;
        RECT 188.695 196.135 190.365 197.225 ;
        RECT 190.995 196.135 191.285 197.300 ;
        RECT 194.860 196.570 195.210 197.820 ;
        RECT 198.560 197.310 198.900 198.140 ;
        RECT 200.380 196.570 200.730 197.820 ;
        RECT 204.080 197.310 204.420 198.140 ;
        RECT 205.900 196.570 206.250 197.820 ;
        RECT 209.600 197.310 209.940 198.140 ;
        RECT 213.535 197.915 216.125 198.685 ;
        RECT 216.755 197.960 217.045 198.685 ;
        RECT 217.215 198.140 222.560 198.685 ;
        RECT 222.735 198.140 228.080 198.685 ;
        RECT 228.255 198.140 233.600 198.685 ;
        RECT 211.420 196.570 211.770 197.820 ;
        RECT 213.535 197.395 214.745 197.915 ;
        RECT 214.915 197.225 216.125 197.745 ;
        RECT 218.800 197.310 219.140 198.140 ;
        RECT 191.455 196.135 196.800 196.570 ;
        RECT 196.975 196.135 202.320 196.570 ;
        RECT 202.495 196.135 207.840 196.570 ;
        RECT 208.015 196.135 213.360 196.570 ;
        RECT 213.535 196.135 216.125 197.225 ;
        RECT 216.755 196.135 217.045 197.300 ;
        RECT 220.620 196.570 220.970 197.820 ;
        RECT 224.320 197.310 224.660 198.140 ;
        RECT 226.140 196.570 226.490 197.820 ;
        RECT 229.840 197.310 230.180 198.140 ;
        RECT 233.775 197.915 237.285 198.685 ;
        RECT 237.915 197.935 239.125 198.685 ;
        RECT 231.660 196.570 232.010 197.820 ;
        RECT 233.775 197.395 235.425 197.915 ;
        RECT 235.595 197.225 237.285 197.745 ;
        RECT 217.215 196.135 222.560 196.570 ;
        RECT 222.735 196.135 228.080 196.570 ;
        RECT 228.255 196.135 233.600 196.570 ;
        RECT 233.775 196.135 237.285 197.225 ;
        RECT 237.915 197.225 238.435 197.765 ;
        RECT 238.605 197.395 239.125 197.935 ;
        RECT 237.915 196.135 239.125 197.225 ;
        RECT 165.150 195.965 239.210 196.135 ;
        RECT 108.630 194.810 153.130 194.980 ;
        RECT 165.235 194.875 166.445 195.965 ;
        RECT 166.615 195.530 171.960 195.965 ;
        RECT 172.135 195.530 177.480 195.965 ;
        RECT 108.630 185.050 108.800 194.810 ;
        RECT 109.585 194.120 110.585 194.290 ;
        RECT 110.875 194.120 111.875 194.290 ;
        RECT 109.355 185.910 109.525 193.950 ;
        RECT 110.645 185.910 110.815 193.950 ;
        RECT 111.935 185.910 112.105 193.950 ;
        RECT 109.585 185.570 110.585 185.740 ;
        RECT 110.875 185.570 111.875 185.740 ;
        RECT 112.660 185.050 112.830 194.810 ;
        RECT 113.615 194.120 114.615 194.290 ;
        RECT 114.905 194.120 115.905 194.290 ;
        RECT 113.385 185.910 113.555 193.950 ;
        RECT 114.675 185.910 114.845 193.950 ;
        RECT 115.965 185.910 116.135 193.950 ;
        RECT 113.615 185.570 114.615 185.740 ;
        RECT 114.905 185.570 115.905 185.740 ;
        RECT 116.690 185.050 116.860 194.810 ;
        RECT 117.645 194.120 118.645 194.290 ;
        RECT 118.935 194.120 119.935 194.290 ;
        RECT 117.415 185.910 117.585 193.950 ;
        RECT 118.705 185.910 118.875 193.950 ;
        RECT 119.995 185.910 120.165 193.950 ;
        RECT 117.645 185.570 118.645 185.740 ;
        RECT 118.935 185.570 119.935 185.740 ;
        RECT 120.720 185.050 120.890 194.810 ;
        RECT 121.675 194.120 122.675 194.290 ;
        RECT 122.965 194.120 123.965 194.290 ;
        RECT 121.445 185.910 121.615 193.950 ;
        RECT 122.735 185.910 122.905 193.950 ;
        RECT 124.025 185.910 124.195 193.950 ;
        RECT 121.675 185.570 122.675 185.740 ;
        RECT 122.965 185.570 123.965 185.740 ;
        RECT 124.750 185.050 124.920 194.810 ;
        RECT 125.705 194.120 126.705 194.290 ;
        RECT 126.995 194.120 127.995 194.290 ;
        RECT 125.475 185.910 125.645 193.950 ;
        RECT 126.765 185.910 126.935 193.950 ;
        RECT 128.055 185.910 128.225 193.950 ;
        RECT 125.705 185.570 126.705 185.740 ;
        RECT 126.995 185.570 127.995 185.740 ;
        RECT 128.780 185.050 128.950 194.810 ;
        RECT 129.735 194.120 130.735 194.290 ;
        RECT 131.025 194.120 132.025 194.290 ;
        RECT 129.505 185.910 129.675 193.950 ;
        RECT 130.795 185.910 130.965 193.950 ;
        RECT 132.085 185.910 132.255 193.950 ;
        RECT 129.735 185.570 130.735 185.740 ;
        RECT 131.025 185.570 132.025 185.740 ;
        RECT 132.810 185.050 132.980 194.810 ;
        RECT 133.765 194.120 134.765 194.290 ;
        RECT 135.055 194.120 136.055 194.290 ;
        RECT 133.535 185.910 133.705 193.950 ;
        RECT 134.825 185.910 134.995 193.950 ;
        RECT 136.115 185.910 136.285 193.950 ;
        RECT 133.765 185.570 134.765 185.740 ;
        RECT 135.055 185.570 136.055 185.740 ;
        RECT 136.840 185.050 137.010 194.810 ;
        RECT 137.795 194.120 138.795 194.290 ;
        RECT 139.085 194.120 140.085 194.290 ;
        RECT 137.565 185.910 137.735 193.950 ;
        RECT 138.855 185.910 139.025 193.950 ;
        RECT 140.145 185.910 140.315 193.950 ;
        RECT 137.795 185.570 138.795 185.740 ;
        RECT 139.085 185.570 140.085 185.740 ;
        RECT 140.870 185.050 141.040 194.810 ;
        RECT 141.825 194.120 142.825 194.290 ;
        RECT 143.115 194.120 144.115 194.290 ;
        RECT 141.595 185.910 141.765 193.950 ;
        RECT 142.885 185.910 143.055 193.950 ;
        RECT 144.175 185.910 144.345 193.950 ;
        RECT 141.825 185.570 142.825 185.740 ;
        RECT 143.115 185.570 144.115 185.740 ;
        RECT 144.900 185.050 145.070 194.810 ;
        RECT 145.855 194.120 146.855 194.290 ;
        RECT 147.145 194.120 148.145 194.290 ;
        RECT 145.625 185.910 145.795 193.950 ;
        RECT 146.915 185.910 147.085 193.950 ;
        RECT 148.205 185.910 148.375 193.950 ;
        RECT 145.855 185.570 146.855 185.740 ;
        RECT 147.145 185.570 148.145 185.740 ;
        RECT 148.930 185.050 149.100 194.810 ;
        RECT 149.885 194.120 150.885 194.290 ;
        RECT 151.175 194.120 152.175 194.290 ;
        RECT 149.655 185.910 149.825 193.950 ;
        RECT 150.945 185.910 151.115 193.950 ;
        RECT 152.235 185.910 152.405 193.950 ;
        RECT 149.885 185.570 150.885 185.740 ;
        RECT 151.175 185.570 152.175 185.740 ;
        RECT 152.960 185.050 153.130 194.810 ;
        RECT 165.235 194.165 165.755 194.705 ;
        RECT 165.925 194.335 166.445 194.875 ;
        RECT 165.235 193.415 166.445 194.165 ;
        RECT 168.200 193.960 168.540 194.790 ;
        RECT 170.020 194.280 170.370 195.530 ;
        RECT 173.720 193.960 174.060 194.790 ;
        RECT 175.540 194.280 175.890 195.530 ;
        RECT 178.115 194.800 178.405 195.965 ;
        RECT 178.575 195.530 183.920 195.965 ;
        RECT 166.615 193.415 171.960 193.960 ;
        RECT 172.135 193.415 177.480 193.960 ;
        RECT 178.115 193.415 178.405 194.140 ;
        RECT 180.160 193.960 180.500 194.790 ;
        RECT 181.980 194.280 182.330 195.530 ;
        RECT 184.095 194.875 187.605 195.965 ;
        RECT 187.775 194.875 188.985 195.965 ;
        RECT 184.095 194.185 185.745 194.705 ;
        RECT 185.915 194.355 187.605 194.875 ;
        RECT 178.575 193.415 183.920 193.960 ;
        RECT 184.095 193.415 187.605 194.185 ;
        RECT 187.775 194.165 188.295 194.705 ;
        RECT 188.465 194.335 188.985 194.875 ;
        RECT 189.155 194.360 189.435 195.795 ;
        RECT 189.605 195.190 190.315 195.965 ;
        RECT 190.485 195.020 190.815 195.795 ;
        RECT 189.665 194.805 190.815 195.020 ;
        RECT 187.775 193.415 188.985 194.165 ;
        RECT 189.155 193.585 189.495 194.360 ;
        RECT 189.665 194.235 189.950 194.805 ;
        RECT 190.135 194.405 190.605 194.635 ;
        RECT 191.010 194.605 191.225 195.720 ;
        RECT 191.405 195.245 191.735 195.965 ;
        RECT 191.515 194.605 191.745 194.945 ;
        RECT 191.915 194.875 195.425 195.965 ;
        RECT 190.775 194.425 191.225 194.605 ;
        RECT 190.775 194.405 191.105 194.425 ;
        RECT 191.415 194.405 191.745 194.605 ;
        RECT 189.665 194.045 190.375 194.235 ;
        RECT 190.075 193.905 190.375 194.045 ;
        RECT 190.565 194.045 191.745 194.235 ;
        RECT 190.565 193.965 190.895 194.045 ;
        RECT 190.075 193.895 190.390 193.905 ;
        RECT 190.075 193.885 190.400 193.895 ;
        RECT 190.075 193.880 190.410 193.885 ;
        RECT 189.665 193.415 189.835 193.875 ;
        RECT 190.075 193.870 190.415 193.880 ;
        RECT 190.075 193.865 190.420 193.870 ;
        RECT 190.075 193.855 190.425 193.865 ;
        RECT 190.075 193.850 190.430 193.855 ;
        RECT 190.075 193.585 190.435 193.850 ;
        RECT 191.065 193.415 191.235 193.875 ;
        RECT 191.405 193.585 191.745 194.045 ;
        RECT 191.915 194.185 193.565 194.705 ;
        RECT 193.735 194.355 195.425 194.875 ;
        RECT 195.635 194.825 195.865 195.965 ;
        RECT 196.035 194.815 196.365 195.795 ;
        RECT 196.535 194.825 196.745 195.965 ;
        RECT 196.975 195.530 202.320 195.965 ;
        RECT 195.615 194.405 195.945 194.655 ;
        RECT 191.915 193.415 195.425 194.185 ;
        RECT 195.635 193.415 195.865 194.235 ;
        RECT 196.115 194.215 196.365 194.815 ;
        RECT 196.035 193.585 196.365 194.215 ;
        RECT 196.535 193.415 196.745 194.235 ;
        RECT 198.560 193.960 198.900 194.790 ;
        RECT 200.380 194.280 200.730 195.530 ;
        RECT 202.495 194.875 203.705 195.965 ;
        RECT 202.495 194.165 203.015 194.705 ;
        RECT 203.185 194.335 203.705 194.875 ;
        RECT 203.875 194.800 204.165 195.965 ;
        RECT 204.335 195.530 209.680 195.965 ;
        RECT 209.855 195.530 215.200 195.965 ;
        RECT 215.375 195.530 220.720 195.965 ;
        RECT 220.895 195.530 226.240 195.965 ;
        RECT 196.975 193.415 202.320 193.960 ;
        RECT 202.495 193.415 203.705 194.165 ;
        RECT 203.875 193.415 204.165 194.140 ;
        RECT 205.920 193.960 206.260 194.790 ;
        RECT 207.740 194.280 208.090 195.530 ;
        RECT 211.440 193.960 211.780 194.790 ;
        RECT 213.260 194.280 213.610 195.530 ;
        RECT 216.960 193.960 217.300 194.790 ;
        RECT 218.780 194.280 219.130 195.530 ;
        RECT 222.480 193.960 222.820 194.790 ;
        RECT 224.300 194.280 224.650 195.530 ;
        RECT 226.415 194.875 229.005 195.965 ;
        RECT 226.415 194.185 227.625 194.705 ;
        RECT 227.795 194.355 229.005 194.875 ;
        RECT 229.635 194.800 229.925 195.965 ;
        RECT 230.095 195.530 235.440 195.965 ;
        RECT 204.335 193.415 209.680 193.960 ;
        RECT 209.855 193.415 215.200 193.960 ;
        RECT 215.375 193.415 220.720 193.960 ;
        RECT 220.895 193.415 226.240 193.960 ;
        RECT 226.415 193.415 229.005 194.185 ;
        RECT 229.635 193.415 229.925 194.140 ;
        RECT 231.680 193.960 232.020 194.790 ;
        RECT 233.500 194.280 233.850 195.530 ;
        RECT 235.615 194.875 237.285 195.965 ;
        RECT 235.615 194.185 236.365 194.705 ;
        RECT 236.535 194.355 237.285 194.875 ;
        RECT 237.915 194.875 239.125 195.965 ;
        RECT 237.915 194.335 238.435 194.875 ;
        RECT 230.095 193.415 235.440 193.960 ;
        RECT 235.615 193.415 237.285 194.185 ;
        RECT 238.605 194.165 239.125 194.705 ;
        RECT 237.915 193.415 239.125 194.165 ;
        RECT 165.150 193.245 239.210 193.415 ;
        RECT 165.235 192.495 166.445 193.245 ;
        RECT 166.615 192.700 171.960 193.245 ;
        RECT 165.235 191.955 165.755 192.495 ;
        RECT 165.925 191.785 166.445 192.325 ;
        RECT 168.200 191.870 168.540 192.700 ;
        RECT 172.135 192.475 173.805 193.245 ;
        RECT 174.435 192.570 174.695 193.075 ;
        RECT 174.875 192.865 175.205 193.245 ;
        RECT 175.385 192.695 175.555 193.075 ;
        RECT 165.235 190.695 166.445 191.785 ;
        RECT 170.020 191.130 170.370 192.380 ;
        RECT 172.135 191.955 172.885 192.475 ;
        RECT 173.055 191.785 173.805 192.305 ;
        RECT 166.615 190.695 171.960 191.130 ;
        RECT 172.135 190.695 173.805 191.785 ;
        RECT 174.435 191.770 174.605 192.570 ;
        RECT 174.890 192.525 175.555 192.695 ;
        RECT 176.275 192.570 176.535 193.075 ;
        RECT 176.715 192.865 177.045 193.245 ;
        RECT 177.225 192.695 177.395 193.075 ;
        RECT 174.890 192.270 175.060 192.525 ;
        RECT 174.775 191.940 175.060 192.270 ;
        RECT 175.295 191.975 175.625 192.345 ;
        RECT 174.890 191.795 175.060 191.940 ;
        RECT 174.435 190.865 174.705 191.770 ;
        RECT 174.890 191.625 175.555 191.795 ;
        RECT 174.875 190.695 175.205 191.455 ;
        RECT 175.385 190.865 175.555 191.625 ;
        RECT 176.275 191.770 176.445 192.570 ;
        RECT 176.730 192.525 177.395 192.695 ;
        RECT 176.730 192.270 176.900 192.525 ;
        RECT 176.615 191.940 176.900 192.270 ;
        RECT 177.135 191.975 177.465 192.345 ;
        RECT 178.115 192.300 178.455 193.075 ;
        RECT 178.625 192.785 178.795 193.245 ;
        RECT 179.035 192.810 179.395 193.075 ;
        RECT 179.035 192.805 179.390 192.810 ;
        RECT 179.035 192.795 179.385 192.805 ;
        RECT 179.035 192.790 179.380 192.795 ;
        RECT 179.035 192.780 179.375 192.790 ;
        RECT 180.025 192.785 180.195 193.245 ;
        RECT 179.035 192.775 179.370 192.780 ;
        RECT 179.035 192.765 179.360 192.775 ;
        RECT 179.035 192.755 179.350 192.765 ;
        RECT 179.035 192.615 179.335 192.755 ;
        RECT 178.625 192.425 179.335 192.615 ;
        RECT 179.525 192.615 179.855 192.695 ;
        RECT 180.365 192.615 180.705 193.075 ;
        RECT 179.525 192.425 180.705 192.615 ;
        RECT 180.900 192.595 181.210 193.065 ;
        RECT 181.380 192.765 182.115 193.245 ;
        RECT 182.285 192.675 182.455 193.025 ;
        RECT 182.625 192.845 183.005 193.245 ;
        RECT 180.900 192.425 181.635 192.595 ;
        RECT 182.285 192.505 183.025 192.675 ;
        RECT 183.195 192.570 183.465 192.915 ;
        RECT 176.730 191.795 176.900 191.940 ;
        RECT 176.275 190.865 176.545 191.770 ;
        RECT 176.730 191.625 177.395 191.795 ;
        RECT 176.715 190.695 177.045 191.455 ;
        RECT 177.225 190.865 177.395 191.625 ;
        RECT 178.115 190.865 178.395 192.300 ;
        RECT 178.625 191.855 178.910 192.425 ;
        RECT 181.385 192.335 181.635 192.425 ;
        RECT 182.855 192.335 183.025 192.505 ;
        RECT 179.095 192.025 179.565 192.255 ;
        RECT 179.735 192.235 180.065 192.255 ;
        RECT 179.735 192.055 180.185 192.235 ;
        RECT 180.375 192.055 180.705 192.255 ;
        RECT 178.625 191.640 179.775 191.855 ;
        RECT 178.565 190.695 179.275 191.470 ;
        RECT 179.445 190.865 179.775 191.640 ;
        RECT 179.970 190.940 180.185 192.055 ;
        RECT 180.475 191.715 180.705 192.055 ;
        RECT 180.880 192.005 181.215 192.255 ;
        RECT 181.385 192.005 182.125 192.335 ;
        RECT 182.855 192.005 183.085 192.335 ;
        RECT 180.365 190.695 180.695 191.415 ;
        RECT 180.880 190.695 181.135 191.835 ;
        RECT 181.385 191.445 181.555 192.005 ;
        RECT 182.855 191.835 183.025 192.005 ;
        RECT 183.295 191.885 183.465 192.570 ;
        RECT 183.725 192.595 183.895 193.075 ;
        RECT 184.065 192.765 184.395 193.245 ;
        RECT 184.620 192.825 186.155 193.075 ;
        RECT 184.620 192.595 184.790 192.825 ;
        RECT 183.725 192.425 184.790 192.595 ;
        RECT 184.970 192.255 185.250 192.655 ;
        RECT 183.640 192.045 183.990 192.255 ;
        RECT 184.160 192.055 184.605 192.255 ;
        RECT 184.775 192.055 185.250 192.255 ;
        RECT 185.520 192.255 185.805 192.655 ;
        RECT 185.985 192.595 186.155 192.825 ;
        RECT 186.325 192.765 186.655 193.245 ;
        RECT 186.870 192.745 187.125 193.075 ;
        RECT 186.915 192.735 187.125 192.745 ;
        RECT 186.940 192.665 187.125 192.735 ;
        RECT 185.985 192.425 186.785 192.595 ;
        RECT 185.520 192.055 185.850 192.255 ;
        RECT 186.020 192.055 186.385 192.255 ;
        RECT 183.235 191.835 183.465 191.885 ;
        RECT 186.615 191.875 186.785 192.425 ;
        RECT 181.780 191.665 183.025 191.835 ;
        RECT 181.780 191.415 182.200 191.665 ;
        RECT 181.330 190.915 182.525 191.245 ;
        RECT 182.705 190.695 182.985 191.495 ;
        RECT 183.195 190.865 183.465 191.835 ;
        RECT 183.725 191.705 186.785 191.875 ;
        RECT 183.725 190.865 183.895 191.705 ;
        RECT 186.955 191.535 187.125 192.665 ;
        RECT 188.260 192.595 188.570 193.065 ;
        RECT 188.740 192.765 189.475 193.245 ;
        RECT 189.645 192.675 189.815 193.025 ;
        RECT 189.985 192.845 190.365 193.245 ;
        RECT 188.260 192.425 188.995 192.595 ;
        RECT 189.645 192.505 190.385 192.675 ;
        RECT 190.555 192.570 190.825 192.915 ;
        RECT 188.745 192.335 188.995 192.425 ;
        RECT 190.215 192.335 190.385 192.505 ;
        RECT 188.240 192.005 188.575 192.255 ;
        RECT 188.745 192.005 189.485 192.335 ;
        RECT 190.215 192.005 190.445 192.335 ;
        RECT 184.065 191.035 184.395 191.535 ;
        RECT 184.565 191.295 186.200 191.535 ;
        RECT 184.565 191.205 184.795 191.295 ;
        RECT 184.905 191.035 185.235 191.075 ;
        RECT 184.065 190.865 185.235 191.035 ;
        RECT 185.425 190.695 185.780 191.115 ;
        RECT 185.950 190.865 186.200 191.295 ;
        RECT 186.370 190.695 186.700 191.455 ;
        RECT 186.870 190.865 187.125 191.535 ;
        RECT 188.240 190.695 188.495 191.835 ;
        RECT 188.745 191.445 188.915 192.005 ;
        RECT 190.215 191.835 190.385 192.005 ;
        RECT 190.655 191.885 190.825 192.570 ;
        RECT 190.995 192.520 191.285 193.245 ;
        RECT 192.465 192.595 192.635 193.075 ;
        RECT 192.805 192.765 193.135 193.245 ;
        RECT 193.360 192.825 194.895 193.075 ;
        RECT 193.360 192.595 193.530 192.825 ;
        RECT 192.465 192.425 193.530 192.595 ;
        RECT 193.710 192.255 193.990 192.655 ;
        RECT 192.380 192.045 192.730 192.255 ;
        RECT 192.900 192.055 193.345 192.255 ;
        RECT 193.515 192.055 193.990 192.255 ;
        RECT 194.260 192.255 194.545 192.655 ;
        RECT 194.725 192.595 194.895 192.825 ;
        RECT 195.065 192.765 195.395 193.245 ;
        RECT 195.610 192.745 195.865 193.075 ;
        RECT 195.680 192.665 195.865 192.745 ;
        RECT 194.725 192.425 195.525 192.595 ;
        RECT 194.260 192.055 194.590 192.255 ;
        RECT 194.760 192.055 195.125 192.255 ;
        RECT 190.595 191.835 190.825 191.885 ;
        RECT 195.355 191.875 195.525 192.425 ;
        RECT 189.140 191.665 190.385 191.835 ;
        RECT 189.140 191.415 189.560 191.665 ;
        RECT 188.690 190.915 189.885 191.245 ;
        RECT 190.065 190.695 190.345 191.495 ;
        RECT 190.555 190.865 190.825 191.835 ;
        RECT 190.995 190.695 191.285 191.860 ;
        RECT 192.465 191.705 195.525 191.875 ;
        RECT 192.465 190.865 192.635 191.705 ;
        RECT 195.695 191.545 195.865 192.665 ;
        RECT 196.055 192.475 198.645 193.245 ;
        RECT 196.055 191.955 197.265 192.475 ;
        RECT 197.435 191.785 198.645 192.305 ;
        RECT 195.655 191.535 195.865 191.545 ;
        RECT 192.805 191.035 193.135 191.535 ;
        RECT 193.305 191.295 194.940 191.535 ;
        RECT 193.305 191.205 193.535 191.295 ;
        RECT 193.645 191.035 193.975 191.075 ;
        RECT 192.805 190.865 193.975 191.035 ;
        RECT 194.165 190.695 194.520 191.115 ;
        RECT 194.690 190.865 194.940 191.295 ;
        RECT 195.110 190.695 195.440 191.455 ;
        RECT 195.610 190.865 195.865 191.535 ;
        RECT 196.055 190.695 198.645 191.785 ;
        RECT 199.275 192.300 199.615 193.075 ;
        RECT 199.785 192.785 199.955 193.245 ;
        RECT 200.195 192.810 200.555 193.075 ;
        RECT 200.195 192.805 200.550 192.810 ;
        RECT 200.195 192.795 200.545 192.805 ;
        RECT 200.195 192.790 200.540 192.795 ;
        RECT 200.195 192.780 200.535 192.790 ;
        RECT 201.185 192.785 201.355 193.245 ;
        RECT 200.195 192.775 200.530 192.780 ;
        RECT 200.195 192.765 200.520 192.775 ;
        RECT 200.195 192.755 200.510 192.765 ;
        RECT 200.195 192.615 200.495 192.755 ;
        RECT 199.785 192.425 200.495 192.615 ;
        RECT 200.685 192.615 201.015 192.695 ;
        RECT 201.525 192.615 201.865 193.075 ;
        RECT 202.035 192.700 207.380 193.245 ;
        RECT 207.555 192.700 212.900 193.245 ;
        RECT 200.685 192.425 201.865 192.615 ;
        RECT 199.275 190.865 199.555 192.300 ;
        RECT 199.785 191.855 200.070 192.425 ;
        RECT 200.255 192.025 200.725 192.255 ;
        RECT 200.895 192.235 201.225 192.255 ;
        RECT 200.895 192.055 201.345 192.235 ;
        RECT 201.535 192.055 201.865 192.255 ;
        RECT 199.785 191.640 200.935 191.855 ;
        RECT 199.725 190.695 200.435 191.470 ;
        RECT 200.605 190.865 200.935 191.640 ;
        RECT 201.130 190.940 201.345 192.055 ;
        RECT 201.635 191.715 201.865 192.055 ;
        RECT 203.620 191.870 203.960 192.700 ;
        RECT 201.525 190.695 201.855 191.415 ;
        RECT 205.440 191.130 205.790 192.380 ;
        RECT 209.140 191.870 209.480 192.700 ;
        RECT 213.075 192.475 216.585 193.245 ;
        RECT 216.755 192.520 217.045 193.245 ;
        RECT 217.215 192.700 222.560 193.245 ;
        RECT 222.735 192.700 228.080 193.245 ;
        RECT 228.255 192.700 233.600 193.245 ;
        RECT 210.960 191.130 211.310 192.380 ;
        RECT 213.075 191.955 214.725 192.475 ;
        RECT 214.895 191.785 216.585 192.305 ;
        RECT 218.800 191.870 219.140 192.700 ;
        RECT 202.035 190.695 207.380 191.130 ;
        RECT 207.555 190.695 212.900 191.130 ;
        RECT 213.075 190.695 216.585 191.785 ;
        RECT 216.755 190.695 217.045 191.860 ;
        RECT 220.620 191.130 220.970 192.380 ;
        RECT 224.320 191.870 224.660 192.700 ;
        RECT 226.140 191.130 226.490 192.380 ;
        RECT 229.840 191.870 230.180 192.700 ;
        RECT 233.775 192.475 237.285 193.245 ;
        RECT 237.915 192.495 239.125 193.245 ;
        RECT 231.660 191.130 232.010 192.380 ;
        RECT 233.775 191.955 235.425 192.475 ;
        RECT 235.595 191.785 237.285 192.305 ;
        RECT 217.215 190.695 222.560 191.130 ;
        RECT 222.735 190.695 228.080 191.130 ;
        RECT 228.255 190.695 233.600 191.130 ;
        RECT 233.775 190.695 237.285 191.785 ;
        RECT 237.915 191.785 238.435 192.325 ;
        RECT 238.605 191.955 239.125 192.495 ;
        RECT 237.915 190.695 239.125 191.785 ;
        RECT 165.150 190.525 239.210 190.695 ;
        RECT 165.235 189.435 166.445 190.525 ;
        RECT 165.235 188.725 165.755 189.265 ;
        RECT 165.925 188.895 166.445 189.435 ;
        RECT 166.695 189.595 166.875 190.355 ;
        RECT 167.055 189.765 167.385 190.525 ;
        RECT 166.695 189.425 167.370 189.595 ;
        RECT 167.555 189.450 167.825 190.355 ;
        RECT 167.200 189.280 167.370 189.425 ;
        RECT 166.635 188.875 166.975 189.245 ;
        RECT 167.200 188.950 167.475 189.280 ;
        RECT 165.235 187.975 166.445 188.725 ;
        RECT 167.200 188.695 167.370 188.950 ;
        RECT 166.705 188.525 167.370 188.695 ;
        RECT 167.645 188.650 167.825 189.450 ;
        RECT 167.995 189.435 171.505 190.525 ;
        RECT 166.705 188.145 166.875 188.525 ;
        RECT 167.055 187.975 167.385 188.355 ;
        RECT 167.565 188.145 167.825 188.650 ;
        RECT 167.995 188.745 169.645 189.265 ;
        RECT 169.815 188.915 171.505 189.435 ;
        RECT 171.765 189.595 171.935 190.355 ;
        RECT 172.115 189.765 172.445 190.525 ;
        RECT 171.765 189.425 172.430 189.595 ;
        RECT 172.615 189.450 172.885 190.355 ;
        RECT 172.260 189.280 172.430 189.425 ;
        RECT 171.695 188.875 172.025 189.245 ;
        RECT 172.260 188.950 172.545 189.280 ;
        RECT 167.995 187.975 171.505 188.745 ;
        RECT 172.260 188.695 172.430 188.950 ;
        RECT 171.765 188.525 172.430 188.695 ;
        RECT 172.715 188.650 172.885 189.450 ;
        RECT 173.270 189.425 173.600 190.525 ;
        RECT 174.075 189.925 174.400 190.355 ;
        RECT 174.570 190.105 174.900 190.525 ;
        RECT 175.645 190.095 176.055 190.525 ;
        RECT 174.075 189.755 176.055 189.925 ;
        RECT 174.075 189.345 174.780 189.755 ;
        RECT 173.055 188.965 173.700 189.175 ;
        RECT 173.870 188.965 174.440 189.175 ;
        RECT 171.765 188.145 171.935 188.525 ;
        RECT 172.115 187.975 172.445 188.355 ;
        RECT 172.625 188.145 172.885 188.650 ;
        RECT 173.210 188.625 174.380 188.795 ;
        RECT 173.210 188.160 173.540 188.625 ;
        RECT 173.710 187.975 173.880 188.445 ;
        RECT 174.050 188.145 174.380 188.625 ;
        RECT 174.610 188.145 174.780 189.345 ;
        RECT 174.950 189.415 175.575 189.585 ;
        RECT 174.950 188.715 175.120 189.415 ;
        RECT 175.790 189.215 176.055 189.755 ;
        RECT 176.225 189.370 176.565 190.355 ;
        RECT 176.825 189.595 176.995 190.355 ;
        RECT 177.175 189.765 177.505 190.525 ;
        RECT 176.825 189.425 177.490 189.595 ;
        RECT 177.675 189.450 177.945 190.355 ;
        RECT 175.290 188.885 175.620 189.215 ;
        RECT 175.790 188.885 176.140 189.215 ;
        RECT 176.310 188.715 176.565 189.370 ;
        RECT 177.320 189.280 177.490 189.425 ;
        RECT 176.755 188.875 177.085 189.245 ;
        RECT 177.320 188.950 177.605 189.280 ;
        RECT 174.950 188.545 175.490 188.715 ;
        RECT 175.320 188.340 175.490 188.545 ;
        RECT 175.770 187.975 175.940 188.715 ;
        RECT 176.205 188.340 176.565 188.715 ;
        RECT 177.320 188.695 177.490 188.950 ;
        RECT 176.825 188.525 177.490 188.695 ;
        RECT 177.775 188.650 177.945 189.450 ;
        RECT 178.115 189.360 178.405 190.525 ;
        RECT 178.575 188.920 178.855 190.355 ;
        RECT 179.025 189.750 179.735 190.525 ;
        RECT 179.905 189.580 180.235 190.355 ;
        RECT 179.085 189.365 180.235 189.580 ;
        RECT 176.335 188.315 176.505 188.340 ;
        RECT 176.825 188.145 176.995 188.525 ;
        RECT 177.175 187.975 177.505 188.355 ;
        RECT 177.685 188.145 177.945 188.650 ;
        RECT 178.115 187.975 178.405 188.700 ;
        RECT 178.575 188.145 178.915 188.920 ;
        RECT 179.085 188.795 179.370 189.365 ;
        RECT 179.555 188.965 180.025 189.195 ;
        RECT 180.430 189.165 180.645 190.280 ;
        RECT 180.825 189.805 181.155 190.525 ;
        RECT 180.935 189.165 181.165 189.505 ;
        RECT 180.195 188.985 180.645 189.165 ;
        RECT 180.195 188.965 180.525 188.985 ;
        RECT 180.835 188.965 181.165 189.165 ;
        RECT 181.795 189.450 182.065 190.355 ;
        RECT 182.235 189.765 182.565 190.525 ;
        RECT 182.745 189.595 182.915 190.355 ;
        RECT 179.085 188.605 179.795 188.795 ;
        RECT 179.495 188.465 179.795 188.605 ;
        RECT 179.985 188.605 181.165 188.795 ;
        RECT 179.985 188.525 180.315 188.605 ;
        RECT 179.495 188.455 179.810 188.465 ;
        RECT 179.495 188.445 179.820 188.455 ;
        RECT 179.495 188.440 179.830 188.445 ;
        RECT 179.085 187.975 179.255 188.435 ;
        RECT 179.495 188.430 179.835 188.440 ;
        RECT 179.495 188.425 179.840 188.430 ;
        RECT 179.495 188.415 179.845 188.425 ;
        RECT 179.495 188.410 179.850 188.415 ;
        RECT 179.495 188.145 179.855 188.410 ;
        RECT 180.485 187.975 180.655 188.435 ;
        RECT 180.825 188.145 181.165 188.605 ;
        RECT 181.795 188.650 181.965 189.450 ;
        RECT 182.250 189.425 182.915 189.595 ;
        RECT 183.725 189.595 183.895 190.355 ;
        RECT 184.075 189.765 184.405 190.525 ;
        RECT 183.725 189.425 184.390 189.595 ;
        RECT 184.575 189.450 184.845 190.355 ;
        RECT 182.250 189.280 182.420 189.425 ;
        RECT 182.135 188.950 182.420 189.280 ;
        RECT 184.220 189.280 184.390 189.425 ;
        RECT 182.250 188.695 182.420 188.950 ;
        RECT 182.655 188.875 182.985 189.245 ;
        RECT 183.655 188.875 183.985 189.245 ;
        RECT 184.220 188.950 184.505 189.280 ;
        RECT 184.220 188.695 184.390 188.950 ;
        RECT 181.795 188.145 182.055 188.650 ;
        RECT 182.250 188.525 182.915 188.695 ;
        RECT 182.235 187.975 182.565 188.355 ;
        RECT 182.745 188.145 182.915 188.525 ;
        RECT 183.725 188.525 184.390 188.695 ;
        RECT 184.675 188.650 184.845 189.450 ;
        RECT 185.565 189.595 185.735 190.355 ;
        RECT 185.915 189.765 186.245 190.525 ;
        RECT 185.565 189.425 186.230 189.595 ;
        RECT 186.415 189.450 186.685 190.355 ;
        RECT 186.060 189.280 186.230 189.425 ;
        RECT 185.495 188.875 185.825 189.245 ;
        RECT 186.060 188.950 186.345 189.280 ;
        RECT 186.060 188.695 186.230 188.950 ;
        RECT 183.725 188.145 183.895 188.525 ;
        RECT 184.075 187.975 184.405 188.355 ;
        RECT 184.585 188.145 184.845 188.650 ;
        RECT 185.565 188.525 186.230 188.695 ;
        RECT 186.515 188.650 186.685 189.450 ;
        RECT 187.405 189.595 187.575 190.355 ;
        RECT 187.755 189.765 188.085 190.525 ;
        RECT 187.405 189.425 188.070 189.595 ;
        RECT 188.255 189.450 188.525 190.355 ;
        RECT 187.900 189.280 188.070 189.425 ;
        RECT 187.335 188.875 187.665 189.245 ;
        RECT 187.900 188.950 188.185 189.280 ;
        RECT 187.900 188.695 188.070 188.950 ;
        RECT 185.565 188.145 185.735 188.525 ;
        RECT 185.915 187.975 186.245 188.355 ;
        RECT 186.425 188.145 186.685 188.650 ;
        RECT 187.405 188.525 188.070 188.695 ;
        RECT 188.355 188.650 188.525 189.450 ;
        RECT 187.405 188.145 187.575 188.525 ;
        RECT 187.755 187.975 188.085 188.355 ;
        RECT 188.265 188.145 188.525 188.650 ;
        RECT 188.695 189.450 188.965 190.355 ;
        RECT 189.135 189.765 189.465 190.525 ;
        RECT 189.645 189.595 189.815 190.355 ;
        RECT 188.695 188.650 188.865 189.450 ;
        RECT 189.150 189.425 189.815 189.595 ;
        RECT 189.150 189.280 189.320 189.425 ;
        RECT 190.080 189.385 190.335 190.525 ;
        RECT 190.530 189.975 191.725 190.305 ;
        RECT 189.035 188.950 189.320 189.280 ;
        RECT 189.150 188.695 189.320 188.950 ;
        RECT 189.555 188.875 189.885 189.245 ;
        RECT 190.585 189.215 190.755 189.775 ;
        RECT 190.980 189.555 191.400 189.805 ;
        RECT 191.905 189.725 192.185 190.525 ;
        RECT 190.980 189.385 192.225 189.555 ;
        RECT 192.395 189.385 192.665 190.355 ;
        RECT 192.925 189.595 193.095 190.355 ;
        RECT 193.275 189.765 193.605 190.525 ;
        RECT 192.925 189.425 193.590 189.595 ;
        RECT 193.775 189.450 194.045 190.355 ;
        RECT 192.055 189.215 192.225 189.385 ;
        RECT 192.435 189.335 192.665 189.385 ;
        RECT 190.080 188.965 190.415 189.215 ;
        RECT 190.585 188.885 191.325 189.215 ;
        RECT 192.055 188.885 192.285 189.215 ;
        RECT 190.585 188.795 190.835 188.885 ;
        RECT 188.695 188.145 188.955 188.650 ;
        RECT 189.150 188.525 189.815 188.695 ;
        RECT 189.135 187.975 189.465 188.355 ;
        RECT 189.645 188.145 189.815 188.525 ;
        RECT 190.100 188.625 190.835 188.795 ;
        RECT 192.055 188.715 192.225 188.885 ;
        RECT 190.100 188.155 190.410 188.625 ;
        RECT 191.485 188.545 192.225 188.715 ;
        RECT 192.495 188.650 192.665 189.335 ;
        RECT 193.420 189.280 193.590 189.425 ;
        RECT 192.855 188.875 193.185 189.245 ;
        RECT 193.420 188.950 193.705 189.280 ;
        RECT 193.420 188.695 193.590 188.950 ;
        RECT 190.580 187.975 191.315 188.455 ;
        RECT 191.485 188.195 191.655 188.545 ;
        RECT 191.825 187.975 192.205 188.375 ;
        RECT 192.395 188.305 192.665 188.650 ;
        RECT 192.925 188.525 193.590 188.695 ;
        RECT 193.875 188.650 194.045 189.450 ;
        RECT 194.305 189.515 194.475 190.355 ;
        RECT 194.645 190.185 195.815 190.355 ;
        RECT 194.645 189.685 194.975 190.185 ;
        RECT 195.485 190.145 195.815 190.185 ;
        RECT 196.005 190.105 196.360 190.525 ;
        RECT 195.145 189.925 195.375 190.015 ;
        RECT 196.530 189.925 196.780 190.355 ;
        RECT 195.145 189.685 196.780 189.925 ;
        RECT 196.950 189.765 197.280 190.525 ;
        RECT 197.450 189.685 197.705 190.355 ;
        RECT 197.495 189.675 197.705 189.685 ;
        RECT 194.305 189.345 197.365 189.515 ;
        RECT 194.220 188.965 194.570 189.175 ;
        RECT 194.740 188.965 195.185 189.165 ;
        RECT 195.355 188.965 195.830 189.165 ;
        RECT 192.925 188.145 193.095 188.525 ;
        RECT 193.275 187.975 193.605 188.355 ;
        RECT 193.785 188.145 194.045 188.650 ;
        RECT 194.305 188.625 195.370 188.795 ;
        RECT 194.305 188.145 194.475 188.625 ;
        RECT 194.645 187.975 194.975 188.455 ;
        RECT 195.200 188.395 195.370 188.625 ;
        RECT 195.550 188.565 195.830 188.965 ;
        RECT 196.100 188.965 196.430 189.165 ;
        RECT 196.600 188.965 196.965 189.165 ;
        RECT 196.100 188.565 196.385 188.965 ;
        RECT 197.195 188.795 197.365 189.345 ;
        RECT 196.565 188.625 197.365 188.795 ;
        RECT 196.565 188.395 196.735 188.625 ;
        RECT 197.535 188.555 197.705 189.675 ;
        RECT 197.520 188.475 197.705 188.555 ;
        RECT 195.200 188.145 196.735 188.395 ;
        RECT 196.905 187.975 197.235 188.455 ;
        RECT 197.450 188.145 197.705 188.475 ;
        RECT 197.895 189.450 198.165 190.355 ;
        RECT 198.335 189.765 198.665 190.525 ;
        RECT 198.845 189.595 199.015 190.355 ;
        RECT 197.895 188.650 198.065 189.450 ;
        RECT 198.350 189.425 199.015 189.595 ;
        RECT 199.275 189.435 202.785 190.525 ;
        RECT 198.350 189.280 198.520 189.425 ;
        RECT 198.235 188.950 198.520 189.280 ;
        RECT 198.350 188.695 198.520 188.950 ;
        RECT 198.755 188.875 199.085 189.245 ;
        RECT 199.275 188.745 200.925 189.265 ;
        RECT 201.095 188.915 202.785 189.435 ;
        RECT 203.875 189.360 204.165 190.525 ;
        RECT 204.335 189.435 207.845 190.525 ;
        RECT 204.335 188.745 205.985 189.265 ;
        RECT 206.155 188.915 207.845 189.435 ;
        RECT 208.475 188.920 208.755 190.355 ;
        RECT 208.925 189.750 209.635 190.525 ;
        RECT 209.805 189.580 210.135 190.355 ;
        RECT 208.985 189.365 210.135 189.580 ;
        RECT 197.895 188.145 198.155 188.650 ;
        RECT 198.350 188.525 199.015 188.695 ;
        RECT 198.335 187.975 198.665 188.355 ;
        RECT 198.845 188.145 199.015 188.525 ;
        RECT 199.275 187.975 202.785 188.745 ;
        RECT 203.875 187.975 204.165 188.700 ;
        RECT 204.335 187.975 207.845 188.745 ;
        RECT 208.475 188.145 208.815 188.920 ;
        RECT 208.985 188.795 209.270 189.365 ;
        RECT 209.455 188.965 209.925 189.195 ;
        RECT 210.330 189.165 210.545 190.280 ;
        RECT 210.725 189.805 211.055 190.525 ;
        RECT 211.235 190.090 216.580 190.525 ;
        RECT 216.755 190.090 222.100 190.525 ;
        RECT 210.835 189.165 211.065 189.505 ;
        RECT 210.095 188.985 210.545 189.165 ;
        RECT 210.095 188.965 210.425 188.985 ;
        RECT 210.735 188.965 211.065 189.165 ;
        RECT 208.985 188.605 209.695 188.795 ;
        RECT 209.395 188.465 209.695 188.605 ;
        RECT 209.885 188.605 211.065 188.795 ;
        RECT 209.885 188.525 210.215 188.605 ;
        RECT 209.395 188.455 209.710 188.465 ;
        RECT 209.395 188.445 209.720 188.455 ;
        RECT 209.395 188.440 209.730 188.445 ;
        RECT 208.985 187.975 209.155 188.435 ;
        RECT 209.395 188.430 209.735 188.440 ;
        RECT 209.395 188.425 209.740 188.430 ;
        RECT 209.395 188.415 209.745 188.425 ;
        RECT 209.395 188.410 209.750 188.415 ;
        RECT 209.395 188.145 209.755 188.410 ;
        RECT 210.385 187.975 210.555 188.435 ;
        RECT 210.725 188.145 211.065 188.605 ;
        RECT 212.820 188.520 213.160 189.350 ;
        RECT 214.640 188.840 214.990 190.090 ;
        RECT 218.340 188.520 218.680 189.350 ;
        RECT 220.160 188.840 220.510 190.090 ;
        RECT 222.275 189.435 225.785 190.525 ;
        RECT 222.275 188.745 223.925 189.265 ;
        RECT 224.095 188.915 225.785 189.435 ;
        RECT 226.415 188.920 226.695 190.355 ;
        RECT 226.865 189.750 227.575 190.525 ;
        RECT 227.745 189.580 228.075 190.355 ;
        RECT 226.925 189.365 228.075 189.580 ;
        RECT 211.235 187.975 216.580 188.520 ;
        RECT 216.755 187.975 222.100 188.520 ;
        RECT 222.275 187.975 225.785 188.745 ;
        RECT 226.415 188.145 226.755 188.920 ;
        RECT 226.925 188.795 227.210 189.365 ;
        RECT 227.395 188.965 227.865 189.195 ;
        RECT 228.270 189.165 228.485 190.280 ;
        RECT 228.665 189.805 228.995 190.525 ;
        RECT 228.775 189.165 229.005 189.505 ;
        RECT 229.635 189.360 229.925 190.525 ;
        RECT 230.095 189.450 230.365 190.355 ;
        RECT 230.535 189.765 230.865 190.525 ;
        RECT 231.045 189.595 231.215 190.355 ;
        RECT 228.035 188.985 228.485 189.165 ;
        RECT 228.035 188.965 228.365 188.985 ;
        RECT 228.675 188.965 229.005 189.165 ;
        RECT 226.925 188.605 227.635 188.795 ;
        RECT 227.335 188.465 227.635 188.605 ;
        RECT 227.825 188.605 229.005 188.795 ;
        RECT 227.825 188.525 228.155 188.605 ;
        RECT 227.335 188.455 227.650 188.465 ;
        RECT 227.335 188.445 227.660 188.455 ;
        RECT 227.335 188.440 227.670 188.445 ;
        RECT 226.925 187.975 227.095 188.435 ;
        RECT 227.335 188.430 227.675 188.440 ;
        RECT 227.335 188.425 227.680 188.430 ;
        RECT 227.335 188.415 227.685 188.425 ;
        RECT 227.335 188.410 227.690 188.415 ;
        RECT 227.335 188.145 227.695 188.410 ;
        RECT 228.325 187.975 228.495 188.435 ;
        RECT 228.665 188.145 229.005 188.605 ;
        RECT 229.635 187.975 229.925 188.700 ;
        RECT 230.095 188.650 230.265 189.450 ;
        RECT 230.550 189.425 231.215 189.595 ;
        RECT 231.565 189.595 231.735 190.355 ;
        RECT 231.915 189.765 232.245 190.525 ;
        RECT 231.565 189.425 232.230 189.595 ;
        RECT 232.415 189.450 232.685 190.355 ;
        RECT 230.550 189.280 230.720 189.425 ;
        RECT 230.435 188.950 230.720 189.280 ;
        RECT 232.060 189.280 232.230 189.425 ;
        RECT 230.550 188.695 230.720 188.950 ;
        RECT 230.955 188.875 231.285 189.245 ;
        RECT 231.495 188.875 231.825 189.245 ;
        RECT 232.060 188.950 232.345 189.280 ;
        RECT 232.060 188.695 232.230 188.950 ;
        RECT 230.095 188.145 230.355 188.650 ;
        RECT 230.550 188.525 231.215 188.695 ;
        RECT 230.535 187.975 230.865 188.355 ;
        RECT 231.045 188.145 231.215 188.525 ;
        RECT 231.565 188.525 232.230 188.695 ;
        RECT 232.515 188.650 232.685 189.450 ;
        RECT 231.565 188.145 231.735 188.525 ;
        RECT 231.915 187.975 232.245 188.355 ;
        RECT 232.425 188.145 232.685 188.650 ;
        RECT 232.855 189.450 233.125 190.355 ;
        RECT 233.295 189.765 233.625 190.525 ;
        RECT 233.805 189.595 233.975 190.355 ;
        RECT 232.855 188.650 233.025 189.450 ;
        RECT 233.310 189.425 233.975 189.595 ;
        RECT 234.235 189.435 237.745 190.525 ;
        RECT 233.310 189.280 233.480 189.425 ;
        RECT 233.195 188.950 233.480 189.280 ;
        RECT 233.310 188.695 233.480 188.950 ;
        RECT 233.715 188.875 234.045 189.245 ;
        RECT 234.235 188.745 235.885 189.265 ;
        RECT 236.055 188.915 237.745 189.435 ;
        RECT 237.915 189.435 239.125 190.525 ;
        RECT 237.915 188.895 238.435 189.435 ;
        RECT 232.855 188.145 233.115 188.650 ;
        RECT 233.310 188.525 233.975 188.695 ;
        RECT 233.295 187.975 233.625 188.355 ;
        RECT 233.805 188.145 233.975 188.525 ;
        RECT 234.235 187.975 237.745 188.745 ;
        RECT 238.605 188.725 239.125 189.265 ;
        RECT 237.915 187.975 239.125 188.725 ;
        RECT 165.150 187.805 239.210 187.975 ;
        RECT 165.235 187.055 166.445 187.805 ;
        RECT 165.235 186.515 165.755 187.055 ;
        RECT 166.615 187.035 168.285 187.805 ;
        RECT 168.545 187.255 168.715 187.635 ;
        RECT 168.895 187.425 169.225 187.805 ;
        RECT 168.545 187.085 169.210 187.255 ;
        RECT 169.405 187.130 169.665 187.635 ;
        RECT 165.925 186.345 166.445 186.885 ;
        RECT 166.615 186.515 167.365 187.035 ;
        RECT 167.535 186.345 168.285 186.865 ;
        RECT 168.475 186.535 168.805 186.905 ;
        RECT 169.040 186.830 169.210 187.085 ;
        RECT 169.040 186.500 169.325 186.830 ;
        RECT 169.040 186.355 169.210 186.500 ;
        RECT 165.235 185.255 166.445 186.345 ;
        RECT 166.615 185.255 168.285 186.345 ;
        RECT 168.545 186.185 169.210 186.355 ;
        RECT 169.495 186.330 169.665 187.130 ;
        RECT 169.925 187.255 170.095 187.635 ;
        RECT 170.275 187.425 170.605 187.805 ;
        RECT 169.925 187.085 170.590 187.255 ;
        RECT 170.785 187.130 171.045 187.635 ;
        RECT 169.855 186.535 170.185 186.905 ;
        RECT 170.420 186.830 170.590 187.085 ;
        RECT 170.420 186.500 170.705 186.830 ;
        RECT 170.420 186.355 170.590 186.500 ;
        RECT 168.545 185.425 168.715 186.185 ;
        RECT 168.895 185.255 169.225 186.015 ;
        RECT 169.395 185.425 169.665 186.330 ;
        RECT 169.925 186.185 170.590 186.355 ;
        RECT 170.875 186.330 171.045 187.130 ;
        RECT 171.305 187.255 171.475 187.635 ;
        RECT 171.690 187.425 172.020 187.805 ;
        RECT 171.305 187.085 172.020 187.255 ;
        RECT 171.215 186.535 171.570 186.905 ;
        RECT 171.850 186.895 172.020 187.085 ;
        RECT 172.190 187.060 172.445 187.635 ;
        RECT 171.850 186.565 172.105 186.895 ;
        RECT 171.850 186.355 172.020 186.565 ;
        RECT 169.925 185.425 170.095 186.185 ;
        RECT 170.275 185.255 170.605 186.015 ;
        RECT 170.775 185.425 171.045 186.330 ;
        RECT 171.305 186.185 172.020 186.355 ;
        RECT 172.275 186.330 172.445 187.060 ;
        RECT 172.620 186.965 172.880 187.805 ;
        RECT 173.210 187.155 173.540 187.620 ;
        RECT 173.710 187.335 173.880 187.805 ;
        RECT 174.050 187.155 174.380 187.635 ;
        RECT 173.210 186.985 174.380 187.155 ;
        RECT 173.055 186.605 173.700 186.815 ;
        RECT 173.870 186.605 174.440 186.815 ;
        RECT 174.610 186.435 174.780 187.635 ;
        RECT 175.320 187.235 175.490 187.440 ;
        RECT 171.305 185.425 171.475 186.185 ;
        RECT 171.690 185.255 172.020 186.015 ;
        RECT 172.190 185.425 172.445 186.330 ;
        RECT 172.620 185.255 172.880 186.405 ;
        RECT 173.270 185.255 173.600 186.355 ;
        RECT 174.075 186.025 174.780 186.435 ;
        RECT 174.950 187.065 175.490 187.235 ;
        RECT 175.770 187.065 175.940 187.805 ;
        RECT 176.205 187.065 176.565 187.440 ;
        RECT 174.950 186.365 175.120 187.065 ;
        RECT 175.290 186.565 175.620 186.895 ;
        RECT 175.790 186.565 176.140 186.895 ;
        RECT 174.950 186.195 175.575 186.365 ;
        RECT 175.790 186.025 176.055 186.565 ;
        RECT 176.310 186.410 176.565 187.065 ;
        RECT 176.890 187.155 177.220 187.620 ;
        RECT 177.390 187.335 177.560 187.805 ;
        RECT 177.730 187.155 178.060 187.635 ;
        RECT 176.890 186.985 178.060 187.155 ;
        RECT 176.735 186.605 177.380 186.815 ;
        RECT 177.550 186.605 178.120 186.815 ;
        RECT 178.290 186.435 178.460 187.635 ;
        RECT 179.000 187.235 179.170 187.440 ;
        RECT 174.075 185.855 176.055 186.025 ;
        RECT 174.075 185.425 174.400 185.855 ;
        RECT 174.570 185.255 174.900 185.675 ;
        RECT 175.645 185.255 176.055 185.685 ;
        RECT 176.225 185.425 176.565 186.410 ;
        RECT 176.950 185.255 177.280 186.355 ;
        RECT 177.755 186.025 178.460 186.435 ;
        RECT 178.630 187.065 179.170 187.235 ;
        RECT 179.450 187.065 179.620 187.805 ;
        RECT 179.885 187.065 180.245 187.440 ;
        RECT 181.425 187.255 181.595 187.635 ;
        RECT 181.775 187.425 182.105 187.805 ;
        RECT 181.425 187.085 182.090 187.255 ;
        RECT 182.285 187.130 182.545 187.635 ;
        RECT 178.630 186.365 178.800 187.065 ;
        RECT 178.970 186.565 179.300 186.895 ;
        RECT 179.470 186.565 179.820 186.895 ;
        RECT 178.630 186.195 179.255 186.365 ;
        RECT 179.470 186.025 179.735 186.565 ;
        RECT 179.990 186.410 180.245 187.065 ;
        RECT 181.355 186.535 181.685 186.905 ;
        RECT 181.920 186.830 182.090 187.085 ;
        RECT 177.755 185.855 179.735 186.025 ;
        RECT 177.755 185.425 178.080 185.855 ;
        RECT 178.250 185.255 178.580 185.675 ;
        RECT 179.325 185.255 179.735 185.685 ;
        RECT 179.905 185.425 180.245 186.410 ;
        RECT 181.920 186.500 182.205 186.830 ;
        RECT 181.920 186.355 182.090 186.500 ;
        RECT 181.425 186.185 182.090 186.355 ;
        RECT 182.375 186.330 182.545 187.130 ;
        RECT 182.805 187.255 182.975 187.635 ;
        RECT 183.155 187.425 183.485 187.805 ;
        RECT 182.805 187.085 183.470 187.255 ;
        RECT 183.665 187.130 183.925 187.635 ;
        RECT 182.735 186.535 183.065 186.905 ;
        RECT 183.300 186.830 183.470 187.085 ;
        RECT 183.300 186.500 183.585 186.830 ;
        RECT 183.300 186.355 183.470 186.500 ;
        RECT 181.425 185.425 181.595 186.185 ;
        RECT 181.775 185.255 182.105 186.015 ;
        RECT 182.275 185.425 182.545 186.330 ;
        RECT 182.805 186.185 183.470 186.355 ;
        RECT 183.755 186.330 183.925 187.130 ;
        RECT 182.805 185.425 182.975 186.185 ;
        RECT 183.155 185.255 183.485 186.015 ;
        RECT 183.655 185.425 183.925 186.330 ;
        RECT 184.095 187.130 184.355 187.635 ;
        RECT 184.535 187.425 184.865 187.805 ;
        RECT 185.045 187.255 185.215 187.635 ;
        RECT 184.095 186.330 184.265 187.130 ;
        RECT 184.550 187.085 185.215 187.255 ;
        RECT 185.565 187.255 185.735 187.635 ;
        RECT 185.915 187.425 186.245 187.805 ;
        RECT 185.565 187.085 186.230 187.255 ;
        RECT 186.425 187.130 186.685 187.635 ;
        RECT 184.550 186.830 184.720 187.085 ;
        RECT 184.435 186.500 184.720 186.830 ;
        RECT 184.955 186.535 185.285 186.905 ;
        RECT 185.495 186.535 185.825 186.905 ;
        RECT 186.060 186.830 186.230 187.085 ;
        RECT 184.550 186.355 184.720 186.500 ;
        RECT 186.060 186.500 186.345 186.830 ;
        RECT 186.060 186.355 186.230 186.500 ;
        RECT 184.095 185.425 184.365 186.330 ;
        RECT 184.550 186.185 185.215 186.355 ;
        RECT 184.535 185.255 184.865 186.015 ;
        RECT 185.045 185.425 185.215 186.185 ;
        RECT 185.565 186.185 186.230 186.355 ;
        RECT 186.515 186.330 186.685 187.130 ;
        RECT 186.945 187.255 187.115 187.635 ;
        RECT 187.295 187.425 187.625 187.805 ;
        RECT 186.945 187.085 187.610 187.255 ;
        RECT 187.805 187.130 188.065 187.635 ;
        RECT 186.875 186.535 187.205 186.905 ;
        RECT 187.440 186.830 187.610 187.085 ;
        RECT 187.440 186.500 187.725 186.830 ;
        RECT 187.440 186.355 187.610 186.500 ;
        RECT 185.565 185.425 185.735 186.185 ;
        RECT 185.915 185.255 186.245 186.015 ;
        RECT 186.415 185.425 186.685 186.330 ;
        RECT 186.945 186.185 187.610 186.355 ;
        RECT 187.895 186.330 188.065 187.130 ;
        RECT 188.260 187.155 188.570 187.625 ;
        RECT 188.740 187.325 189.475 187.805 ;
        RECT 189.645 187.235 189.815 187.585 ;
        RECT 189.985 187.405 190.365 187.805 ;
        RECT 188.260 186.985 188.995 187.155 ;
        RECT 189.645 187.065 190.385 187.235 ;
        RECT 190.555 187.130 190.825 187.475 ;
        RECT 188.745 186.895 188.995 186.985 ;
        RECT 190.215 186.895 190.385 187.065 ;
        RECT 188.240 186.565 188.575 186.815 ;
        RECT 188.745 186.565 189.485 186.895 ;
        RECT 190.215 186.565 190.445 186.895 ;
        RECT 186.945 185.425 187.115 186.185 ;
        RECT 187.295 185.255 187.625 186.015 ;
        RECT 187.795 185.425 188.065 186.330 ;
        RECT 188.240 185.255 188.495 186.395 ;
        RECT 188.745 186.005 188.915 186.565 ;
        RECT 190.215 186.395 190.385 186.565 ;
        RECT 190.655 186.395 190.825 187.130 ;
        RECT 190.995 187.080 191.285 187.805 ;
        RECT 192.465 187.155 192.635 187.635 ;
        RECT 192.805 187.325 193.135 187.805 ;
        RECT 193.360 187.385 194.895 187.635 ;
        RECT 193.360 187.155 193.530 187.385 ;
        RECT 192.465 186.985 193.530 187.155 ;
        RECT 193.710 186.815 193.990 187.215 ;
        RECT 192.380 186.605 192.730 186.815 ;
        RECT 192.900 186.615 193.345 186.815 ;
        RECT 193.515 186.615 193.990 186.815 ;
        RECT 194.260 186.815 194.545 187.215 ;
        RECT 194.725 187.155 194.895 187.385 ;
        RECT 195.065 187.325 195.395 187.805 ;
        RECT 195.610 187.305 195.865 187.635 ;
        RECT 195.655 187.295 195.865 187.305 ;
        RECT 195.680 187.225 195.865 187.295 ;
        RECT 194.725 186.985 195.525 187.155 ;
        RECT 194.260 186.615 194.590 186.815 ;
        RECT 194.760 186.615 195.125 186.815 ;
        RECT 195.355 186.435 195.525 186.985 ;
        RECT 189.140 186.225 190.385 186.395 ;
        RECT 189.140 185.975 189.560 186.225 ;
        RECT 188.690 185.475 189.885 185.805 ;
        RECT 190.065 185.255 190.345 186.055 ;
        RECT 190.555 185.425 190.825 186.395 ;
        RECT 190.995 185.255 191.285 186.420 ;
        RECT 192.465 186.265 195.525 186.435 ;
        RECT 192.465 185.425 192.635 186.265 ;
        RECT 195.695 186.095 195.865 187.225 ;
        RECT 196.145 187.155 196.315 187.635 ;
        RECT 196.485 187.325 196.815 187.805 ;
        RECT 197.040 187.385 198.575 187.635 ;
        RECT 197.040 187.155 197.210 187.385 ;
        RECT 196.145 186.985 197.210 187.155 ;
        RECT 197.390 186.815 197.670 187.215 ;
        RECT 196.060 186.605 196.410 186.815 ;
        RECT 196.580 186.615 197.025 186.815 ;
        RECT 197.195 186.615 197.670 186.815 ;
        RECT 197.940 186.815 198.225 187.215 ;
        RECT 198.405 187.155 198.575 187.385 ;
        RECT 198.745 187.325 199.075 187.805 ;
        RECT 199.290 187.305 199.545 187.635 ;
        RECT 199.360 187.225 199.545 187.305 ;
        RECT 198.405 186.985 199.205 187.155 ;
        RECT 197.940 186.615 198.270 186.815 ;
        RECT 198.440 186.615 198.805 186.815 ;
        RECT 199.035 186.435 199.205 186.985 ;
        RECT 192.805 185.595 193.135 186.095 ;
        RECT 193.305 185.855 194.940 186.095 ;
        RECT 193.305 185.765 193.535 185.855 ;
        RECT 193.645 185.595 193.975 185.635 ;
        RECT 192.805 185.425 193.975 185.595 ;
        RECT 194.165 185.255 194.520 185.675 ;
        RECT 194.690 185.425 194.940 185.855 ;
        RECT 195.110 185.255 195.440 186.015 ;
        RECT 195.610 185.425 195.865 186.095 ;
        RECT 196.145 186.265 199.205 186.435 ;
        RECT 196.145 185.425 196.315 186.265 ;
        RECT 199.375 186.105 199.545 187.225 ;
        RECT 199.825 187.155 199.995 187.635 ;
        RECT 200.165 187.325 200.495 187.805 ;
        RECT 200.720 187.385 202.255 187.635 ;
        RECT 200.720 187.155 200.890 187.385 ;
        RECT 199.825 186.985 200.890 187.155 ;
        RECT 201.070 186.815 201.350 187.215 ;
        RECT 199.740 186.605 200.090 186.815 ;
        RECT 200.260 186.615 200.705 186.815 ;
        RECT 200.875 186.615 201.350 186.815 ;
        RECT 201.620 186.815 201.905 187.215 ;
        RECT 202.085 187.155 202.255 187.385 ;
        RECT 202.425 187.325 202.755 187.805 ;
        RECT 202.970 187.305 203.225 187.635 ;
        RECT 203.015 187.295 203.225 187.305 ;
        RECT 203.040 187.225 203.225 187.295 ;
        RECT 203.415 187.260 208.760 187.805 ;
        RECT 202.085 186.985 202.885 187.155 ;
        RECT 201.620 186.615 201.950 186.815 ;
        RECT 202.120 186.615 202.485 186.815 ;
        RECT 202.715 186.435 202.885 186.985 ;
        RECT 199.335 186.095 199.545 186.105 ;
        RECT 196.485 185.595 196.815 186.095 ;
        RECT 196.985 185.855 198.620 186.095 ;
        RECT 196.985 185.765 197.215 185.855 ;
        RECT 197.325 185.595 197.655 185.635 ;
        RECT 196.485 185.425 197.655 185.595 ;
        RECT 197.845 185.255 198.200 185.675 ;
        RECT 198.370 185.425 198.620 185.855 ;
        RECT 198.790 185.255 199.120 186.015 ;
        RECT 199.290 185.425 199.545 186.095 ;
        RECT 199.825 186.265 202.885 186.435 ;
        RECT 199.825 185.425 199.995 186.265 ;
        RECT 203.055 186.095 203.225 187.225 ;
        RECT 205.000 186.430 205.340 187.260 ;
        RECT 209.025 187.255 209.195 187.635 ;
        RECT 209.410 187.425 209.740 187.805 ;
        RECT 209.025 187.085 209.740 187.255 ;
        RECT 200.165 185.595 200.495 186.095 ;
        RECT 200.665 185.855 202.300 186.095 ;
        RECT 200.665 185.765 200.895 185.855 ;
        RECT 201.005 185.595 201.335 185.635 ;
        RECT 200.165 185.425 201.335 185.595 ;
        RECT 201.525 185.255 201.880 185.675 ;
        RECT 202.050 185.425 202.300 185.855 ;
        RECT 202.470 185.255 202.800 186.015 ;
        RECT 202.970 185.425 203.225 186.095 ;
        RECT 206.820 185.690 207.170 186.940 ;
        RECT 208.935 186.535 209.290 186.905 ;
        RECT 209.570 186.895 209.740 187.085 ;
        RECT 209.910 187.060 210.165 187.635 ;
        RECT 209.570 186.565 209.825 186.895 ;
        RECT 209.570 186.355 209.740 186.565 ;
        RECT 209.025 186.185 209.740 186.355 ;
        RECT 209.995 186.330 210.165 187.060 ;
        RECT 210.340 186.965 210.600 187.805 ;
        RECT 210.865 187.255 211.035 187.635 ;
        RECT 211.215 187.425 211.545 187.805 ;
        RECT 210.865 187.085 211.530 187.255 ;
        RECT 211.725 187.130 211.985 187.635 ;
        RECT 210.795 186.535 211.125 186.905 ;
        RECT 211.360 186.830 211.530 187.085 ;
        RECT 211.360 186.500 211.645 186.830 ;
        RECT 203.415 185.255 208.760 185.690 ;
        RECT 209.025 185.425 209.195 186.185 ;
        RECT 209.410 185.255 209.740 186.015 ;
        RECT 209.910 185.425 210.165 186.330 ;
        RECT 210.340 185.255 210.600 186.405 ;
        RECT 211.360 186.355 211.530 186.500 ;
        RECT 210.865 186.185 211.530 186.355 ;
        RECT 211.815 186.330 211.985 187.130 ;
        RECT 212.245 187.255 212.415 187.635 ;
        RECT 212.595 187.425 212.925 187.805 ;
        RECT 212.245 187.085 212.910 187.255 ;
        RECT 213.105 187.130 213.365 187.635 ;
        RECT 212.175 186.535 212.505 186.905 ;
        RECT 212.740 186.830 212.910 187.085 ;
        RECT 212.740 186.500 213.025 186.830 ;
        RECT 212.740 186.355 212.910 186.500 ;
        RECT 210.865 185.425 211.035 186.185 ;
        RECT 211.215 185.255 211.545 186.015 ;
        RECT 211.715 185.425 211.985 186.330 ;
        RECT 212.245 186.185 212.910 186.355 ;
        RECT 213.195 186.330 213.365 187.130 ;
        RECT 213.625 187.255 213.795 187.635 ;
        RECT 213.975 187.425 214.305 187.805 ;
        RECT 213.625 187.085 214.290 187.255 ;
        RECT 214.485 187.130 214.745 187.635 ;
        RECT 213.555 186.535 213.885 186.905 ;
        RECT 214.120 186.830 214.290 187.085 ;
        RECT 214.120 186.500 214.405 186.830 ;
        RECT 214.120 186.355 214.290 186.500 ;
        RECT 212.245 185.425 212.415 186.185 ;
        RECT 212.595 185.255 212.925 186.015 ;
        RECT 213.095 185.425 213.365 186.330 ;
        RECT 213.625 186.185 214.290 186.355 ;
        RECT 214.575 186.330 214.745 187.130 ;
        RECT 215.005 187.255 215.175 187.635 ;
        RECT 215.355 187.425 215.685 187.805 ;
        RECT 215.005 187.085 215.670 187.255 ;
        RECT 215.865 187.130 216.125 187.635 ;
        RECT 214.935 186.535 215.265 186.905 ;
        RECT 215.500 186.830 215.670 187.085 ;
        RECT 215.500 186.500 215.785 186.830 ;
        RECT 215.500 186.355 215.670 186.500 ;
        RECT 213.625 185.425 213.795 186.185 ;
        RECT 213.975 185.255 214.305 186.015 ;
        RECT 214.475 185.425 214.745 186.330 ;
        RECT 215.005 186.185 215.670 186.355 ;
        RECT 215.955 186.330 216.125 187.130 ;
        RECT 216.755 187.080 217.045 187.805 ;
        RECT 217.215 186.860 217.555 187.635 ;
        RECT 217.725 187.345 217.895 187.805 ;
        RECT 218.135 187.370 218.495 187.635 ;
        RECT 218.135 187.365 218.490 187.370 ;
        RECT 218.135 187.355 218.485 187.365 ;
        RECT 218.135 187.350 218.480 187.355 ;
        RECT 218.135 187.340 218.475 187.350 ;
        RECT 219.125 187.345 219.295 187.805 ;
        RECT 218.135 187.335 218.470 187.340 ;
        RECT 218.135 187.325 218.460 187.335 ;
        RECT 218.135 187.315 218.450 187.325 ;
        RECT 218.135 187.175 218.435 187.315 ;
        RECT 217.725 186.985 218.435 187.175 ;
        RECT 218.625 187.175 218.955 187.255 ;
        RECT 219.465 187.175 219.805 187.635 ;
        RECT 218.625 186.985 219.805 187.175 ;
        RECT 220.065 187.255 220.235 187.635 ;
        RECT 220.415 187.425 220.745 187.805 ;
        RECT 220.065 187.085 220.730 187.255 ;
        RECT 220.925 187.130 221.185 187.635 ;
        RECT 215.005 185.425 215.175 186.185 ;
        RECT 215.355 185.255 215.685 186.015 ;
        RECT 215.855 185.425 216.125 186.330 ;
        RECT 216.755 185.255 217.045 186.420 ;
        RECT 217.215 185.425 217.495 186.860 ;
        RECT 217.725 186.415 218.010 186.985 ;
        RECT 218.195 186.585 218.665 186.815 ;
        RECT 218.835 186.795 219.165 186.815 ;
        RECT 218.835 186.615 219.285 186.795 ;
        RECT 219.475 186.615 219.805 186.815 ;
        RECT 217.725 186.200 218.875 186.415 ;
        RECT 217.665 185.255 218.375 186.030 ;
        RECT 218.545 185.425 218.875 186.200 ;
        RECT 219.070 185.500 219.285 186.615 ;
        RECT 219.575 186.275 219.805 186.615 ;
        RECT 219.995 186.535 220.325 186.905 ;
        RECT 220.560 186.830 220.730 187.085 ;
        RECT 220.560 186.500 220.845 186.830 ;
        RECT 220.560 186.355 220.730 186.500 ;
        RECT 220.065 186.185 220.730 186.355 ;
        RECT 221.015 186.330 221.185 187.130 ;
        RECT 219.465 185.255 219.795 185.975 ;
        RECT 220.065 185.425 220.235 186.185 ;
        RECT 220.415 185.255 220.745 186.015 ;
        RECT 220.915 185.425 221.185 186.330 ;
        RECT 221.355 187.130 221.615 187.635 ;
        RECT 221.795 187.425 222.125 187.805 ;
        RECT 222.305 187.255 222.475 187.635 ;
        RECT 221.355 186.330 221.525 187.130 ;
        RECT 221.810 187.085 222.475 187.255 ;
        RECT 222.825 187.255 222.995 187.630 ;
        RECT 223.165 187.425 223.495 187.805 ;
        RECT 223.665 187.465 224.740 187.635 ;
        RECT 223.665 187.255 223.835 187.465 ;
        RECT 222.825 187.085 223.835 187.255 ;
        RECT 224.060 187.125 224.400 187.295 ;
        RECT 224.570 187.130 224.740 187.465 ;
        RECT 221.810 186.830 221.980 187.085 ;
        RECT 224.060 186.955 224.350 187.125 ;
        RECT 221.695 186.500 221.980 186.830 ;
        RECT 222.215 186.535 222.545 186.905 ;
        RECT 221.810 186.355 221.980 186.500 ;
        RECT 222.800 186.445 223.145 186.895 ;
        RECT 221.355 185.425 221.625 186.330 ;
        RECT 221.810 186.185 222.475 186.355 ;
        RECT 222.795 186.275 223.145 186.445 ;
        RECT 223.455 186.275 223.890 186.895 ;
        RECT 224.060 186.435 224.230 186.955 ;
        RECT 224.910 186.785 225.270 187.460 ;
        RECT 225.450 187.085 225.740 187.805 ;
        RECT 226.030 187.465 227.630 187.635 ;
        RECT 226.030 187.095 226.200 187.465 ;
        RECT 227.275 187.425 227.630 187.465 ;
        RECT 227.800 187.345 227.970 187.805 ;
        RECT 226.370 187.045 226.700 187.295 ;
        RECT 226.385 186.970 226.700 187.045 ;
        RECT 226.870 187.175 227.040 187.295 ;
        RECT 228.145 187.175 228.390 187.595 ;
        RECT 228.660 187.425 228.990 187.805 ;
        RECT 229.160 187.235 229.335 187.565 ;
        RECT 229.680 187.475 229.850 187.635 ;
        RECT 229.680 187.305 230.210 187.475 ;
        RECT 230.380 187.465 231.375 187.635 ;
        RECT 230.380 187.305 230.550 187.465 ;
        RECT 226.870 187.005 228.390 187.175 ;
        RECT 224.730 186.605 225.270 186.785 ;
        RECT 224.910 186.495 225.270 186.605 ;
        RECT 224.060 186.265 224.695 186.435 ;
        RECT 224.910 186.265 225.715 186.495 ;
        RECT 221.795 185.255 222.125 186.015 ;
        RECT 222.305 185.425 222.475 186.185 ;
        RECT 222.825 185.925 224.355 186.095 ;
        RECT 222.825 185.425 222.995 185.925 ;
        RECT 224.185 185.765 224.355 185.925 ;
        RECT 224.525 185.935 224.695 186.265 ;
        RECT 224.525 185.765 224.855 185.935 ;
        RECT 223.165 185.255 223.495 185.635 ;
        RECT 223.665 185.595 223.835 185.755 ;
        RECT 225.025 185.595 225.195 186.095 ;
        RECT 223.665 185.425 225.195 185.595 ;
        RECT 225.365 185.425 225.715 186.265 ;
        RECT 225.915 185.895 226.215 186.895 ;
        RECT 226.385 186.445 226.555 186.970 ;
        RECT 226.870 186.965 227.040 187.005 ;
        RECT 226.725 186.785 227.055 186.795 ;
        RECT 227.450 186.785 227.695 186.835 ;
        RECT 226.725 186.625 227.110 186.785 ;
        RECT 226.940 186.615 227.110 186.625 ;
        RECT 227.395 186.615 227.695 186.785 ;
        RECT 226.385 186.275 227.145 186.445 ;
        RECT 225.885 185.255 226.215 185.635 ;
        RECT 226.475 185.595 226.645 186.105 ;
        RECT 226.815 185.765 227.145 186.275 ;
        RECT 227.450 186.215 227.695 186.615 ;
        RECT 227.900 186.785 228.230 186.835 ;
        RECT 227.900 186.615 228.255 186.785 ;
        RECT 227.900 186.215 228.230 186.615 ;
        RECT 228.705 186.215 228.995 186.895 ;
        RECT 229.165 186.785 229.335 187.235 ;
        RECT 229.630 186.955 229.870 187.125 ;
        RECT 229.165 186.615 229.455 186.785 ;
        RECT 227.315 185.805 228.380 185.975 ;
        RECT 227.315 185.595 227.485 185.805 ;
        RECT 226.475 185.425 227.485 185.595 ;
        RECT 227.710 185.255 228.040 185.635 ;
        RECT 228.210 185.425 228.380 185.805 ;
        RECT 229.165 185.755 229.335 186.615 ;
        RECT 228.630 185.255 228.980 185.635 ;
        RECT 229.150 185.425 229.335 185.755 ;
        RECT 229.630 185.755 229.800 186.955 ;
        RECT 230.040 186.135 230.210 187.305 ;
        RECT 230.860 187.125 231.035 187.295 ;
        RECT 230.620 186.965 231.035 187.125 ;
        RECT 231.205 187.175 231.375 187.465 ;
        RECT 231.545 187.345 231.715 187.805 ;
        RECT 231.205 187.005 231.775 187.175 ;
        RECT 230.620 186.955 231.030 186.965 ;
        RECT 230.840 186.615 231.295 186.785 ;
        RECT 231.605 186.225 231.775 187.005 ;
        RECT 230.040 185.905 230.825 186.135 ;
        RECT 230.495 185.765 230.825 185.905 ;
        RECT 231.125 186.055 231.775 186.225 ;
        RECT 229.630 185.425 229.840 185.755 ;
        RECT 230.010 185.595 230.340 185.635 ;
        RECT 231.125 185.595 231.295 186.055 ;
        RECT 230.010 185.425 231.295 185.595 ;
        RECT 231.465 185.255 231.795 185.635 ;
        RECT 231.965 185.425 232.225 187.635 ;
        RECT 232.395 187.175 232.735 187.635 ;
        RECT 232.905 187.345 233.075 187.805 ;
        RECT 233.705 187.370 234.065 187.635 ;
        RECT 233.710 187.365 234.065 187.370 ;
        RECT 233.715 187.355 234.065 187.365 ;
        RECT 233.720 187.350 234.065 187.355 ;
        RECT 233.725 187.340 234.065 187.350 ;
        RECT 234.305 187.345 234.475 187.805 ;
        RECT 233.730 187.335 234.065 187.340 ;
        RECT 233.740 187.325 234.065 187.335 ;
        RECT 233.750 187.315 234.065 187.325 ;
        RECT 233.245 187.175 233.575 187.255 ;
        RECT 232.395 186.985 233.575 187.175 ;
        RECT 233.765 187.175 234.065 187.315 ;
        RECT 233.765 186.985 234.475 187.175 ;
        RECT 232.395 186.615 232.725 186.815 ;
        RECT 233.035 186.795 233.365 186.815 ;
        RECT 232.915 186.615 233.365 186.795 ;
        RECT 232.395 186.275 232.625 186.615 ;
        RECT 232.405 185.255 232.735 185.975 ;
        RECT 232.915 185.500 233.130 186.615 ;
        RECT 233.535 186.585 234.005 186.815 ;
        RECT 234.190 186.415 234.475 186.985 ;
        RECT 234.645 186.860 234.985 187.635 ;
        RECT 233.325 186.200 234.475 186.415 ;
        RECT 233.325 185.425 233.655 186.200 ;
        RECT 233.825 185.255 234.535 186.030 ;
        RECT 234.705 185.425 234.985 186.860 ;
        RECT 235.155 187.130 235.415 187.635 ;
        RECT 235.595 187.425 235.925 187.805 ;
        RECT 236.105 187.255 236.275 187.635 ;
        RECT 235.155 186.330 235.325 187.130 ;
        RECT 235.610 187.085 236.275 187.255 ;
        RECT 236.535 187.130 236.795 187.635 ;
        RECT 236.975 187.425 237.305 187.805 ;
        RECT 237.485 187.255 237.655 187.635 ;
        RECT 235.610 186.830 235.780 187.085 ;
        RECT 235.495 186.500 235.780 186.830 ;
        RECT 236.015 186.535 236.345 186.905 ;
        RECT 235.610 186.355 235.780 186.500 ;
        RECT 235.155 185.425 235.425 186.330 ;
        RECT 235.610 186.185 236.275 186.355 ;
        RECT 235.595 185.255 235.925 186.015 ;
        RECT 236.105 185.425 236.275 186.185 ;
        RECT 236.535 186.330 236.705 187.130 ;
        RECT 236.990 187.085 237.655 187.255 ;
        RECT 236.990 186.830 237.160 187.085 ;
        RECT 237.915 187.055 239.125 187.805 ;
        RECT 236.875 186.500 237.160 186.830 ;
        RECT 237.395 186.535 237.725 186.905 ;
        RECT 236.990 186.355 237.160 186.500 ;
        RECT 236.535 185.425 236.805 186.330 ;
        RECT 236.990 186.185 237.655 186.355 ;
        RECT 236.975 185.255 237.305 186.015 ;
        RECT 237.485 185.425 237.655 186.185 ;
        RECT 237.915 186.345 238.435 186.885 ;
        RECT 238.605 186.515 239.125 187.055 ;
        RECT 237.915 185.255 239.125 186.345 ;
        RECT 165.150 185.085 239.210 185.255 ;
        RECT 108.630 184.880 153.130 185.050 ;
        RECT 165.235 183.995 166.445 185.085 ;
        RECT 165.235 183.285 165.755 183.825 ;
        RECT 165.925 183.455 166.445 183.995 ;
        RECT 166.705 184.155 166.875 184.915 ;
        RECT 167.055 184.325 167.385 185.085 ;
        RECT 166.705 183.985 167.370 184.155 ;
        RECT 167.555 184.010 167.825 184.915 ;
        RECT 167.200 183.840 167.370 183.985 ;
        RECT 166.635 183.435 166.965 183.805 ;
        RECT 167.200 183.510 167.485 183.840 ;
        RECT 165.235 182.535 166.445 183.285 ;
        RECT 167.200 183.255 167.370 183.510 ;
        RECT 166.705 183.085 167.370 183.255 ;
        RECT 167.655 183.210 167.825 184.010 ;
        RECT 168.085 184.155 168.255 184.915 ;
        RECT 168.435 184.325 168.765 185.085 ;
        RECT 168.085 183.985 168.750 184.155 ;
        RECT 168.935 184.010 169.205 184.915 ;
        RECT 168.580 183.840 168.750 183.985 ;
        RECT 168.015 183.435 168.345 183.805 ;
        RECT 168.580 183.510 168.865 183.840 ;
        RECT 168.580 183.255 168.750 183.510 ;
        RECT 166.705 182.705 166.875 183.085 ;
        RECT 167.055 182.535 167.385 182.915 ;
        RECT 167.565 182.705 167.825 183.210 ;
        RECT 168.085 183.085 168.750 183.255 ;
        RECT 169.035 183.210 169.205 184.010 ;
        RECT 169.465 184.155 169.635 184.915 ;
        RECT 169.815 184.325 170.145 185.085 ;
        RECT 169.465 183.985 170.130 184.155 ;
        RECT 170.315 184.010 170.585 184.915 ;
        RECT 169.960 183.840 170.130 183.985 ;
        RECT 169.395 183.435 169.725 183.805 ;
        RECT 169.960 183.510 170.245 183.840 ;
        RECT 169.960 183.255 170.130 183.510 ;
        RECT 168.085 182.705 168.255 183.085 ;
        RECT 168.435 182.535 168.765 182.915 ;
        RECT 168.945 182.705 169.205 183.210 ;
        RECT 169.465 183.085 170.130 183.255 ;
        RECT 170.415 183.210 170.585 184.010 ;
        RECT 170.970 183.985 171.300 185.085 ;
        RECT 171.775 184.485 172.100 184.915 ;
        RECT 172.270 184.665 172.600 185.085 ;
        RECT 173.345 184.655 173.755 185.085 ;
        RECT 171.775 184.315 173.755 184.485 ;
        RECT 171.775 183.905 172.480 184.315 ;
        RECT 170.755 183.525 171.400 183.735 ;
        RECT 171.570 183.525 172.140 183.735 ;
        RECT 169.465 182.705 169.635 183.085 ;
        RECT 169.815 182.535 170.145 182.915 ;
        RECT 170.325 182.705 170.585 183.210 ;
        RECT 170.910 183.185 172.080 183.355 ;
        RECT 170.910 182.720 171.240 183.185 ;
        RECT 171.410 182.535 171.580 183.005 ;
        RECT 171.750 182.705 172.080 183.185 ;
        RECT 172.310 182.705 172.480 183.905 ;
        RECT 172.650 183.975 173.275 184.145 ;
        RECT 172.650 183.275 172.820 183.975 ;
        RECT 173.490 183.775 173.755 184.315 ;
        RECT 173.925 183.930 174.265 184.915 ;
        RECT 172.990 183.445 173.320 183.775 ;
        RECT 173.490 183.445 173.840 183.775 ;
        RECT 174.010 183.275 174.265 183.930 ;
        RECT 172.650 183.105 173.190 183.275 ;
        RECT 173.020 182.900 173.190 183.105 ;
        RECT 173.470 182.535 173.640 183.275 ;
        RECT 173.905 182.900 174.265 183.275 ;
        RECT 174.455 184.245 174.710 184.915 ;
        RECT 174.880 184.325 175.210 185.085 ;
        RECT 175.380 184.485 175.630 184.915 ;
        RECT 175.800 184.665 176.155 185.085 ;
        RECT 176.345 184.745 177.515 184.915 ;
        RECT 176.345 184.705 176.675 184.745 ;
        RECT 176.785 184.485 177.015 184.575 ;
        RECT 175.380 184.245 177.015 184.485 ;
        RECT 177.185 184.245 177.515 184.745 ;
        RECT 174.455 184.235 174.665 184.245 ;
        RECT 174.455 183.115 174.625 184.235 ;
        RECT 177.685 184.075 177.855 184.915 ;
        RECT 174.795 183.905 177.855 184.075 ;
        RECT 178.115 183.920 178.405 185.085 ;
        RECT 178.595 184.245 178.850 184.915 ;
        RECT 179.020 184.325 179.350 185.085 ;
        RECT 179.520 184.485 179.770 184.915 ;
        RECT 179.940 184.665 180.295 185.085 ;
        RECT 180.485 184.745 181.655 184.915 ;
        RECT 180.485 184.705 180.815 184.745 ;
        RECT 180.925 184.485 181.155 184.575 ;
        RECT 179.520 184.245 181.155 184.485 ;
        RECT 181.325 184.245 181.655 184.745 ;
        RECT 174.795 183.355 174.965 183.905 ;
        RECT 175.195 183.525 175.560 183.725 ;
        RECT 175.730 183.525 176.060 183.725 ;
        RECT 174.795 183.185 175.595 183.355 ;
        RECT 174.455 183.035 174.640 183.115 ;
        RECT 174.455 182.705 174.710 183.035 ;
        RECT 174.925 182.535 175.255 183.015 ;
        RECT 175.425 182.955 175.595 183.185 ;
        RECT 175.775 183.125 176.060 183.525 ;
        RECT 176.330 183.525 176.805 183.725 ;
        RECT 176.975 183.525 177.420 183.725 ;
        RECT 177.590 183.525 177.940 183.735 ;
        RECT 176.330 183.125 176.610 183.525 ;
        RECT 176.790 183.185 177.855 183.355 ;
        RECT 176.790 182.955 176.960 183.185 ;
        RECT 175.425 182.705 176.960 182.955 ;
        RECT 177.185 182.535 177.515 183.015 ;
        RECT 177.685 182.705 177.855 183.185 ;
        RECT 178.115 182.535 178.405 183.260 ;
        RECT 178.595 183.115 178.765 184.245 ;
        RECT 181.825 184.075 181.995 184.915 ;
        RECT 178.935 183.905 181.995 184.075 ;
        RECT 182.470 183.985 182.800 185.085 ;
        RECT 183.275 184.485 183.600 184.915 ;
        RECT 183.770 184.665 184.100 185.085 ;
        RECT 184.845 184.655 185.255 185.085 ;
        RECT 183.275 184.315 185.255 184.485 ;
        RECT 183.275 183.905 183.980 184.315 ;
        RECT 178.935 183.355 179.105 183.905 ;
        RECT 179.335 183.525 179.700 183.725 ;
        RECT 179.870 183.525 180.200 183.725 ;
        RECT 178.935 183.185 179.735 183.355 ;
        RECT 178.595 183.035 178.780 183.115 ;
        RECT 178.595 182.705 178.850 183.035 ;
        RECT 179.065 182.535 179.395 183.015 ;
        RECT 179.565 182.955 179.735 183.185 ;
        RECT 179.915 183.125 180.200 183.525 ;
        RECT 180.470 183.525 180.945 183.725 ;
        RECT 181.115 183.525 181.560 183.725 ;
        RECT 181.730 183.525 182.080 183.735 ;
        RECT 182.255 183.525 182.900 183.735 ;
        RECT 183.070 183.525 183.640 183.735 ;
        RECT 180.470 183.125 180.750 183.525 ;
        RECT 180.930 183.185 181.995 183.355 ;
        RECT 180.930 182.955 181.100 183.185 ;
        RECT 179.565 182.705 181.100 182.955 ;
        RECT 181.325 182.535 181.655 183.015 ;
        RECT 181.825 182.705 181.995 183.185 ;
        RECT 182.410 183.185 183.580 183.355 ;
        RECT 182.410 182.720 182.740 183.185 ;
        RECT 182.910 182.535 183.080 183.005 ;
        RECT 183.250 182.705 183.580 183.185 ;
        RECT 183.810 182.705 183.980 183.905 ;
        RECT 184.150 183.975 184.775 184.145 ;
        RECT 184.150 183.275 184.320 183.975 ;
        RECT 184.990 183.775 185.255 184.315 ;
        RECT 185.425 183.930 185.765 184.915 ;
        RECT 186.945 184.155 187.115 184.915 ;
        RECT 187.295 184.325 187.625 185.085 ;
        RECT 186.945 183.985 187.610 184.155 ;
        RECT 187.795 184.010 188.065 184.915 ;
        RECT 184.490 183.445 184.820 183.775 ;
        RECT 184.990 183.445 185.340 183.775 ;
        RECT 185.510 183.275 185.765 183.930 ;
        RECT 187.440 183.840 187.610 183.985 ;
        RECT 186.875 183.435 187.205 183.805 ;
        RECT 187.440 183.510 187.725 183.840 ;
        RECT 184.150 183.105 184.690 183.275 ;
        RECT 184.520 182.900 184.690 183.105 ;
        RECT 184.970 182.535 185.140 183.275 ;
        RECT 185.405 182.900 185.765 183.275 ;
        RECT 187.440 183.255 187.610 183.510 ;
        RECT 186.945 183.085 187.610 183.255 ;
        RECT 187.895 183.210 188.065 184.010 ;
        RECT 188.240 183.945 188.495 185.085 ;
        RECT 188.690 184.535 189.885 184.865 ;
        RECT 188.745 183.775 188.915 184.335 ;
        RECT 189.140 184.115 189.560 184.365 ;
        RECT 190.065 184.285 190.345 185.085 ;
        RECT 189.140 183.945 190.385 184.115 ;
        RECT 190.555 183.945 190.825 184.915 ;
        RECT 191.000 183.945 191.255 185.085 ;
        RECT 191.450 184.535 192.645 184.865 ;
        RECT 190.215 183.775 190.385 183.945 ;
        RECT 188.240 183.525 188.575 183.775 ;
        RECT 188.745 183.445 189.485 183.775 ;
        RECT 190.215 183.445 190.445 183.775 ;
        RECT 188.745 183.355 188.995 183.445 ;
        RECT 186.945 182.705 187.115 183.085 ;
        RECT 187.295 182.535 187.625 182.915 ;
        RECT 187.805 182.705 188.065 183.210 ;
        RECT 188.260 183.185 188.995 183.355 ;
        RECT 190.215 183.275 190.385 183.445 ;
        RECT 188.260 182.715 188.570 183.185 ;
        RECT 189.645 183.105 190.385 183.275 ;
        RECT 190.655 183.210 190.825 183.945 ;
        RECT 191.505 183.775 191.675 184.335 ;
        RECT 191.900 184.115 192.320 184.365 ;
        RECT 192.825 184.285 193.105 185.085 ;
        RECT 191.900 183.945 193.145 184.115 ;
        RECT 193.315 183.945 193.585 184.915 ;
        RECT 192.975 183.775 193.145 183.945 ;
        RECT 191.000 183.525 191.335 183.775 ;
        RECT 191.505 183.445 192.245 183.775 ;
        RECT 192.975 183.445 193.205 183.775 ;
        RECT 191.505 183.355 191.755 183.445 ;
        RECT 188.740 182.535 189.475 183.015 ;
        RECT 189.645 182.755 189.815 183.105 ;
        RECT 189.985 182.535 190.365 182.935 ;
        RECT 190.555 182.865 190.825 183.210 ;
        RECT 191.020 183.185 191.755 183.355 ;
        RECT 192.975 183.275 193.145 183.445 ;
        RECT 191.020 182.715 191.330 183.185 ;
        RECT 192.405 183.105 193.145 183.275 ;
        RECT 193.415 183.210 193.585 183.945 ;
        RECT 191.500 182.535 192.235 183.015 ;
        RECT 192.405 182.755 192.575 183.105 ;
        RECT 192.745 182.535 193.125 182.935 ;
        RECT 193.315 182.865 193.585 183.210 ;
        RECT 194.680 183.945 195.015 184.915 ;
        RECT 195.185 183.945 195.355 185.085 ;
        RECT 195.525 184.745 197.555 184.915 ;
        RECT 194.680 183.275 194.850 183.945 ;
        RECT 195.525 183.775 195.695 184.745 ;
        RECT 195.020 183.445 195.275 183.775 ;
        RECT 195.500 183.445 195.695 183.775 ;
        RECT 195.865 184.405 196.990 184.575 ;
        RECT 195.105 183.275 195.275 183.445 ;
        RECT 195.865 183.275 196.035 184.405 ;
        RECT 194.680 182.705 194.935 183.275 ;
        RECT 195.105 183.105 196.035 183.275 ;
        RECT 196.205 184.065 197.215 184.235 ;
        RECT 196.205 183.265 196.375 184.065 ;
        RECT 196.580 183.385 196.855 183.865 ;
        RECT 196.575 183.215 196.855 183.385 ;
        RECT 195.860 183.070 196.035 183.105 ;
        RECT 195.105 182.535 195.435 182.935 ;
        RECT 195.860 182.705 196.390 183.070 ;
        RECT 196.580 182.705 196.855 183.215 ;
        RECT 197.025 182.705 197.215 184.065 ;
        RECT 197.385 184.080 197.555 184.745 ;
        RECT 197.725 184.325 197.895 185.085 ;
        RECT 198.130 184.325 198.645 184.735 ;
        RECT 197.385 183.890 198.135 184.080 ;
        RECT 198.305 183.515 198.645 184.325 ;
        RECT 197.415 183.345 198.645 183.515 ;
        RECT 198.815 184.115 199.125 184.915 ;
        RECT 199.295 184.285 199.605 185.085 ;
        RECT 199.775 184.455 200.035 184.915 ;
        RECT 200.205 184.625 200.460 185.085 ;
        RECT 200.635 184.455 200.895 184.915 ;
        RECT 199.775 184.285 200.895 184.455 ;
        RECT 198.815 183.945 199.845 184.115 ;
        RECT 197.395 182.535 197.905 183.070 ;
        RECT 198.125 182.740 198.370 183.345 ;
        RECT 198.815 183.035 198.985 183.945 ;
        RECT 199.155 183.205 199.505 183.775 ;
        RECT 199.675 183.695 199.845 183.945 ;
        RECT 200.635 184.035 200.895 184.285 ;
        RECT 201.065 184.215 201.350 185.085 ;
        RECT 200.635 183.865 201.390 184.035 ;
        RECT 199.675 183.525 200.815 183.695 ;
        RECT 200.985 183.355 201.390 183.865 ;
        RECT 199.740 183.185 201.390 183.355 ;
        RECT 202.035 184.010 202.305 184.915 ;
        RECT 202.475 184.325 202.805 185.085 ;
        RECT 202.985 184.155 203.155 184.915 ;
        RECT 202.035 183.210 202.205 184.010 ;
        RECT 202.490 183.985 203.155 184.155 ;
        RECT 202.490 183.840 202.660 183.985 ;
        RECT 203.875 183.920 204.165 185.085 ;
        RECT 204.425 184.155 204.595 184.915 ;
        RECT 204.775 184.325 205.105 185.085 ;
        RECT 204.425 183.985 205.090 184.155 ;
        RECT 205.275 184.010 205.545 184.915 ;
        RECT 202.375 183.510 202.660 183.840 ;
        RECT 204.920 183.840 205.090 183.985 ;
        RECT 202.490 183.255 202.660 183.510 ;
        RECT 202.895 183.435 203.225 183.805 ;
        RECT 204.355 183.435 204.685 183.805 ;
        RECT 204.920 183.510 205.205 183.840 ;
        RECT 198.815 182.705 199.115 183.035 ;
        RECT 199.285 182.535 199.560 183.015 ;
        RECT 199.740 182.795 200.035 183.185 ;
        RECT 200.205 182.535 200.460 183.015 ;
        RECT 200.635 182.795 200.895 183.185 ;
        RECT 201.065 182.535 201.345 183.015 ;
        RECT 202.035 182.705 202.295 183.210 ;
        RECT 202.490 183.085 203.155 183.255 ;
        RECT 202.475 182.535 202.805 182.915 ;
        RECT 202.985 182.705 203.155 183.085 ;
        RECT 203.875 182.535 204.165 183.260 ;
        RECT 204.920 183.255 205.090 183.510 ;
        RECT 204.425 183.085 205.090 183.255 ;
        RECT 205.375 183.210 205.545 184.010 ;
        RECT 206.265 184.155 206.435 184.915 ;
        RECT 206.615 184.325 206.945 185.085 ;
        RECT 206.265 183.985 206.930 184.155 ;
        RECT 207.115 184.010 207.385 184.915 ;
        RECT 206.760 183.840 206.930 183.985 ;
        RECT 206.195 183.435 206.525 183.805 ;
        RECT 206.760 183.510 207.045 183.840 ;
        RECT 206.760 183.255 206.930 183.510 ;
        RECT 204.425 182.705 204.595 183.085 ;
        RECT 204.775 182.535 205.105 182.915 ;
        RECT 205.285 182.705 205.545 183.210 ;
        RECT 206.265 183.085 206.930 183.255 ;
        RECT 207.215 183.210 207.385 184.010 ;
        RECT 206.265 182.705 206.435 183.085 ;
        RECT 206.615 182.535 206.945 182.915 ;
        RECT 207.125 182.705 207.385 183.210 ;
        RECT 207.555 182.705 207.815 184.915 ;
        RECT 207.985 184.705 208.315 185.085 ;
        RECT 208.485 184.745 209.770 184.915 ;
        RECT 208.485 184.285 208.655 184.745 ;
        RECT 209.440 184.705 209.770 184.745 ;
        RECT 209.940 184.585 210.150 184.915 ;
        RECT 208.005 184.115 208.655 184.285 ;
        RECT 208.955 184.435 209.285 184.575 ;
        RECT 208.955 184.205 209.740 184.435 ;
        RECT 208.005 183.335 208.175 184.115 ;
        RECT 208.485 183.555 208.940 183.725 ;
        RECT 208.750 183.375 209.160 183.385 ;
        RECT 208.005 183.165 208.575 183.335 ;
        RECT 208.065 182.535 208.235 182.995 ;
        RECT 208.405 182.875 208.575 183.165 ;
        RECT 208.745 183.215 209.160 183.375 ;
        RECT 208.745 183.045 208.920 183.215 ;
        RECT 209.570 183.035 209.740 184.205 ;
        RECT 209.980 183.385 210.150 184.585 ;
        RECT 210.445 184.585 210.630 184.915 ;
        RECT 210.800 184.705 211.150 185.085 ;
        RECT 210.445 183.725 210.615 184.585 ;
        RECT 211.400 184.535 211.570 184.915 ;
        RECT 211.740 184.705 212.070 185.085 ;
        RECT 212.295 184.745 213.305 184.915 ;
        RECT 212.295 184.535 212.465 184.745 ;
        RECT 211.400 184.365 212.465 184.535 ;
        RECT 210.325 183.555 210.615 183.725 ;
        RECT 209.910 183.215 210.150 183.385 ;
        RECT 210.445 183.105 210.615 183.555 ;
        RECT 210.785 183.445 211.075 184.125 ;
        RECT 211.550 183.505 211.880 184.125 ;
        RECT 212.085 184.065 212.330 184.125 ;
        RECT 212.635 184.065 212.965 184.575 ;
        RECT 213.135 184.235 213.305 184.745 ;
        RECT 213.565 184.705 213.895 185.085 ;
        RECT 212.085 183.895 212.385 184.065 ;
        RECT 212.635 183.895 213.395 184.065 ;
        RECT 212.085 183.505 212.330 183.895 ;
        RECT 212.670 183.715 212.840 183.725 ;
        RECT 212.670 183.555 213.055 183.715 ;
        RECT 212.725 183.545 213.055 183.555 ;
        RECT 212.740 183.335 212.910 183.375 ;
        RECT 213.225 183.370 213.395 183.895 ;
        RECT 213.565 183.445 213.865 184.445 ;
        RECT 214.065 184.075 214.415 184.915 ;
        RECT 214.585 184.745 216.115 184.915 ;
        RECT 214.585 184.245 214.755 184.745 ;
        RECT 215.945 184.585 216.115 184.745 ;
        RECT 216.285 184.705 216.615 185.085 ;
        RECT 214.925 184.405 215.255 184.575 ;
        RECT 215.085 184.075 215.255 184.405 ;
        RECT 215.425 184.415 215.595 184.575 ;
        RECT 216.785 184.415 216.955 184.915 ;
        RECT 215.425 184.245 216.955 184.415 ;
        RECT 214.065 183.845 214.870 184.075 ;
        RECT 215.085 183.905 215.720 184.075 ;
        RECT 214.510 183.735 214.870 183.845 ;
        RECT 214.510 183.555 215.050 183.735 ;
        RECT 211.390 183.165 212.910 183.335 ;
        RECT 209.230 182.875 209.400 183.035 ;
        RECT 208.405 182.705 209.400 182.875 ;
        RECT 209.570 182.865 210.100 183.035 ;
        RECT 209.930 182.705 210.100 182.865 ;
        RECT 210.445 182.775 210.620 183.105 ;
        RECT 210.790 182.535 211.120 182.915 ;
        RECT 211.390 182.745 211.635 183.165 ;
        RECT 212.740 183.045 212.910 183.165 ;
        RECT 213.080 183.295 213.395 183.370 ;
        RECT 213.080 183.045 213.410 183.295 ;
        RECT 211.810 182.535 211.980 182.995 ;
        RECT 212.150 182.875 212.505 182.915 ;
        RECT 213.580 182.875 213.750 183.245 ;
        RECT 212.150 182.705 213.750 182.875 ;
        RECT 214.040 182.535 214.330 183.255 ;
        RECT 214.510 182.880 214.870 183.555 ;
        RECT 215.550 183.385 215.720 183.905 ;
        RECT 215.890 183.445 216.325 184.065 ;
        RECT 216.635 183.895 216.985 184.065 ;
        RECT 217.215 184.010 217.485 184.915 ;
        RECT 217.655 184.325 217.985 185.085 ;
        RECT 218.165 184.155 218.335 184.915 ;
        RECT 216.635 183.445 216.980 183.895 ;
        RECT 215.430 183.215 215.720 183.385 ;
        RECT 215.040 182.875 215.210 183.210 ;
        RECT 215.380 183.045 215.720 183.215 ;
        RECT 215.945 183.085 216.955 183.255 ;
        RECT 215.945 182.875 216.115 183.085 ;
        RECT 215.040 182.705 216.115 182.875 ;
        RECT 216.285 182.535 216.615 182.915 ;
        RECT 216.785 182.710 216.955 183.085 ;
        RECT 217.215 183.210 217.385 184.010 ;
        RECT 217.670 183.985 218.335 184.155 ;
        RECT 218.685 184.155 218.855 184.915 ;
        RECT 219.035 184.325 219.365 185.085 ;
        RECT 218.685 183.985 219.350 184.155 ;
        RECT 219.535 184.010 219.805 184.915 ;
        RECT 220.065 184.415 220.235 184.915 ;
        RECT 220.405 184.705 220.735 185.085 ;
        RECT 220.905 184.745 222.435 184.915 ;
        RECT 220.905 184.585 221.075 184.745 ;
        RECT 221.425 184.415 221.595 184.575 ;
        RECT 220.065 184.245 221.595 184.415 ;
        RECT 221.765 184.405 222.095 184.575 ;
        RECT 221.765 184.075 221.935 184.405 ;
        RECT 222.265 184.245 222.435 184.745 ;
        RECT 222.605 184.075 222.955 184.915 ;
        RECT 223.125 184.705 223.455 185.085 ;
        RECT 223.715 184.745 224.725 184.915 ;
        RECT 217.670 183.840 217.840 183.985 ;
        RECT 217.555 183.510 217.840 183.840 ;
        RECT 219.180 183.840 219.350 183.985 ;
        RECT 217.670 183.255 217.840 183.510 ;
        RECT 218.075 183.435 218.405 183.805 ;
        RECT 218.615 183.435 218.945 183.805 ;
        RECT 219.180 183.510 219.465 183.840 ;
        RECT 219.180 183.255 219.350 183.510 ;
        RECT 217.215 182.705 217.475 183.210 ;
        RECT 217.670 183.085 218.335 183.255 ;
        RECT 217.655 182.535 217.985 182.915 ;
        RECT 218.165 182.705 218.335 183.085 ;
        RECT 218.685 183.085 219.350 183.255 ;
        RECT 219.635 183.210 219.805 184.010 ;
        RECT 220.040 183.725 220.385 184.065 ;
        RECT 220.035 183.555 220.385 183.725 ;
        RECT 220.040 183.445 220.385 183.555 ;
        RECT 220.695 183.445 221.130 184.065 ;
        RECT 221.300 183.905 221.935 184.075 ;
        RECT 221.300 183.385 221.470 183.905 ;
        RECT 222.150 183.845 222.955 184.075 ;
        RECT 222.150 183.735 222.510 183.845 ;
        RECT 221.970 183.555 222.510 183.735 ;
        RECT 218.685 182.705 218.855 183.085 ;
        RECT 219.035 182.535 219.365 182.915 ;
        RECT 219.545 182.705 219.805 183.210 ;
        RECT 220.065 183.085 221.075 183.255 ;
        RECT 220.065 182.710 220.235 183.085 ;
        RECT 220.405 182.535 220.735 182.915 ;
        RECT 220.905 182.875 221.075 183.085 ;
        RECT 221.300 183.215 221.590 183.385 ;
        RECT 221.300 183.045 221.640 183.215 ;
        RECT 221.810 182.875 221.980 183.210 ;
        RECT 222.150 182.880 222.510 183.555 ;
        RECT 223.155 183.445 223.455 184.445 ;
        RECT 223.715 184.235 223.885 184.745 ;
        RECT 224.055 184.065 224.385 184.575 ;
        RECT 224.555 184.535 224.725 184.745 ;
        RECT 224.950 184.705 225.280 185.085 ;
        RECT 225.450 184.535 225.620 184.915 ;
        RECT 225.870 184.705 226.220 185.085 ;
        RECT 226.390 184.585 226.575 184.915 ;
        RECT 224.555 184.365 225.620 184.535 ;
        RECT 224.690 184.065 224.935 184.125 ;
        RECT 223.625 183.895 224.385 184.065 ;
        RECT 224.635 183.895 224.935 184.065 ;
        RECT 223.625 183.370 223.795 183.895 ;
        RECT 224.180 183.715 224.350 183.725 ;
        RECT 223.965 183.555 224.350 183.715 ;
        RECT 223.965 183.545 224.295 183.555 ;
        RECT 224.690 183.505 224.935 183.895 ;
        RECT 225.140 184.065 225.470 184.125 ;
        RECT 225.140 183.895 225.495 184.065 ;
        RECT 225.140 183.505 225.470 183.895 ;
        RECT 225.945 183.445 226.235 184.125 ;
        RECT 226.405 183.725 226.575 184.585 ;
        RECT 226.870 184.585 227.080 184.915 ;
        RECT 227.250 184.745 228.535 184.915 ;
        RECT 227.250 184.705 227.580 184.745 ;
        RECT 226.405 183.555 226.695 183.725 ;
        RECT 223.625 183.295 223.940 183.370 ;
        RECT 220.905 182.705 221.980 182.875 ;
        RECT 222.690 182.535 222.980 183.255 ;
        RECT 223.270 182.875 223.440 183.245 ;
        RECT 223.610 183.045 223.940 183.295 ;
        RECT 224.110 183.335 224.280 183.375 ;
        RECT 224.110 183.165 225.630 183.335 ;
        RECT 224.110 183.045 224.280 183.165 ;
        RECT 224.515 182.875 224.870 182.915 ;
        RECT 223.270 182.705 224.870 182.875 ;
        RECT 225.040 182.535 225.210 182.995 ;
        RECT 225.385 182.745 225.630 183.165 ;
        RECT 226.405 183.105 226.575 183.555 ;
        RECT 226.870 183.385 227.040 184.585 ;
        RECT 227.735 184.435 228.065 184.575 ;
        RECT 227.280 184.205 228.065 184.435 ;
        RECT 228.365 184.285 228.535 184.745 ;
        RECT 228.705 184.705 229.035 185.085 ;
        RECT 226.870 183.215 227.110 183.385 ;
        RECT 225.900 182.535 226.230 182.915 ;
        RECT 226.400 182.775 226.575 183.105 ;
        RECT 227.280 183.035 227.450 184.205 ;
        RECT 228.365 184.115 229.015 184.285 ;
        RECT 228.080 183.555 228.535 183.725 ;
        RECT 227.860 183.375 228.270 183.385 ;
        RECT 227.860 183.215 228.275 183.375 ;
        RECT 228.845 183.335 229.015 184.115 ;
        RECT 228.100 183.045 228.275 183.215 ;
        RECT 228.445 183.165 229.015 183.335 ;
        RECT 226.920 182.865 227.450 183.035 ;
        RECT 227.620 182.875 227.790 183.035 ;
        RECT 228.445 182.875 228.615 183.165 ;
        RECT 226.920 182.705 227.090 182.865 ;
        RECT 227.620 182.705 228.615 182.875 ;
        RECT 228.785 182.535 228.955 182.995 ;
        RECT 229.205 182.705 229.465 184.915 ;
        RECT 229.635 183.920 229.925 185.085 ;
        RECT 230.185 184.155 230.355 184.915 ;
        RECT 230.535 184.325 230.865 185.085 ;
        RECT 230.185 183.985 230.850 184.155 ;
        RECT 231.035 184.010 231.305 184.915 ;
        RECT 230.680 183.840 230.850 183.985 ;
        RECT 230.115 183.435 230.445 183.805 ;
        RECT 230.680 183.510 230.965 183.840 ;
        RECT 229.635 182.535 229.925 183.260 ;
        RECT 230.680 183.255 230.850 183.510 ;
        RECT 230.185 183.085 230.850 183.255 ;
        RECT 231.135 183.210 231.305 184.010 ;
        RECT 230.185 182.705 230.355 183.085 ;
        RECT 230.535 182.535 230.865 182.915 ;
        RECT 231.045 182.705 231.305 183.210 ;
        RECT 231.475 184.010 231.745 184.915 ;
        RECT 231.915 184.325 232.245 185.085 ;
        RECT 232.425 184.155 232.595 184.915 ;
        RECT 231.475 183.210 231.645 184.010 ;
        RECT 231.930 183.985 232.595 184.155 ;
        RECT 232.855 184.010 233.125 184.915 ;
        RECT 233.295 184.325 233.625 185.085 ;
        RECT 233.805 184.155 233.975 184.915 ;
        RECT 231.930 183.840 232.100 183.985 ;
        RECT 231.815 183.510 232.100 183.840 ;
        RECT 231.930 183.255 232.100 183.510 ;
        RECT 232.335 183.435 232.665 183.805 ;
        RECT 231.475 182.705 231.735 183.210 ;
        RECT 231.930 183.085 232.595 183.255 ;
        RECT 231.915 182.535 232.245 182.915 ;
        RECT 232.425 182.705 232.595 183.085 ;
        RECT 232.855 183.210 233.025 184.010 ;
        RECT 233.310 183.985 233.975 184.155 ;
        RECT 234.235 184.010 234.505 184.915 ;
        RECT 234.675 184.325 235.005 185.085 ;
        RECT 235.185 184.155 235.355 184.915 ;
        RECT 233.310 183.840 233.480 183.985 ;
        RECT 233.195 183.510 233.480 183.840 ;
        RECT 233.310 183.255 233.480 183.510 ;
        RECT 233.715 183.435 234.045 183.805 ;
        RECT 232.855 182.705 233.115 183.210 ;
        RECT 233.310 183.085 233.975 183.255 ;
        RECT 233.295 182.535 233.625 182.915 ;
        RECT 233.805 182.705 233.975 183.085 ;
        RECT 234.235 183.210 234.405 184.010 ;
        RECT 234.690 183.985 235.355 184.155 ;
        RECT 235.615 184.010 235.885 184.915 ;
        RECT 236.055 184.325 236.385 185.085 ;
        RECT 236.565 184.155 236.735 184.915 ;
        RECT 234.690 183.840 234.860 183.985 ;
        RECT 234.575 183.510 234.860 183.840 ;
        RECT 234.690 183.255 234.860 183.510 ;
        RECT 235.095 183.435 235.425 183.805 ;
        RECT 234.235 182.705 234.495 183.210 ;
        RECT 234.690 183.085 235.355 183.255 ;
        RECT 234.675 182.535 235.005 182.915 ;
        RECT 235.185 182.705 235.355 183.085 ;
        RECT 235.615 183.210 235.785 184.010 ;
        RECT 236.070 183.985 236.735 184.155 ;
        RECT 237.915 183.995 239.125 185.085 ;
        RECT 236.070 183.840 236.240 183.985 ;
        RECT 235.955 183.510 236.240 183.840 ;
        RECT 236.070 183.255 236.240 183.510 ;
        RECT 236.475 183.435 236.805 183.805 ;
        RECT 237.915 183.455 238.435 183.995 ;
        RECT 238.605 183.285 239.125 183.825 ;
        RECT 235.615 182.705 235.875 183.210 ;
        RECT 236.070 183.085 236.735 183.255 ;
        RECT 236.055 182.535 236.385 182.915 ;
        RECT 236.565 182.705 236.735 183.085 ;
        RECT 237.915 182.535 239.125 183.285 ;
        RECT 165.150 182.365 239.210 182.535 ;
        RECT 165.235 181.615 166.445 182.365 ;
        RECT 166.615 181.865 166.875 182.195 ;
        RECT 167.085 181.885 167.360 182.365 ;
        RECT 165.235 181.075 165.755 181.615 ;
        RECT 102.225 180.620 155.700 181.020 ;
        RECT 165.925 180.905 166.445 181.445 ;
        RECT 62.895 180.305 99.045 180.475 ;
        RECT 9.330 178.450 52.060 178.620 ;
        RECT 9.330 168.690 9.500 178.450 ;
        RECT 10.230 177.760 12.230 177.930 ;
        RECT 12.520 177.760 14.520 177.930 ;
        RECT 14.810 177.760 16.810 177.930 ;
        RECT 17.100 177.760 19.100 177.930 ;
        RECT 19.390 177.760 21.390 177.930 ;
        RECT 21.680 177.760 23.680 177.930 ;
        RECT 23.970 177.760 25.970 177.930 ;
        RECT 26.260 177.760 28.260 177.930 ;
        RECT 28.550 177.760 30.550 177.930 ;
        RECT 30.840 177.760 32.840 177.930 ;
        RECT 33.130 177.760 35.130 177.930 ;
        RECT 35.420 177.760 37.420 177.930 ;
        RECT 37.710 177.760 39.710 177.930 ;
        RECT 40.000 177.760 42.000 177.930 ;
        RECT 42.290 177.760 44.290 177.930 ;
        RECT 44.580 177.760 46.580 177.930 ;
        RECT 46.870 177.760 48.870 177.930 ;
        RECT 49.160 177.760 51.160 177.930 ;
        RECT 10.000 169.550 10.170 177.590 ;
        RECT 12.290 169.550 12.460 177.590 ;
        RECT 14.580 169.550 14.750 177.590 ;
        RECT 16.870 169.550 17.040 177.590 ;
        RECT 19.160 169.550 19.330 177.590 ;
        RECT 21.450 169.550 21.620 177.590 ;
        RECT 23.740 169.550 23.910 177.590 ;
        RECT 26.030 169.550 26.200 177.590 ;
        RECT 28.320 169.550 28.490 177.590 ;
        RECT 30.610 169.550 30.780 177.590 ;
        RECT 32.900 169.550 33.070 177.590 ;
        RECT 35.190 169.550 35.360 177.590 ;
        RECT 37.480 169.550 37.650 177.590 ;
        RECT 39.770 169.550 39.940 177.590 ;
        RECT 42.060 169.550 42.230 177.590 ;
        RECT 44.350 169.550 44.520 177.590 ;
        RECT 46.640 169.550 46.810 177.590 ;
        RECT 48.930 169.550 49.100 177.590 ;
        RECT 51.220 169.550 51.390 177.590 ;
        RECT 10.230 169.210 12.230 169.380 ;
        RECT 12.520 169.210 14.520 169.380 ;
        RECT 14.810 169.210 16.810 169.380 ;
        RECT 17.100 169.210 19.100 169.380 ;
        RECT 19.390 169.210 21.390 169.380 ;
        RECT 21.680 169.210 23.680 169.380 ;
        RECT 23.970 169.210 25.970 169.380 ;
        RECT 26.260 169.210 28.260 169.380 ;
        RECT 28.550 169.210 30.550 169.380 ;
        RECT 30.840 169.210 32.840 169.380 ;
        RECT 33.130 169.210 35.130 169.380 ;
        RECT 35.420 169.210 37.420 169.380 ;
        RECT 37.710 169.210 39.710 169.380 ;
        RECT 40.000 169.210 42.000 169.380 ;
        RECT 42.290 169.210 44.290 169.380 ;
        RECT 44.580 169.210 46.580 169.380 ;
        RECT 46.870 169.210 48.870 169.380 ;
        RECT 49.160 169.210 51.160 169.380 ;
        RECT 51.890 168.690 52.060 178.450 ;
        RECT 62.895 177.455 63.425 180.305 ;
        RECT 64.155 179.615 80.155 179.785 ;
        RECT 63.925 178.360 64.095 179.400 ;
        RECT 80.215 178.360 80.385 179.400 ;
        RECT 64.155 177.975 80.155 178.145 ;
        RECT 80.885 177.455 81.055 180.305 ;
        RECT 81.785 179.615 97.785 179.785 ;
        RECT 81.555 178.360 81.725 179.400 ;
        RECT 97.845 178.360 98.015 179.400 ;
        RECT 81.785 177.975 97.785 178.145 ;
        RECT 98.515 177.455 99.045 180.305 ;
        RECT 62.895 177.285 99.045 177.455 ;
        RECT 62.895 174.435 63.425 177.285 ;
        RECT 64.155 176.595 80.155 176.765 ;
        RECT 63.925 175.340 64.095 176.380 ;
        RECT 80.215 175.340 80.385 176.380 ;
        RECT 64.155 174.955 80.155 175.125 ;
        RECT 80.885 174.435 81.055 177.285 ;
        RECT 81.785 176.595 97.785 176.765 ;
        RECT 81.555 175.340 81.725 176.380 ;
        RECT 97.845 175.340 98.015 176.380 ;
        RECT 81.785 174.955 97.785 175.125 ;
        RECT 98.515 174.435 99.045 177.285 ;
        RECT 62.895 174.265 99.045 174.435 ;
        RECT 62.895 171.415 63.425 174.265 ;
        RECT 63.925 173.575 80.385 173.745 ;
        RECT 63.925 172.105 64.155 173.575 ;
        RECT 80.155 172.105 80.385 173.575 ;
        RECT 63.925 171.935 80.385 172.105 ;
        RECT 80.885 171.415 81.055 174.265 ;
        RECT 81.555 173.575 98.015 173.745 ;
        RECT 81.555 172.105 81.785 173.575 ;
        RECT 97.785 172.105 98.015 173.575 ;
        RECT 81.555 171.935 98.015 172.105 ;
        RECT 98.515 171.415 99.045 174.265 ;
        RECT 113.860 176.355 151.710 176.885 ;
        RECT 62.895 170.885 99.045 171.415 ;
        RECT 102.740 172.330 110.970 172.500 ;
        RECT 9.330 168.520 52.060 168.690 ;
        RECT 9.330 167.860 51.780 168.030 ;
        RECT 9.330 158.100 9.500 167.860 ;
        RECT 10.290 167.170 12.290 167.340 ;
        RECT 12.580 167.170 14.580 167.340 ;
        RECT 10.060 158.960 10.230 167.000 ;
        RECT 12.350 158.960 12.520 167.000 ;
        RECT 14.640 158.960 14.810 167.000 ;
        RECT 10.290 158.620 12.290 158.790 ;
        RECT 12.580 158.620 14.580 158.790 ;
        RECT 15.370 158.100 15.540 167.860 ;
        RECT 16.330 167.170 18.330 167.340 ;
        RECT 18.620 167.170 20.620 167.340 ;
        RECT 16.100 158.960 16.270 167.000 ;
        RECT 18.390 158.960 18.560 167.000 ;
        RECT 20.680 158.960 20.850 167.000 ;
        RECT 16.330 158.620 18.330 158.790 ;
        RECT 18.620 158.620 20.620 158.790 ;
        RECT 21.410 158.100 21.580 167.860 ;
        RECT 22.370 167.170 24.370 167.340 ;
        RECT 24.660 167.170 26.660 167.340 ;
        RECT 22.140 158.960 22.310 167.000 ;
        RECT 24.430 158.960 24.600 167.000 ;
        RECT 26.720 158.960 26.890 167.000 ;
        RECT 22.370 158.620 24.370 158.790 ;
        RECT 24.660 158.620 26.660 158.790 ;
        RECT 27.450 158.100 27.620 167.860 ;
        RECT 28.410 167.170 30.410 167.340 ;
        RECT 30.700 167.170 32.700 167.340 ;
        RECT 28.180 158.960 28.350 167.000 ;
        RECT 30.470 158.960 30.640 167.000 ;
        RECT 32.760 158.960 32.930 167.000 ;
        RECT 28.410 158.620 30.410 158.790 ;
        RECT 30.700 158.620 32.700 158.790 ;
        RECT 33.490 158.100 33.660 167.860 ;
        RECT 34.450 167.170 36.450 167.340 ;
        RECT 36.740 167.170 38.740 167.340 ;
        RECT 34.220 158.960 34.390 167.000 ;
        RECT 36.510 158.960 36.680 167.000 ;
        RECT 38.800 158.960 38.970 167.000 ;
        RECT 34.450 158.620 36.450 158.790 ;
        RECT 36.740 158.620 38.740 158.790 ;
        RECT 39.530 158.100 39.700 167.860 ;
        RECT 40.490 167.170 42.490 167.340 ;
        RECT 42.780 167.170 44.780 167.340 ;
        RECT 40.260 158.960 40.430 167.000 ;
        RECT 42.550 158.960 42.720 167.000 ;
        RECT 44.840 158.960 45.010 167.000 ;
        RECT 40.490 158.620 42.490 158.790 ;
        RECT 42.780 158.620 44.780 158.790 ;
        RECT 45.570 158.100 45.740 167.860 ;
        RECT 46.530 167.170 48.530 167.340 ;
        RECT 48.820 167.170 50.820 167.340 ;
        RECT 46.300 158.960 46.470 167.000 ;
        RECT 48.590 158.960 48.760 167.000 ;
        RECT 50.880 158.960 51.050 167.000 ;
        RECT 46.530 158.620 48.530 158.790 ;
        RECT 48.820 158.620 50.820 158.790 ;
        RECT 51.610 158.100 51.780 167.860 ;
        RECT 9.330 157.930 51.780 158.100 ;
        RECT 9.330 148.170 9.500 157.930 ;
        RECT 10.290 157.240 12.290 157.410 ;
        RECT 12.580 157.240 14.580 157.410 ;
        RECT 10.060 149.030 10.230 157.070 ;
        RECT 12.350 149.030 12.520 157.070 ;
        RECT 14.640 149.030 14.810 157.070 ;
        RECT 10.290 148.690 12.290 148.860 ;
        RECT 12.580 148.690 14.580 148.860 ;
        RECT 15.370 148.170 15.540 157.930 ;
        RECT 16.330 157.240 18.330 157.410 ;
        RECT 18.620 157.240 20.620 157.410 ;
        RECT 16.100 149.030 16.270 157.070 ;
        RECT 18.390 149.030 18.560 157.070 ;
        RECT 20.680 149.030 20.850 157.070 ;
        RECT 16.330 148.690 18.330 148.860 ;
        RECT 18.620 148.690 20.620 148.860 ;
        RECT 21.410 148.170 21.580 157.930 ;
        RECT 22.370 157.240 24.370 157.410 ;
        RECT 24.660 157.240 26.660 157.410 ;
        RECT 22.140 149.030 22.310 157.070 ;
        RECT 24.430 149.030 24.600 157.070 ;
        RECT 26.720 149.030 26.890 157.070 ;
        RECT 22.370 148.690 24.370 148.860 ;
        RECT 24.660 148.690 26.660 148.860 ;
        RECT 27.450 148.170 27.620 157.930 ;
        RECT 28.410 157.240 30.410 157.410 ;
        RECT 30.700 157.240 32.700 157.410 ;
        RECT 28.180 149.030 28.350 157.070 ;
        RECT 30.470 149.030 30.640 157.070 ;
        RECT 32.760 149.030 32.930 157.070 ;
        RECT 28.410 148.690 30.410 148.860 ;
        RECT 30.700 148.690 32.700 148.860 ;
        RECT 33.490 148.170 33.660 157.930 ;
        RECT 34.450 157.240 36.450 157.410 ;
        RECT 36.740 157.240 38.740 157.410 ;
        RECT 34.220 149.030 34.390 157.070 ;
        RECT 36.510 149.030 36.680 157.070 ;
        RECT 38.800 149.030 38.970 157.070 ;
        RECT 34.450 148.690 36.450 148.860 ;
        RECT 36.740 148.690 38.740 148.860 ;
        RECT 39.530 148.170 39.700 157.930 ;
        RECT 40.490 157.240 42.490 157.410 ;
        RECT 42.780 157.240 44.780 157.410 ;
        RECT 40.260 149.030 40.430 157.070 ;
        RECT 42.550 149.030 42.720 157.070 ;
        RECT 44.840 149.030 45.010 157.070 ;
        RECT 40.490 148.690 42.490 148.860 ;
        RECT 42.780 148.690 44.780 148.860 ;
        RECT 45.570 148.170 45.740 157.930 ;
        RECT 46.530 157.240 48.530 157.410 ;
        RECT 48.820 157.240 50.820 157.410 ;
        RECT 46.300 149.030 46.470 157.070 ;
        RECT 48.590 149.030 48.760 157.070 ;
        RECT 50.880 149.030 51.050 157.070 ;
        RECT 46.530 148.690 48.530 148.860 ;
        RECT 48.820 148.690 50.820 148.860 ;
        RECT 51.610 148.170 51.780 157.930 ;
        RECT 9.330 148.000 51.780 148.170 ;
        RECT 64.100 166.025 96.940 166.425 ;
        RECT 23.195 143.155 58.705 143.745 ;
        RECT 23.195 140.745 23.785 143.155 ;
        RECT 24.515 142.465 32.515 142.635 ;
        RECT 32.805 142.465 40.805 142.635 ;
        RECT 41.095 142.465 49.095 142.635 ;
        RECT 49.385 142.465 57.385 142.635 ;
        RECT 24.285 141.255 24.455 142.295 ;
        RECT 32.575 141.255 32.745 142.295 ;
        RECT 40.865 141.255 41.035 142.295 ;
        RECT 49.155 141.255 49.325 142.295 ;
        RECT 57.445 141.255 57.615 142.295 ;
        RECT 24.515 140.915 32.515 141.085 ;
        RECT 32.805 140.915 40.805 141.085 ;
        RECT 41.095 140.915 49.095 141.085 ;
        RECT 49.385 140.915 57.385 141.085 ;
        RECT 23.195 139.705 24.455 140.745 ;
        RECT 32.575 139.705 32.745 140.745 ;
        RECT 40.865 139.705 41.035 140.745 ;
        RECT 49.155 139.705 49.325 140.745 ;
        RECT 57.445 139.705 57.615 140.745 ;
        RECT 23.195 139.195 23.785 139.705 ;
        RECT 24.515 139.365 32.515 139.535 ;
        RECT 32.805 139.365 40.805 139.535 ;
        RECT 41.095 139.365 49.095 139.535 ;
        RECT 49.385 139.365 57.385 139.535 ;
        RECT 9.430 137.955 20.720 138.485 ;
        RECT 9.430 135.195 9.960 137.955 ;
        RECT 10.995 137.265 11.995 137.435 ;
        RECT 10.765 136.055 10.935 137.095 ;
        RECT 12.055 136.055 12.225 137.095 ;
        RECT 13.030 135.195 13.200 137.955 ;
        RECT 13.930 137.265 14.930 137.435 ;
        RECT 15.220 137.265 16.220 137.435 ;
        RECT 13.700 136.055 13.870 137.095 ;
        RECT 14.990 136.055 15.160 137.095 ;
        RECT 16.280 136.055 16.450 137.095 ;
        RECT 16.950 135.195 17.120 137.955 ;
        RECT 18.155 137.265 19.155 137.435 ;
        RECT 17.925 136.055 18.095 137.095 ;
        RECT 19.215 136.055 19.385 137.095 ;
        RECT 20.190 135.195 20.720 137.955 ;
        RECT 9.430 134.665 20.720 135.195 ;
        RECT 23.195 138.155 24.455 139.195 ;
        RECT 32.575 138.155 32.745 139.195 ;
        RECT 40.865 138.155 41.035 139.195 ;
        RECT 49.155 138.155 49.325 139.195 ;
        RECT 57.445 138.155 57.615 139.195 ;
        RECT 23.195 135.745 23.785 138.155 ;
        RECT 24.515 137.815 32.515 137.985 ;
        RECT 32.805 137.815 40.805 137.985 ;
        RECT 41.095 137.815 49.095 137.985 ;
        RECT 49.385 137.815 57.385 137.985 ;
        RECT 24.285 136.605 24.455 137.645 ;
        RECT 32.575 136.605 32.745 137.645 ;
        RECT 40.865 136.605 41.035 137.645 ;
        RECT 49.155 136.605 49.325 137.645 ;
        RECT 57.445 136.605 57.615 137.645 ;
        RECT 24.515 136.265 32.515 136.435 ;
        RECT 32.805 136.265 40.805 136.435 ;
        RECT 41.095 136.265 49.095 136.435 ;
        RECT 49.385 136.265 57.385 136.435 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 23.195 135.155 58.705 135.745 ;
        RECT 64.100 133.985 64.500 166.025 ;
        RECT 69.635 160.720 91.405 160.890 ;
        RECT 69.635 139.290 69.805 160.720 ;
        RECT 71.220 158.800 89.820 159.305 ;
        RECT 71.220 156.090 71.725 158.800 ;
        RECT 72.035 158.130 74.125 158.490 ;
        RECT 72.035 156.760 72.395 158.130 ;
        RECT 72.685 157.050 73.475 157.840 ;
        RECT 73.765 156.760 74.125 158.130 ;
        RECT 72.035 156.400 74.125 156.760 ;
        RECT 74.435 156.090 75.445 158.800 ;
        RECT 75.755 158.130 77.845 158.490 ;
        RECT 75.755 156.760 76.115 158.130 ;
        RECT 76.405 157.050 77.195 157.840 ;
        RECT 77.485 156.760 77.845 158.130 ;
        RECT 75.755 156.400 77.845 156.760 ;
        RECT 78.155 156.090 79.165 158.800 ;
        RECT 79.475 158.130 81.565 158.490 ;
        RECT 79.475 156.760 79.835 158.130 ;
        RECT 80.125 157.050 80.915 157.840 ;
        RECT 81.205 156.760 81.565 158.130 ;
        RECT 79.475 156.400 81.565 156.760 ;
        RECT 81.875 156.090 82.885 158.800 ;
        RECT 83.195 158.130 85.285 158.490 ;
        RECT 83.195 156.760 83.555 158.130 ;
        RECT 83.845 157.050 84.635 157.840 ;
        RECT 84.925 156.760 85.285 158.130 ;
        RECT 83.195 156.400 85.285 156.760 ;
        RECT 85.595 156.090 86.605 158.800 ;
        RECT 86.915 158.130 89.005 158.490 ;
        RECT 86.915 156.760 87.275 158.130 ;
        RECT 87.565 157.050 88.355 157.840 ;
        RECT 88.645 156.760 89.005 158.130 ;
        RECT 86.915 156.400 89.005 156.760 ;
        RECT 89.315 156.090 89.820 158.800 ;
        RECT 71.220 155.080 89.820 156.090 ;
        RECT 71.220 152.370 71.725 155.080 ;
        RECT 72.035 154.410 74.125 154.770 ;
        RECT 72.035 153.040 72.395 154.410 ;
        RECT 72.685 153.330 73.475 154.120 ;
        RECT 73.765 153.040 74.125 154.410 ;
        RECT 72.035 152.680 74.125 153.040 ;
        RECT 74.435 152.370 75.445 155.080 ;
        RECT 75.755 154.410 77.845 154.770 ;
        RECT 75.755 153.040 76.115 154.410 ;
        RECT 76.405 153.330 77.195 154.120 ;
        RECT 77.485 153.040 77.845 154.410 ;
        RECT 75.755 152.680 77.845 153.040 ;
        RECT 78.155 152.370 79.165 155.080 ;
        RECT 79.475 154.410 81.565 154.770 ;
        RECT 79.475 153.040 79.835 154.410 ;
        RECT 80.125 153.330 80.915 154.120 ;
        RECT 81.205 153.040 81.565 154.410 ;
        RECT 79.475 152.680 81.565 153.040 ;
        RECT 81.875 152.370 82.885 155.080 ;
        RECT 83.195 154.410 85.285 154.770 ;
        RECT 83.195 153.040 83.555 154.410 ;
        RECT 83.845 153.330 84.635 154.120 ;
        RECT 84.925 153.040 85.285 154.410 ;
        RECT 83.195 152.680 85.285 153.040 ;
        RECT 85.595 152.370 86.605 155.080 ;
        RECT 86.915 154.410 89.005 154.770 ;
        RECT 86.915 153.040 87.275 154.410 ;
        RECT 87.565 153.330 88.355 154.120 ;
        RECT 88.645 153.040 89.005 154.410 ;
        RECT 86.915 152.680 89.005 153.040 ;
        RECT 89.315 152.370 89.820 155.080 ;
        RECT 71.220 151.360 89.820 152.370 ;
        RECT 71.220 148.650 71.725 151.360 ;
        RECT 72.035 150.690 74.125 151.050 ;
        RECT 72.035 149.320 72.395 150.690 ;
        RECT 72.685 149.610 73.475 150.400 ;
        RECT 73.765 149.320 74.125 150.690 ;
        RECT 72.035 148.960 74.125 149.320 ;
        RECT 74.435 148.650 75.445 151.360 ;
        RECT 75.755 150.690 77.845 151.050 ;
        RECT 75.755 149.320 76.115 150.690 ;
        RECT 76.405 149.610 77.195 150.400 ;
        RECT 77.485 149.320 77.845 150.690 ;
        RECT 75.755 148.960 77.845 149.320 ;
        RECT 78.155 148.650 79.165 151.360 ;
        RECT 79.475 150.690 81.565 151.050 ;
        RECT 79.475 149.320 79.835 150.690 ;
        RECT 80.125 149.610 80.915 150.400 ;
        RECT 81.205 149.320 81.565 150.690 ;
        RECT 79.475 148.960 81.565 149.320 ;
        RECT 81.875 148.650 82.885 151.360 ;
        RECT 83.195 150.690 85.285 151.050 ;
        RECT 83.195 149.320 83.555 150.690 ;
        RECT 83.845 149.610 84.635 150.400 ;
        RECT 84.925 149.320 85.285 150.690 ;
        RECT 83.195 148.960 85.285 149.320 ;
        RECT 85.595 148.650 86.605 151.360 ;
        RECT 86.915 150.690 89.005 151.050 ;
        RECT 86.915 149.320 87.275 150.690 ;
        RECT 87.565 149.610 88.355 150.400 ;
        RECT 88.645 149.320 89.005 150.690 ;
        RECT 86.915 148.960 89.005 149.320 ;
        RECT 89.315 148.650 89.820 151.360 ;
        RECT 71.220 147.640 89.820 148.650 ;
        RECT 71.220 144.930 71.725 147.640 ;
        RECT 72.035 146.970 74.125 147.330 ;
        RECT 72.035 145.600 72.395 146.970 ;
        RECT 72.685 145.890 73.475 146.680 ;
        RECT 73.765 145.600 74.125 146.970 ;
        RECT 72.035 145.240 74.125 145.600 ;
        RECT 74.435 144.930 75.445 147.640 ;
        RECT 75.755 146.970 77.845 147.330 ;
        RECT 75.755 145.600 76.115 146.970 ;
        RECT 76.405 145.890 77.195 146.680 ;
        RECT 77.485 145.600 77.845 146.970 ;
        RECT 75.755 145.240 77.845 145.600 ;
        RECT 78.155 144.930 79.165 147.640 ;
        RECT 79.475 146.970 81.565 147.330 ;
        RECT 79.475 145.600 79.835 146.970 ;
        RECT 80.125 145.890 80.915 146.680 ;
        RECT 81.205 145.600 81.565 146.970 ;
        RECT 79.475 145.240 81.565 145.600 ;
        RECT 81.875 144.930 82.885 147.640 ;
        RECT 83.195 146.970 85.285 147.330 ;
        RECT 83.195 145.600 83.555 146.970 ;
        RECT 83.845 145.890 84.635 146.680 ;
        RECT 84.925 145.600 85.285 146.970 ;
        RECT 83.195 145.240 85.285 145.600 ;
        RECT 85.595 144.930 86.605 147.640 ;
        RECT 86.915 146.970 89.005 147.330 ;
        RECT 86.915 145.600 87.275 146.970 ;
        RECT 87.565 145.890 88.355 146.680 ;
        RECT 88.645 145.600 89.005 146.970 ;
        RECT 86.915 145.240 89.005 145.600 ;
        RECT 89.315 144.930 89.820 147.640 ;
        RECT 71.220 143.920 89.820 144.930 ;
        RECT 71.220 141.210 71.725 143.920 ;
        RECT 72.035 143.250 74.125 143.610 ;
        RECT 72.035 141.880 72.395 143.250 ;
        RECT 72.685 142.170 73.475 142.960 ;
        RECT 73.765 141.880 74.125 143.250 ;
        RECT 72.035 141.520 74.125 141.880 ;
        RECT 74.435 141.210 75.445 143.920 ;
        RECT 75.755 143.250 77.845 143.610 ;
        RECT 75.755 141.880 76.115 143.250 ;
        RECT 76.405 142.170 77.195 142.960 ;
        RECT 77.485 141.880 77.845 143.250 ;
        RECT 75.755 141.520 77.845 141.880 ;
        RECT 78.155 141.210 79.165 143.920 ;
        RECT 79.475 143.250 81.565 143.610 ;
        RECT 79.475 141.880 79.835 143.250 ;
        RECT 80.125 142.170 80.915 142.960 ;
        RECT 81.205 141.880 81.565 143.250 ;
        RECT 79.475 141.520 81.565 141.880 ;
        RECT 81.875 141.210 82.885 143.920 ;
        RECT 83.195 143.250 85.285 143.610 ;
        RECT 83.195 141.880 83.555 143.250 ;
        RECT 83.845 142.170 84.635 142.960 ;
        RECT 84.925 141.880 85.285 143.250 ;
        RECT 83.195 141.520 85.285 141.880 ;
        RECT 85.595 141.210 86.605 143.920 ;
        RECT 86.915 143.250 89.005 143.610 ;
        RECT 86.915 141.880 87.275 143.250 ;
        RECT 87.565 142.170 88.355 142.960 ;
        RECT 88.645 141.880 89.005 143.250 ;
        RECT 86.915 141.520 89.005 141.880 ;
        RECT 89.315 141.210 89.820 143.920 ;
        RECT 71.220 140.705 89.820 141.210 ;
        RECT 91.235 139.290 91.405 160.720 ;
        RECT 69.635 139.120 91.405 139.290 ;
        RECT 96.540 133.985 96.940 166.025 ;
        RECT 102.740 162.570 102.910 172.330 ;
        RECT 103.695 171.640 104.695 171.810 ;
        RECT 104.985 171.640 105.985 171.810 ;
        RECT 103.465 163.430 103.635 171.470 ;
        RECT 104.755 163.430 104.925 171.470 ;
        RECT 106.045 163.430 106.215 171.470 ;
        RECT 103.695 163.090 104.695 163.260 ;
        RECT 104.985 163.090 105.985 163.260 ;
        RECT 106.770 162.570 106.940 172.330 ;
        RECT 107.725 171.640 108.725 171.810 ;
        RECT 109.015 171.640 110.015 171.810 ;
        RECT 107.495 163.430 107.665 171.470 ;
        RECT 108.785 163.430 108.955 171.470 ;
        RECT 110.075 163.430 110.245 171.470 ;
        RECT 107.725 163.090 108.725 163.260 ;
        RECT 109.015 163.090 110.015 163.260 ;
        RECT 110.800 162.570 110.970 172.330 ;
        RECT 113.860 166.595 114.390 176.355 ;
        RECT 115.180 175.665 115.680 175.835 ;
        RECT 115.970 175.665 116.470 175.835 ;
        RECT 116.760 175.665 117.260 175.835 ;
        RECT 117.550 175.665 118.050 175.835 ;
        RECT 114.950 167.455 115.120 175.495 ;
        RECT 115.740 167.455 115.910 175.495 ;
        RECT 116.530 167.455 116.700 175.495 ;
        RECT 117.320 167.455 117.490 175.495 ;
        RECT 118.110 167.455 118.280 175.495 ;
        RECT 115.180 167.115 115.680 167.285 ;
        RECT 115.970 167.115 116.470 167.285 ;
        RECT 116.760 167.115 117.260 167.285 ;
        RECT 117.550 167.115 118.050 167.285 ;
        RECT 118.840 166.595 119.010 176.355 ;
        RECT 119.800 175.665 120.300 175.835 ;
        RECT 120.590 175.665 121.090 175.835 ;
        RECT 121.380 175.665 121.880 175.835 ;
        RECT 122.170 175.665 122.670 175.835 ;
        RECT 119.570 167.455 119.740 175.495 ;
        RECT 120.360 167.455 120.530 175.495 ;
        RECT 121.150 167.455 121.320 175.495 ;
        RECT 121.940 167.455 122.110 175.495 ;
        RECT 122.730 167.455 122.900 175.495 ;
        RECT 119.800 167.115 120.300 167.285 ;
        RECT 120.590 167.115 121.090 167.285 ;
        RECT 121.380 167.115 121.880 167.285 ;
        RECT 122.170 167.115 122.670 167.285 ;
        RECT 123.460 166.595 123.630 176.355 ;
        RECT 124.420 175.665 124.920 175.835 ;
        RECT 125.210 175.665 125.710 175.835 ;
        RECT 126.000 175.665 126.500 175.835 ;
        RECT 126.790 175.665 127.290 175.835 ;
        RECT 124.190 167.455 124.360 175.495 ;
        RECT 124.980 167.455 125.150 175.495 ;
        RECT 125.770 167.455 125.940 175.495 ;
        RECT 126.560 167.455 126.730 175.495 ;
        RECT 127.350 167.455 127.520 175.495 ;
        RECT 124.420 167.115 124.920 167.285 ;
        RECT 125.210 167.115 125.710 167.285 ;
        RECT 126.000 167.115 126.500 167.285 ;
        RECT 126.790 167.115 127.290 167.285 ;
        RECT 128.080 166.595 128.250 176.355 ;
        RECT 129.040 175.665 129.540 175.835 ;
        RECT 129.830 175.665 130.330 175.835 ;
        RECT 130.620 175.665 131.120 175.835 ;
        RECT 131.410 175.665 131.910 175.835 ;
        RECT 128.810 167.455 128.980 175.495 ;
        RECT 129.600 167.455 129.770 175.495 ;
        RECT 130.390 167.455 130.560 175.495 ;
        RECT 131.180 167.455 131.350 175.495 ;
        RECT 131.970 167.455 132.140 175.495 ;
        RECT 129.040 167.115 129.540 167.285 ;
        RECT 129.830 167.115 130.330 167.285 ;
        RECT 130.620 167.115 131.120 167.285 ;
        RECT 131.410 167.115 131.910 167.285 ;
        RECT 132.700 166.595 132.870 176.355 ;
        RECT 133.660 175.665 134.160 175.835 ;
        RECT 134.450 175.665 134.950 175.835 ;
        RECT 135.240 175.665 135.740 175.835 ;
        RECT 136.030 175.665 136.530 175.835 ;
        RECT 133.430 167.455 133.600 175.495 ;
        RECT 134.220 167.455 134.390 175.495 ;
        RECT 135.010 167.455 135.180 175.495 ;
        RECT 135.800 167.455 135.970 175.495 ;
        RECT 136.590 167.455 136.760 175.495 ;
        RECT 133.660 167.115 134.160 167.285 ;
        RECT 134.450 167.115 134.950 167.285 ;
        RECT 135.240 167.115 135.740 167.285 ;
        RECT 136.030 167.115 136.530 167.285 ;
        RECT 137.320 166.595 137.490 176.355 ;
        RECT 138.280 175.665 138.780 175.835 ;
        RECT 139.070 175.665 139.570 175.835 ;
        RECT 139.860 175.665 140.360 175.835 ;
        RECT 140.650 175.665 141.150 175.835 ;
        RECT 138.050 167.455 138.220 175.495 ;
        RECT 138.840 167.455 139.010 175.495 ;
        RECT 139.630 167.455 139.800 175.495 ;
        RECT 140.420 167.455 140.590 175.495 ;
        RECT 141.210 167.455 141.380 175.495 ;
        RECT 138.280 167.115 138.780 167.285 ;
        RECT 139.070 167.115 139.570 167.285 ;
        RECT 139.860 167.115 140.360 167.285 ;
        RECT 140.650 167.115 141.150 167.285 ;
        RECT 141.940 166.595 142.110 176.355 ;
        RECT 142.900 175.665 143.400 175.835 ;
        RECT 143.690 175.665 144.190 175.835 ;
        RECT 144.480 175.665 144.980 175.835 ;
        RECT 145.270 175.665 145.770 175.835 ;
        RECT 142.670 167.455 142.840 175.495 ;
        RECT 143.460 167.455 143.630 175.495 ;
        RECT 144.250 167.455 144.420 175.495 ;
        RECT 145.040 167.455 145.210 175.495 ;
        RECT 145.830 167.455 146.000 175.495 ;
        RECT 142.900 167.115 143.400 167.285 ;
        RECT 143.690 167.115 144.190 167.285 ;
        RECT 144.480 167.115 144.980 167.285 ;
        RECT 145.270 167.115 145.770 167.285 ;
        RECT 146.560 166.595 146.730 176.355 ;
        RECT 147.520 175.665 148.020 175.835 ;
        RECT 148.310 175.665 148.810 175.835 ;
        RECT 149.100 175.665 149.600 175.835 ;
        RECT 149.890 175.665 150.390 175.835 ;
        RECT 147.290 167.455 147.460 175.495 ;
        RECT 148.080 167.455 148.250 175.495 ;
        RECT 148.870 167.455 149.040 175.495 ;
        RECT 149.660 167.455 149.830 175.495 ;
        RECT 150.450 167.455 150.620 175.495 ;
        RECT 147.520 167.115 148.020 167.285 ;
        RECT 148.310 167.115 148.810 167.285 ;
        RECT 149.100 167.115 149.600 167.285 ;
        RECT 149.890 167.115 150.390 167.285 ;
        RECT 151.180 166.595 151.710 176.355 ;
        RECT 113.860 166.065 151.710 166.595 ;
        RECT 102.740 162.400 110.970 162.570 ;
        RECT 102.740 158.640 102.910 162.400 ;
        RECT 103.465 159.500 103.635 161.540 ;
        RECT 104.755 159.500 104.925 161.540 ;
        RECT 106.045 159.500 106.215 161.540 ;
        RECT 103.695 159.160 104.695 159.330 ;
        RECT 104.985 159.160 105.985 159.330 ;
        RECT 106.770 158.640 106.940 162.400 ;
        RECT 107.495 159.500 107.665 161.540 ;
        RECT 108.785 159.500 108.955 161.540 ;
        RECT 110.075 159.500 110.245 161.540 ;
        RECT 107.725 159.160 108.725 159.330 ;
        RECT 109.015 159.160 110.015 159.330 ;
        RECT 110.800 158.640 110.970 162.400 ;
        RECT 102.740 158.470 110.970 158.640 ;
        RECT 116.015 157.500 149.445 158.030 ;
        RECT 102.740 155.775 110.970 155.945 ;
        RECT 102.740 151.925 102.910 155.775 ;
        RECT 103.695 155.085 104.695 155.255 ;
        RECT 104.985 155.085 105.985 155.255 ;
        RECT 103.465 152.830 103.635 154.870 ;
        RECT 104.755 152.830 104.925 154.870 ;
        RECT 106.045 152.830 106.215 154.870 ;
        RECT 106.770 151.925 106.940 155.775 ;
        RECT 107.725 155.085 108.725 155.255 ;
        RECT 109.015 155.085 110.015 155.255 ;
        RECT 107.495 152.830 107.665 154.870 ;
        RECT 108.785 152.830 108.955 154.870 ;
        RECT 110.075 152.830 110.245 154.870 ;
        RECT 110.800 151.925 110.970 155.775 ;
        RECT 102.740 151.755 110.970 151.925 ;
        RECT 102.740 141.905 102.910 151.755 ;
        RECT 103.695 151.065 104.695 151.235 ;
        RECT 104.985 151.065 105.985 151.235 ;
        RECT 103.465 142.810 103.635 150.850 ;
        RECT 104.755 142.810 104.925 150.850 ;
        RECT 106.045 142.810 106.215 150.850 ;
        RECT 103.695 142.425 104.695 142.595 ;
        RECT 104.985 142.425 105.985 142.595 ;
        RECT 106.770 141.905 106.940 151.755 ;
        RECT 107.725 151.065 108.725 151.235 ;
        RECT 109.015 151.065 110.015 151.235 ;
        RECT 107.495 142.810 107.665 150.850 ;
        RECT 108.785 142.810 108.955 150.850 ;
        RECT 110.075 142.810 110.245 150.850 ;
        RECT 107.725 142.425 108.725 142.595 ;
        RECT 109.015 142.425 110.015 142.595 ;
        RECT 110.800 141.905 110.970 151.755 ;
        RECT 102.740 141.735 110.970 141.905 ;
        RECT 116.015 140.250 116.545 157.500 ;
        RECT 117.130 156.135 119.290 156.825 ;
        RECT 117.130 154.965 119.290 155.655 ;
        RECT 117.130 153.795 119.290 154.485 ;
        RECT 117.130 152.625 119.290 153.315 ;
        RECT 117.130 151.455 119.290 152.145 ;
        RECT 117.130 150.285 119.290 150.975 ;
        RECT 117.130 149.115 119.290 149.805 ;
        RECT 117.130 147.945 119.290 148.635 ;
        RECT 117.130 146.775 119.290 147.465 ;
        RECT 117.130 145.605 119.290 146.295 ;
        RECT 117.130 144.435 119.290 145.125 ;
        RECT 117.130 143.265 119.290 143.955 ;
        RECT 117.130 142.095 119.290 142.785 ;
        RECT 117.130 140.925 119.290 141.615 ;
        RECT 119.595 140.250 122.075 157.500 ;
        RECT 122.380 156.135 124.540 156.825 ;
        RECT 125.060 156.135 127.220 156.825 ;
        RECT 122.380 154.965 124.540 155.655 ;
        RECT 125.060 154.965 127.220 155.655 ;
        RECT 122.380 153.795 124.540 154.485 ;
        RECT 125.060 153.795 127.220 154.485 ;
        RECT 122.380 152.625 124.540 153.315 ;
        RECT 125.060 152.625 127.220 153.315 ;
        RECT 122.380 151.455 124.540 152.145 ;
        RECT 125.060 151.455 127.220 152.145 ;
        RECT 122.380 150.285 124.540 150.975 ;
        RECT 125.060 150.285 127.220 150.975 ;
        RECT 122.380 149.115 124.540 149.805 ;
        RECT 125.060 149.115 127.220 149.805 ;
        RECT 122.380 147.945 124.540 148.635 ;
        RECT 125.060 147.945 127.220 148.635 ;
        RECT 122.380 146.775 124.540 147.465 ;
        RECT 125.060 146.775 127.220 147.465 ;
        RECT 122.380 145.605 124.540 146.295 ;
        RECT 125.060 145.605 127.220 146.295 ;
        RECT 122.380 144.435 124.540 145.125 ;
        RECT 125.060 144.435 127.220 145.125 ;
        RECT 122.380 143.265 124.540 143.955 ;
        RECT 125.060 143.265 127.220 143.955 ;
        RECT 122.380 142.095 124.540 142.785 ;
        RECT 125.060 142.095 127.220 142.785 ;
        RECT 122.380 140.925 124.540 141.615 ;
        RECT 125.060 140.925 127.220 141.615 ;
        RECT 127.525 140.250 130.005 157.500 ;
        RECT 130.310 156.135 132.470 156.825 ;
        RECT 132.990 156.135 135.150 156.825 ;
        RECT 130.310 154.965 132.470 155.655 ;
        RECT 132.990 154.965 135.150 155.655 ;
        RECT 130.310 153.795 132.470 154.485 ;
        RECT 132.990 153.795 135.150 154.485 ;
        RECT 130.310 152.625 132.470 153.315 ;
        RECT 132.990 152.625 135.150 153.315 ;
        RECT 130.310 151.455 132.470 152.145 ;
        RECT 132.990 151.455 135.150 152.145 ;
        RECT 130.310 150.285 132.470 150.975 ;
        RECT 132.990 150.285 135.150 150.975 ;
        RECT 130.310 149.115 132.470 149.805 ;
        RECT 132.990 149.115 135.150 149.805 ;
        RECT 130.310 147.945 132.470 148.635 ;
        RECT 132.990 147.945 135.150 148.635 ;
        RECT 130.310 146.775 132.470 147.465 ;
        RECT 132.990 146.775 135.150 147.465 ;
        RECT 130.310 145.605 132.470 146.295 ;
        RECT 132.990 145.605 135.150 146.295 ;
        RECT 130.310 144.435 132.470 145.125 ;
        RECT 132.990 144.435 135.150 145.125 ;
        RECT 130.310 143.265 132.470 143.955 ;
        RECT 132.990 143.265 135.150 143.955 ;
        RECT 130.310 142.095 132.470 142.785 ;
        RECT 132.990 142.095 135.150 142.785 ;
        RECT 130.310 140.925 132.470 141.615 ;
        RECT 132.990 140.925 135.150 141.615 ;
        RECT 135.455 140.250 137.935 157.500 ;
        RECT 138.240 156.135 140.400 156.825 ;
        RECT 140.920 156.135 143.080 156.825 ;
        RECT 138.240 154.965 140.400 155.655 ;
        RECT 140.920 154.965 143.080 155.655 ;
        RECT 138.240 153.795 140.400 154.485 ;
        RECT 140.920 153.795 143.080 154.485 ;
        RECT 138.240 152.625 140.400 153.315 ;
        RECT 140.920 152.625 143.080 153.315 ;
        RECT 138.240 151.455 140.400 152.145 ;
        RECT 140.920 151.455 143.080 152.145 ;
        RECT 138.240 150.285 140.400 150.975 ;
        RECT 140.920 150.285 143.080 150.975 ;
        RECT 138.240 149.115 140.400 149.805 ;
        RECT 140.920 149.115 143.080 149.805 ;
        RECT 138.240 147.945 140.400 148.635 ;
        RECT 140.920 147.945 143.080 148.635 ;
        RECT 138.240 146.775 140.400 147.465 ;
        RECT 140.920 146.775 143.080 147.465 ;
        RECT 138.240 145.605 140.400 146.295 ;
        RECT 140.920 145.605 143.080 146.295 ;
        RECT 138.240 144.435 140.400 145.125 ;
        RECT 140.920 144.435 143.080 145.125 ;
        RECT 138.240 143.265 140.400 143.955 ;
        RECT 140.920 143.265 143.080 143.955 ;
        RECT 138.240 142.095 140.400 142.785 ;
        RECT 140.920 142.095 143.080 142.785 ;
        RECT 138.240 140.925 140.400 141.615 ;
        RECT 140.920 140.925 143.080 141.615 ;
        RECT 143.385 140.250 145.865 157.500 ;
        RECT 146.170 156.135 148.330 156.825 ;
        RECT 146.170 154.965 148.330 155.655 ;
        RECT 146.170 153.795 148.330 154.485 ;
        RECT 146.170 152.625 148.330 153.315 ;
        RECT 146.170 151.455 148.330 152.145 ;
        RECT 146.170 150.285 148.330 150.975 ;
        RECT 146.170 149.115 148.330 149.805 ;
        RECT 146.170 147.945 148.330 148.635 ;
        RECT 146.170 146.775 148.330 147.465 ;
        RECT 146.170 145.605 148.330 146.295 ;
        RECT 146.170 144.435 148.330 145.125 ;
        RECT 146.170 143.265 148.330 143.955 ;
        RECT 146.170 142.095 148.330 142.785 ;
        RECT 146.170 140.925 148.330 141.615 ;
        RECT 148.915 140.250 149.445 157.500 ;
        RECT 116.015 139.720 149.445 140.250 ;
        RECT 64.100 133.585 96.940 133.985 ;
        RECT 138.110 134.130 145.930 134.660 ;
        RECT 138.110 130.280 138.640 134.130 ;
        RECT 139.465 133.440 140.465 133.610 ;
        RECT 140.755 133.440 141.755 133.610 ;
        RECT 139.235 131.185 139.405 133.225 ;
        RECT 140.525 131.185 140.695 133.225 ;
        RECT 141.815 131.185 141.985 133.225 ;
        RECT 142.580 130.280 142.750 134.130 ;
        RECT 143.345 131.185 143.515 133.225 ;
        RECT 144.635 131.185 144.805 133.225 ;
        RECT 143.575 130.800 144.575 130.970 ;
        RECT 145.400 130.280 145.930 134.130 ;
        RECT 138.110 129.750 145.930 130.280 ;
        RECT 138.110 128.410 145.930 128.940 ;
        RECT 138.110 124.650 138.640 128.410 ;
        RECT 139.235 125.510 139.405 127.550 ;
        RECT 140.525 125.510 140.695 127.550 ;
        RECT 141.815 125.510 141.985 127.550 ;
        RECT 139.465 125.170 140.465 125.340 ;
        RECT 140.755 125.170 141.755 125.340 ;
        RECT 142.580 124.650 142.750 128.410 ;
        RECT 143.575 127.720 144.575 127.890 ;
        RECT 143.345 125.510 143.515 127.550 ;
        RECT 144.635 125.510 144.805 127.550 ;
        RECT 145.400 124.650 145.930 128.410 ;
        RECT 10.055 123.725 70.145 124.255 ;
        RECT 10.055 113.875 10.585 123.725 ;
        RECT 11.315 123.035 13.315 123.205 ;
        RECT 13.605 123.035 15.605 123.205 ;
        RECT 11.085 114.780 11.255 122.820 ;
        RECT 13.375 114.780 13.545 122.820 ;
        RECT 15.665 114.780 15.835 122.820 ;
        RECT 11.315 114.395 13.315 114.565 ;
        RECT 13.605 114.395 15.605 114.565 ;
        RECT 16.335 113.875 16.505 123.725 ;
        RECT 17.235 123.035 19.235 123.205 ;
        RECT 19.525 123.035 21.525 123.205 ;
        RECT 17.005 114.780 17.175 122.820 ;
        RECT 19.295 114.780 19.465 122.820 ;
        RECT 21.585 114.780 21.755 122.820 ;
        RECT 17.235 114.395 19.235 114.565 ;
        RECT 19.525 114.395 21.525 114.565 ;
        RECT 22.255 113.875 22.425 123.725 ;
        RECT 23.155 123.035 25.155 123.205 ;
        RECT 25.445 123.035 27.445 123.205 ;
        RECT 22.925 114.780 23.095 122.820 ;
        RECT 25.215 114.780 25.385 122.820 ;
        RECT 27.505 114.780 27.675 122.820 ;
        RECT 23.155 114.395 25.155 114.565 ;
        RECT 25.445 114.395 27.445 114.565 ;
        RECT 28.175 113.875 28.345 123.725 ;
        RECT 29.075 123.035 31.075 123.205 ;
        RECT 31.365 123.035 33.365 123.205 ;
        RECT 28.845 114.780 29.015 122.820 ;
        RECT 31.135 114.780 31.305 122.820 ;
        RECT 33.425 114.780 33.595 122.820 ;
        RECT 29.075 114.395 31.075 114.565 ;
        RECT 31.365 114.395 33.365 114.565 ;
        RECT 34.095 113.875 34.265 123.725 ;
        RECT 34.995 123.035 36.995 123.205 ;
        RECT 37.285 123.035 39.285 123.205 ;
        RECT 34.765 114.780 34.935 122.820 ;
        RECT 37.055 114.780 37.225 122.820 ;
        RECT 39.345 114.780 39.515 122.820 ;
        RECT 34.995 114.395 36.995 114.565 ;
        RECT 37.285 114.395 39.285 114.565 ;
        RECT 40.015 113.875 40.185 123.725 ;
        RECT 40.915 123.035 42.915 123.205 ;
        RECT 43.205 123.035 45.205 123.205 ;
        RECT 40.685 114.780 40.855 122.820 ;
        RECT 42.975 114.780 43.145 122.820 ;
        RECT 45.265 114.780 45.435 122.820 ;
        RECT 40.915 114.395 42.915 114.565 ;
        RECT 43.205 114.395 45.205 114.565 ;
        RECT 45.935 113.875 46.105 123.725 ;
        RECT 46.835 123.035 48.835 123.205 ;
        RECT 49.125 123.035 51.125 123.205 ;
        RECT 46.605 114.780 46.775 122.820 ;
        RECT 48.895 114.780 49.065 122.820 ;
        RECT 51.185 114.780 51.355 122.820 ;
        RECT 46.835 114.395 48.835 114.565 ;
        RECT 49.125 114.395 51.125 114.565 ;
        RECT 51.855 113.875 52.025 123.725 ;
        RECT 52.755 123.035 54.755 123.205 ;
        RECT 55.045 123.035 57.045 123.205 ;
        RECT 52.525 114.780 52.695 122.820 ;
        RECT 54.815 114.780 54.985 122.820 ;
        RECT 57.105 114.780 57.275 122.820 ;
        RECT 52.755 114.395 54.755 114.565 ;
        RECT 55.045 114.395 57.045 114.565 ;
        RECT 57.775 113.875 57.945 123.725 ;
        RECT 58.675 123.035 60.675 123.205 ;
        RECT 60.965 123.035 62.965 123.205 ;
        RECT 58.445 114.780 58.615 122.820 ;
        RECT 60.735 114.780 60.905 122.820 ;
        RECT 63.025 114.780 63.195 122.820 ;
        RECT 58.675 114.395 60.675 114.565 ;
        RECT 60.965 114.395 62.965 114.565 ;
        RECT 63.695 113.875 63.865 123.725 ;
        RECT 64.595 123.035 66.595 123.205 ;
        RECT 66.885 123.035 68.885 123.205 ;
        RECT 64.365 114.780 64.535 122.820 ;
        RECT 66.655 114.780 66.825 122.820 ;
        RECT 68.945 114.780 69.115 122.820 ;
        RECT 64.595 114.395 66.595 114.565 ;
        RECT 66.885 114.395 68.885 114.565 ;
        RECT 69.615 113.875 70.145 123.725 ;
        RECT 10.055 113.705 70.145 113.875 ;
        RECT 10.055 103.855 10.585 113.705 ;
        RECT 11.315 113.015 13.315 113.185 ;
        RECT 13.605 113.015 15.605 113.185 ;
        RECT 11.085 104.760 11.255 112.800 ;
        RECT 13.375 104.760 13.545 112.800 ;
        RECT 15.665 104.760 15.835 112.800 ;
        RECT 11.315 104.375 13.315 104.545 ;
        RECT 13.605 104.375 15.605 104.545 ;
        RECT 16.335 103.855 16.505 113.705 ;
        RECT 17.235 113.015 19.235 113.185 ;
        RECT 19.525 113.015 21.525 113.185 ;
        RECT 17.005 104.760 17.175 112.800 ;
        RECT 19.295 104.760 19.465 112.800 ;
        RECT 21.585 104.760 21.755 112.800 ;
        RECT 17.235 104.375 19.235 104.545 ;
        RECT 19.525 104.375 21.525 104.545 ;
        RECT 22.255 103.855 22.425 113.705 ;
        RECT 23.155 113.015 25.155 113.185 ;
        RECT 25.445 113.015 27.445 113.185 ;
        RECT 22.925 104.760 23.095 112.800 ;
        RECT 25.215 104.760 25.385 112.800 ;
        RECT 27.505 104.760 27.675 112.800 ;
        RECT 23.155 104.375 25.155 104.545 ;
        RECT 25.445 104.375 27.445 104.545 ;
        RECT 28.175 103.855 28.345 113.705 ;
        RECT 29.075 113.015 31.075 113.185 ;
        RECT 31.365 113.015 33.365 113.185 ;
        RECT 28.845 104.760 29.015 112.800 ;
        RECT 31.135 104.760 31.305 112.800 ;
        RECT 33.425 104.760 33.595 112.800 ;
        RECT 29.075 104.375 31.075 104.545 ;
        RECT 31.365 104.375 33.365 104.545 ;
        RECT 34.095 103.855 34.265 113.705 ;
        RECT 34.995 113.015 36.995 113.185 ;
        RECT 37.285 113.015 39.285 113.185 ;
        RECT 34.765 104.760 34.935 112.800 ;
        RECT 37.055 104.760 37.225 112.800 ;
        RECT 39.345 104.760 39.515 112.800 ;
        RECT 34.995 104.375 36.995 104.545 ;
        RECT 37.285 104.375 39.285 104.545 ;
        RECT 40.015 103.855 40.185 113.705 ;
        RECT 40.915 113.015 42.915 113.185 ;
        RECT 43.205 113.015 45.205 113.185 ;
        RECT 40.685 104.760 40.855 112.800 ;
        RECT 42.975 104.760 43.145 112.800 ;
        RECT 45.265 104.760 45.435 112.800 ;
        RECT 40.915 104.375 42.915 104.545 ;
        RECT 43.205 104.375 45.205 104.545 ;
        RECT 45.935 103.855 46.105 113.705 ;
        RECT 46.835 113.015 48.835 113.185 ;
        RECT 49.125 113.015 51.125 113.185 ;
        RECT 46.605 104.760 46.775 112.800 ;
        RECT 48.895 104.760 49.065 112.800 ;
        RECT 51.185 104.760 51.355 112.800 ;
        RECT 46.835 104.375 48.835 104.545 ;
        RECT 49.125 104.375 51.125 104.545 ;
        RECT 51.855 103.855 52.025 113.705 ;
        RECT 52.755 113.015 54.755 113.185 ;
        RECT 55.045 113.015 57.045 113.185 ;
        RECT 52.525 104.760 52.695 112.800 ;
        RECT 54.815 104.760 54.985 112.800 ;
        RECT 57.105 104.760 57.275 112.800 ;
        RECT 52.755 104.375 54.755 104.545 ;
        RECT 55.045 104.375 57.045 104.545 ;
        RECT 57.775 103.855 57.945 113.705 ;
        RECT 58.675 113.015 60.675 113.185 ;
        RECT 60.965 113.015 62.965 113.185 ;
        RECT 58.445 104.760 58.615 112.800 ;
        RECT 60.735 104.760 60.905 112.800 ;
        RECT 63.025 104.760 63.195 112.800 ;
        RECT 58.675 104.375 60.675 104.545 ;
        RECT 60.965 104.375 62.965 104.545 ;
        RECT 63.695 103.855 63.865 113.705 ;
        RECT 64.595 113.015 66.595 113.185 ;
        RECT 66.885 113.015 68.885 113.185 ;
        RECT 64.365 104.760 64.535 112.800 ;
        RECT 66.655 104.760 66.825 112.800 ;
        RECT 68.945 104.760 69.115 112.800 ;
        RECT 64.595 104.375 66.595 104.545 ;
        RECT 66.885 104.375 68.885 104.545 ;
        RECT 69.615 103.855 70.145 113.705 ;
        RECT 10.055 103.325 70.145 103.855 ;
        RECT 71.805 123.725 114.135 124.255 ;
        RECT 138.110 124.120 145.930 124.650 ;
        RECT 71.805 113.875 72.335 123.725 ;
        RECT 72.835 122.820 77.585 123.725 ;
        RECT 72.835 114.780 73.005 122.820 ;
        RECT 75.125 114.780 75.295 122.820 ;
        RECT 77.415 114.780 77.585 122.820 ;
        RECT 73.065 114.395 75.065 114.565 ;
        RECT 75.355 114.395 77.355 114.565 ;
        RECT 78.085 113.875 78.255 123.725 ;
        RECT 78.985 123.035 80.985 123.205 ;
        RECT 81.275 123.035 83.275 123.205 ;
        RECT 78.755 114.780 78.925 122.820 ;
        RECT 81.045 114.780 81.215 122.820 ;
        RECT 83.335 114.780 83.505 122.820 ;
        RECT 78.985 114.395 80.985 114.565 ;
        RECT 81.275 114.395 83.275 114.565 ;
        RECT 84.005 113.875 84.175 123.725 ;
        RECT 84.905 123.035 86.905 123.205 ;
        RECT 87.195 123.035 89.195 123.205 ;
        RECT 84.675 114.780 84.845 122.820 ;
        RECT 86.965 114.780 87.135 122.820 ;
        RECT 89.255 114.780 89.425 122.820 ;
        RECT 84.905 114.395 86.905 114.565 ;
        RECT 87.195 114.395 89.195 114.565 ;
        RECT 89.925 113.875 90.095 123.725 ;
        RECT 90.825 123.035 92.825 123.205 ;
        RECT 93.115 123.035 95.115 123.205 ;
        RECT 90.595 114.780 90.765 122.820 ;
        RECT 92.885 114.780 93.055 122.820 ;
        RECT 95.175 114.780 95.345 122.820 ;
        RECT 90.825 114.395 92.825 114.565 ;
        RECT 93.115 114.395 95.115 114.565 ;
        RECT 95.845 113.875 96.015 123.725 ;
        RECT 96.745 123.035 98.745 123.205 ;
        RECT 99.035 123.035 101.035 123.205 ;
        RECT 96.515 114.780 96.685 122.820 ;
        RECT 98.805 114.780 98.975 122.820 ;
        RECT 101.095 114.780 101.265 122.820 ;
        RECT 96.745 114.395 98.745 114.565 ;
        RECT 99.035 114.395 101.035 114.565 ;
        RECT 101.765 113.875 101.935 123.725 ;
        RECT 102.665 123.035 104.665 123.205 ;
        RECT 104.955 123.035 106.955 123.205 ;
        RECT 102.435 114.780 102.605 122.820 ;
        RECT 104.725 114.780 104.895 122.820 ;
        RECT 107.015 114.780 107.185 122.820 ;
        RECT 102.665 114.395 104.665 114.565 ;
        RECT 104.955 114.395 106.955 114.565 ;
        RECT 107.685 113.875 107.855 123.725 ;
        RECT 108.355 122.820 113.105 123.725 ;
        RECT 108.355 114.780 108.525 122.820 ;
        RECT 110.645 114.780 110.815 122.820 ;
        RECT 112.935 114.780 113.105 122.820 ;
        RECT 108.585 114.395 110.585 114.565 ;
        RECT 110.875 114.395 112.875 114.565 ;
        RECT 113.605 113.875 114.135 123.725 ;
        RECT 71.805 113.705 114.135 113.875 ;
        RECT 71.805 103.855 72.335 113.705 ;
        RECT 73.065 113.015 75.065 113.185 ;
        RECT 75.355 113.015 77.355 113.185 ;
        RECT 72.835 104.760 73.005 112.800 ;
        RECT 75.125 104.760 75.295 112.800 ;
        RECT 77.415 104.760 77.585 112.800 ;
        RECT 72.835 103.855 77.585 104.760 ;
        RECT 78.085 103.855 78.255 113.705 ;
        RECT 78.985 113.015 80.985 113.185 ;
        RECT 81.275 113.015 83.275 113.185 ;
        RECT 78.755 104.760 78.925 112.800 ;
        RECT 81.045 104.760 81.215 112.800 ;
        RECT 83.335 104.760 83.505 112.800 ;
        RECT 78.985 104.375 80.985 104.545 ;
        RECT 81.275 104.375 83.275 104.545 ;
        RECT 84.005 103.855 84.175 113.705 ;
        RECT 84.905 113.015 86.905 113.185 ;
        RECT 87.195 113.015 89.195 113.185 ;
        RECT 84.675 104.760 84.845 112.800 ;
        RECT 86.965 104.760 87.135 112.800 ;
        RECT 89.255 104.760 89.425 112.800 ;
        RECT 84.905 104.375 86.905 104.545 ;
        RECT 87.195 104.375 89.195 104.545 ;
        RECT 89.925 103.855 90.095 113.705 ;
        RECT 90.825 113.015 92.825 113.185 ;
        RECT 93.115 113.015 95.115 113.185 ;
        RECT 90.595 104.760 90.765 112.800 ;
        RECT 92.885 104.760 93.055 112.800 ;
        RECT 95.175 104.760 95.345 112.800 ;
        RECT 90.825 104.375 92.825 104.545 ;
        RECT 93.115 104.375 95.115 104.545 ;
        RECT 95.845 103.855 96.015 113.705 ;
        RECT 96.745 113.015 98.745 113.185 ;
        RECT 99.035 113.015 101.035 113.185 ;
        RECT 96.515 104.760 96.685 112.800 ;
        RECT 98.805 104.760 98.975 112.800 ;
        RECT 101.095 104.760 101.265 112.800 ;
        RECT 96.745 104.375 98.745 104.545 ;
        RECT 99.035 104.375 101.035 104.545 ;
        RECT 101.765 103.855 101.935 113.705 ;
        RECT 102.665 113.015 104.665 113.185 ;
        RECT 104.955 113.015 106.955 113.185 ;
        RECT 102.435 104.760 102.605 112.800 ;
        RECT 104.725 104.760 104.895 112.800 ;
        RECT 107.015 104.760 107.185 112.800 ;
        RECT 102.665 104.375 104.665 104.545 ;
        RECT 104.955 104.375 106.955 104.545 ;
        RECT 107.685 103.855 107.855 113.705 ;
        RECT 108.585 113.015 110.585 113.185 ;
        RECT 110.875 113.015 112.875 113.185 ;
        RECT 108.355 104.760 108.525 112.800 ;
        RECT 110.645 104.760 110.815 112.800 ;
        RECT 112.935 104.760 113.105 112.800 ;
        RECT 108.355 103.855 113.105 104.760 ;
        RECT 113.605 103.855 114.135 113.705 ;
        RECT 71.805 103.325 114.135 103.855 ;
        RECT 115.935 122.945 128.905 123.475 ;
        RECT 115.935 113.485 116.465 122.945 ;
        RECT 117.370 122.275 118.410 122.445 ;
        RECT 116.985 114.215 117.155 122.215 ;
        RECT 118.625 114.215 118.795 122.215 ;
        RECT 117.370 113.985 118.410 114.155 ;
        RECT 119.315 113.485 119.485 122.945 ;
        RECT 120.390 122.275 121.430 122.445 ;
        RECT 120.005 114.215 120.175 122.215 ;
        RECT 121.645 114.215 121.815 122.215 ;
        RECT 120.390 113.985 121.430 114.155 ;
        RECT 122.335 113.485 122.505 122.945 ;
        RECT 123.410 122.275 124.450 122.445 ;
        RECT 123.025 114.215 123.195 122.215 ;
        RECT 124.665 114.215 124.835 122.215 ;
        RECT 123.410 113.985 124.450 114.155 ;
        RECT 125.355 113.485 125.525 122.945 ;
        RECT 126.430 122.275 127.470 122.445 ;
        RECT 126.045 114.215 126.215 122.215 ;
        RECT 127.685 114.215 127.855 122.215 ;
        RECT 126.430 113.985 127.470 114.155 ;
        RECT 128.375 113.485 128.905 122.945 ;
        RECT 115.935 113.315 128.905 113.485 ;
        RECT 115.935 103.855 116.465 113.315 ;
        RECT 117.370 112.645 118.410 112.815 ;
        RECT 116.985 104.585 117.155 112.585 ;
        RECT 118.625 104.585 118.795 112.585 ;
        RECT 117.370 104.355 118.410 104.525 ;
        RECT 119.315 103.855 119.485 113.315 ;
        RECT 120.390 112.645 121.430 112.815 ;
        RECT 120.005 104.585 120.175 112.585 ;
        RECT 121.645 104.585 121.815 112.585 ;
        RECT 120.390 104.355 121.430 104.525 ;
        RECT 122.335 103.855 122.505 113.315 ;
        RECT 123.410 112.645 124.450 112.815 ;
        RECT 123.025 104.585 123.195 112.585 ;
        RECT 124.665 104.585 124.835 112.585 ;
        RECT 123.410 104.355 124.450 104.525 ;
        RECT 125.355 103.855 125.525 113.315 ;
        RECT 126.430 112.645 127.470 112.815 ;
        RECT 126.045 104.585 126.215 112.585 ;
        RECT 127.685 104.585 127.855 112.585 ;
        RECT 126.430 104.355 127.470 104.525 ;
        RECT 128.375 103.855 128.905 113.315 ;
        RECT 115.935 103.325 128.905 103.855 ;
        RECT 135.150 104.785 149.540 108.660 ;
        RECT 10.055 102.145 128.905 102.675 ;
        RECT 10.055 92.295 10.585 102.145 ;
        RECT 11.315 101.455 13.315 101.625 ;
        RECT 13.605 101.455 15.605 101.625 ;
        RECT 15.895 101.455 17.895 101.625 ;
        RECT 18.185 101.455 20.185 101.625 ;
        RECT 20.475 101.455 22.475 101.625 ;
        RECT 22.765 101.455 24.765 101.625 ;
        RECT 25.055 101.455 27.055 101.625 ;
        RECT 27.345 101.455 29.345 101.625 ;
        RECT 11.085 93.200 11.255 101.240 ;
        RECT 13.375 93.200 13.545 101.240 ;
        RECT 15.665 93.200 15.835 101.240 ;
        RECT 17.955 93.200 18.125 101.240 ;
        RECT 20.245 93.200 20.415 101.240 ;
        RECT 22.535 93.200 22.705 101.240 ;
        RECT 24.825 93.200 24.995 101.240 ;
        RECT 27.115 93.200 27.285 101.240 ;
        RECT 29.405 93.200 29.575 101.240 ;
        RECT 11.315 92.815 13.315 92.985 ;
        RECT 13.605 92.815 15.605 92.985 ;
        RECT 15.895 92.815 17.895 92.985 ;
        RECT 18.185 92.815 20.185 92.985 ;
        RECT 20.475 92.815 22.475 92.985 ;
        RECT 22.765 92.815 24.765 92.985 ;
        RECT 25.055 92.815 27.055 92.985 ;
        RECT 27.345 92.815 29.345 92.985 ;
        RECT 30.075 92.295 30.245 102.145 ;
        RECT 30.975 101.455 32.975 101.625 ;
        RECT 33.265 101.455 35.265 101.625 ;
        RECT 35.555 101.455 37.555 101.625 ;
        RECT 37.845 101.455 39.845 101.625 ;
        RECT 40.135 101.455 42.135 101.625 ;
        RECT 42.425 101.455 44.425 101.625 ;
        RECT 44.715 101.455 46.715 101.625 ;
        RECT 47.005 101.455 49.005 101.625 ;
        RECT 30.745 93.200 30.915 101.240 ;
        RECT 33.035 93.200 33.205 101.240 ;
        RECT 35.325 93.200 35.495 101.240 ;
        RECT 37.615 93.200 37.785 101.240 ;
        RECT 39.905 93.200 40.075 101.240 ;
        RECT 42.195 93.200 42.365 101.240 ;
        RECT 44.485 93.200 44.655 101.240 ;
        RECT 46.775 93.200 46.945 101.240 ;
        RECT 49.065 93.200 49.235 101.240 ;
        RECT 30.975 92.815 32.975 92.985 ;
        RECT 33.265 92.815 35.265 92.985 ;
        RECT 35.555 92.815 37.555 92.985 ;
        RECT 37.845 92.815 39.845 92.985 ;
        RECT 40.135 92.815 42.135 92.985 ;
        RECT 42.425 92.815 44.425 92.985 ;
        RECT 44.715 92.815 46.715 92.985 ;
        RECT 47.005 92.815 49.005 92.985 ;
        RECT 49.735 92.295 49.905 102.145 ;
        RECT 50.635 101.455 52.635 101.625 ;
        RECT 52.925 101.455 54.925 101.625 ;
        RECT 55.215 101.455 57.215 101.625 ;
        RECT 57.505 101.455 59.505 101.625 ;
        RECT 59.795 101.455 61.795 101.625 ;
        RECT 62.085 101.455 64.085 101.625 ;
        RECT 64.375 101.455 66.375 101.625 ;
        RECT 66.665 101.455 68.665 101.625 ;
        RECT 50.405 93.200 50.575 101.240 ;
        RECT 52.695 93.200 52.865 101.240 ;
        RECT 54.985 93.200 55.155 101.240 ;
        RECT 57.275 93.200 57.445 101.240 ;
        RECT 59.565 93.200 59.735 101.240 ;
        RECT 61.855 93.200 62.025 101.240 ;
        RECT 64.145 93.200 64.315 101.240 ;
        RECT 66.435 93.200 66.605 101.240 ;
        RECT 68.725 93.200 68.895 101.240 ;
        RECT 50.635 92.815 52.635 92.985 ;
        RECT 52.925 92.815 54.925 92.985 ;
        RECT 55.215 92.815 57.215 92.985 ;
        RECT 57.505 92.815 59.505 92.985 ;
        RECT 59.795 92.815 61.795 92.985 ;
        RECT 62.085 92.815 64.085 92.985 ;
        RECT 64.375 92.815 66.375 92.985 ;
        RECT 66.665 92.815 68.665 92.985 ;
        RECT 69.395 92.295 69.565 102.145 ;
        RECT 70.295 101.455 72.295 101.625 ;
        RECT 72.585 101.455 74.585 101.625 ;
        RECT 74.875 101.455 76.875 101.625 ;
        RECT 77.165 101.455 79.165 101.625 ;
        RECT 79.455 101.455 81.455 101.625 ;
        RECT 81.745 101.455 83.745 101.625 ;
        RECT 84.035 101.455 86.035 101.625 ;
        RECT 86.325 101.455 88.325 101.625 ;
        RECT 70.065 93.200 70.235 101.240 ;
        RECT 72.355 93.200 72.525 101.240 ;
        RECT 74.645 93.200 74.815 101.240 ;
        RECT 76.935 93.200 77.105 101.240 ;
        RECT 79.225 93.200 79.395 101.240 ;
        RECT 81.515 93.200 81.685 101.240 ;
        RECT 83.805 93.200 83.975 101.240 ;
        RECT 86.095 93.200 86.265 101.240 ;
        RECT 88.385 93.200 88.555 101.240 ;
        RECT 70.295 92.815 72.295 92.985 ;
        RECT 72.585 92.815 74.585 92.985 ;
        RECT 74.875 92.815 76.875 92.985 ;
        RECT 77.165 92.815 79.165 92.985 ;
        RECT 79.455 92.815 81.455 92.985 ;
        RECT 81.745 92.815 83.745 92.985 ;
        RECT 84.035 92.815 86.035 92.985 ;
        RECT 86.325 92.815 88.325 92.985 ;
        RECT 89.055 92.295 89.225 102.145 ;
        RECT 89.955 101.455 91.955 101.625 ;
        RECT 92.245 101.455 94.245 101.625 ;
        RECT 94.535 101.455 96.535 101.625 ;
        RECT 96.825 101.455 98.825 101.625 ;
        RECT 99.115 101.455 101.115 101.625 ;
        RECT 101.405 101.455 103.405 101.625 ;
        RECT 103.695 101.455 105.695 101.625 ;
        RECT 105.985 101.455 107.985 101.625 ;
        RECT 89.725 93.200 89.895 101.240 ;
        RECT 92.015 93.200 92.185 101.240 ;
        RECT 94.305 93.200 94.475 101.240 ;
        RECT 96.595 93.200 96.765 101.240 ;
        RECT 98.885 93.200 99.055 101.240 ;
        RECT 101.175 93.200 101.345 101.240 ;
        RECT 103.465 93.200 103.635 101.240 ;
        RECT 105.755 93.200 105.925 101.240 ;
        RECT 108.045 93.200 108.215 101.240 ;
        RECT 89.955 92.815 91.955 92.985 ;
        RECT 92.245 92.815 94.245 92.985 ;
        RECT 94.535 92.815 96.535 92.985 ;
        RECT 96.825 92.815 98.825 92.985 ;
        RECT 99.115 92.815 101.115 92.985 ;
        RECT 101.405 92.815 103.405 92.985 ;
        RECT 103.695 92.815 105.695 92.985 ;
        RECT 105.985 92.815 107.985 92.985 ;
        RECT 108.715 92.295 108.885 102.145 ;
        RECT 109.615 101.455 111.615 101.625 ;
        RECT 111.905 101.455 113.905 101.625 ;
        RECT 114.195 101.455 116.195 101.625 ;
        RECT 116.485 101.455 118.485 101.625 ;
        RECT 118.775 101.455 120.775 101.625 ;
        RECT 121.065 101.455 123.065 101.625 ;
        RECT 123.355 101.455 125.355 101.625 ;
        RECT 125.645 101.455 127.645 101.625 ;
        RECT 109.385 93.200 109.555 101.240 ;
        RECT 111.675 93.200 111.845 101.240 ;
        RECT 113.965 93.200 114.135 101.240 ;
        RECT 116.255 93.200 116.425 101.240 ;
        RECT 118.545 93.200 118.715 101.240 ;
        RECT 120.835 93.200 121.005 101.240 ;
        RECT 123.125 93.200 123.295 101.240 ;
        RECT 125.415 93.200 125.585 101.240 ;
        RECT 127.705 93.200 127.875 101.240 ;
        RECT 109.615 92.815 111.615 92.985 ;
        RECT 111.905 92.815 113.905 92.985 ;
        RECT 114.195 92.815 116.195 92.985 ;
        RECT 116.485 92.815 118.485 92.985 ;
        RECT 118.775 92.815 120.775 92.985 ;
        RECT 121.065 92.815 123.065 92.985 ;
        RECT 123.355 92.815 125.355 92.985 ;
        RECT 125.645 92.815 127.645 92.985 ;
        RECT 128.375 92.295 128.905 102.145 ;
        RECT 10.055 92.125 128.905 92.295 ;
        RECT 10.055 82.275 10.585 92.125 ;
        RECT 11.315 91.435 13.315 91.605 ;
        RECT 13.605 91.435 15.605 91.605 ;
        RECT 15.895 91.435 17.895 91.605 ;
        RECT 18.185 91.435 20.185 91.605 ;
        RECT 20.475 91.435 22.475 91.605 ;
        RECT 22.765 91.435 24.765 91.605 ;
        RECT 25.055 91.435 27.055 91.605 ;
        RECT 27.345 91.435 29.345 91.605 ;
        RECT 11.085 83.180 11.255 91.220 ;
        RECT 13.375 83.180 13.545 91.220 ;
        RECT 15.665 83.180 15.835 91.220 ;
        RECT 17.955 83.180 18.125 91.220 ;
        RECT 20.245 83.180 20.415 91.220 ;
        RECT 22.535 83.180 22.705 91.220 ;
        RECT 24.825 83.180 24.995 91.220 ;
        RECT 27.115 83.180 27.285 91.220 ;
        RECT 29.405 83.180 29.575 91.220 ;
        RECT 11.315 82.795 13.315 82.965 ;
        RECT 13.605 82.795 15.605 82.965 ;
        RECT 15.895 82.795 17.895 82.965 ;
        RECT 18.185 82.795 20.185 82.965 ;
        RECT 20.475 82.795 22.475 82.965 ;
        RECT 22.765 82.795 24.765 82.965 ;
        RECT 25.055 82.795 27.055 82.965 ;
        RECT 27.345 82.795 29.345 82.965 ;
        RECT 30.075 82.275 30.245 92.125 ;
        RECT 30.975 91.435 32.975 91.605 ;
        RECT 33.265 91.435 35.265 91.605 ;
        RECT 35.555 91.435 37.555 91.605 ;
        RECT 37.845 91.435 39.845 91.605 ;
        RECT 40.135 91.435 42.135 91.605 ;
        RECT 42.425 91.435 44.425 91.605 ;
        RECT 44.715 91.435 46.715 91.605 ;
        RECT 47.005 91.435 49.005 91.605 ;
        RECT 30.745 83.180 30.915 91.220 ;
        RECT 33.035 83.180 33.205 91.220 ;
        RECT 35.325 83.180 35.495 91.220 ;
        RECT 37.615 83.180 37.785 91.220 ;
        RECT 39.905 83.180 40.075 91.220 ;
        RECT 42.195 83.180 42.365 91.220 ;
        RECT 44.485 83.180 44.655 91.220 ;
        RECT 46.775 83.180 46.945 91.220 ;
        RECT 49.065 83.180 49.235 91.220 ;
        RECT 30.975 82.795 32.975 82.965 ;
        RECT 33.265 82.795 35.265 82.965 ;
        RECT 35.555 82.795 37.555 82.965 ;
        RECT 37.845 82.795 39.845 82.965 ;
        RECT 40.135 82.795 42.135 82.965 ;
        RECT 42.425 82.795 44.425 82.965 ;
        RECT 44.715 82.795 46.715 82.965 ;
        RECT 47.005 82.795 49.005 82.965 ;
        RECT 49.735 82.275 49.905 92.125 ;
        RECT 50.635 91.435 52.635 91.605 ;
        RECT 52.925 91.435 54.925 91.605 ;
        RECT 55.215 91.435 57.215 91.605 ;
        RECT 57.505 91.435 59.505 91.605 ;
        RECT 59.795 91.435 61.795 91.605 ;
        RECT 62.085 91.435 64.085 91.605 ;
        RECT 64.375 91.435 66.375 91.605 ;
        RECT 66.665 91.435 68.665 91.605 ;
        RECT 50.405 83.180 50.575 91.220 ;
        RECT 52.695 83.180 52.865 91.220 ;
        RECT 54.985 83.180 55.155 91.220 ;
        RECT 57.275 83.180 57.445 91.220 ;
        RECT 59.565 83.180 59.735 91.220 ;
        RECT 61.855 83.180 62.025 91.220 ;
        RECT 64.145 83.180 64.315 91.220 ;
        RECT 66.435 83.180 66.605 91.220 ;
        RECT 68.725 83.180 68.895 91.220 ;
        RECT 50.635 82.795 52.635 82.965 ;
        RECT 52.925 82.795 54.925 82.965 ;
        RECT 55.215 82.795 57.215 82.965 ;
        RECT 57.505 82.795 59.505 82.965 ;
        RECT 59.795 82.795 61.795 82.965 ;
        RECT 62.085 82.795 64.085 82.965 ;
        RECT 64.375 82.795 66.375 82.965 ;
        RECT 66.665 82.795 68.665 82.965 ;
        RECT 69.395 82.275 69.565 92.125 ;
        RECT 70.295 91.435 72.295 91.605 ;
        RECT 72.585 91.435 74.585 91.605 ;
        RECT 74.875 91.435 76.875 91.605 ;
        RECT 77.165 91.435 79.165 91.605 ;
        RECT 79.455 91.435 81.455 91.605 ;
        RECT 81.745 91.435 83.745 91.605 ;
        RECT 84.035 91.435 86.035 91.605 ;
        RECT 86.325 91.435 88.325 91.605 ;
        RECT 70.065 83.180 70.235 91.220 ;
        RECT 72.355 83.180 72.525 91.220 ;
        RECT 74.645 83.180 74.815 91.220 ;
        RECT 76.935 83.180 77.105 91.220 ;
        RECT 79.225 83.180 79.395 91.220 ;
        RECT 81.515 83.180 81.685 91.220 ;
        RECT 83.805 83.180 83.975 91.220 ;
        RECT 86.095 83.180 86.265 91.220 ;
        RECT 88.385 83.180 88.555 91.220 ;
        RECT 70.295 82.795 72.295 82.965 ;
        RECT 72.585 82.795 74.585 82.965 ;
        RECT 74.875 82.795 76.875 82.965 ;
        RECT 77.165 82.795 79.165 82.965 ;
        RECT 79.455 82.795 81.455 82.965 ;
        RECT 81.745 82.795 83.745 82.965 ;
        RECT 84.035 82.795 86.035 82.965 ;
        RECT 86.325 82.795 88.325 82.965 ;
        RECT 89.055 82.275 89.225 92.125 ;
        RECT 89.955 91.435 91.955 91.605 ;
        RECT 92.245 91.435 94.245 91.605 ;
        RECT 94.535 91.435 96.535 91.605 ;
        RECT 96.825 91.435 98.825 91.605 ;
        RECT 99.115 91.435 101.115 91.605 ;
        RECT 101.405 91.435 103.405 91.605 ;
        RECT 103.695 91.435 105.695 91.605 ;
        RECT 105.985 91.435 107.985 91.605 ;
        RECT 89.725 83.180 89.895 91.220 ;
        RECT 92.015 83.180 92.185 91.220 ;
        RECT 94.305 83.180 94.475 91.220 ;
        RECT 96.595 83.180 96.765 91.220 ;
        RECT 98.885 83.180 99.055 91.220 ;
        RECT 101.175 83.180 101.345 91.220 ;
        RECT 103.465 83.180 103.635 91.220 ;
        RECT 105.755 83.180 105.925 91.220 ;
        RECT 108.045 83.180 108.215 91.220 ;
        RECT 89.955 82.795 91.955 82.965 ;
        RECT 92.245 82.795 94.245 82.965 ;
        RECT 94.535 82.795 96.535 82.965 ;
        RECT 96.825 82.795 98.825 82.965 ;
        RECT 99.115 82.795 101.115 82.965 ;
        RECT 101.405 82.795 103.405 82.965 ;
        RECT 103.695 82.795 105.695 82.965 ;
        RECT 105.985 82.795 107.985 82.965 ;
        RECT 108.715 82.275 108.885 92.125 ;
        RECT 109.615 91.435 111.615 91.605 ;
        RECT 111.905 91.435 113.905 91.605 ;
        RECT 114.195 91.435 116.195 91.605 ;
        RECT 116.485 91.435 118.485 91.605 ;
        RECT 118.775 91.435 120.775 91.605 ;
        RECT 121.065 91.435 123.065 91.605 ;
        RECT 123.355 91.435 125.355 91.605 ;
        RECT 125.645 91.435 127.645 91.605 ;
        RECT 109.385 83.180 109.555 91.220 ;
        RECT 111.675 83.180 111.845 91.220 ;
        RECT 113.965 83.180 114.135 91.220 ;
        RECT 116.255 83.180 116.425 91.220 ;
        RECT 118.545 83.180 118.715 91.220 ;
        RECT 120.835 83.180 121.005 91.220 ;
        RECT 123.125 83.180 123.295 91.220 ;
        RECT 125.415 83.180 125.585 91.220 ;
        RECT 127.705 83.180 127.875 91.220 ;
        RECT 109.615 82.795 111.615 82.965 ;
        RECT 111.905 82.795 113.905 82.965 ;
        RECT 114.195 82.795 116.195 82.965 ;
        RECT 116.485 82.795 118.485 82.965 ;
        RECT 118.775 82.795 120.775 82.965 ;
        RECT 121.065 82.795 123.065 82.965 ;
        RECT 123.355 82.795 125.355 82.965 ;
        RECT 125.645 82.795 127.645 82.965 ;
        RECT 128.375 82.275 128.905 92.125 ;
        RECT 10.055 82.105 128.905 82.275 ;
        RECT 10.055 72.255 10.585 82.105 ;
        RECT 11.315 81.415 13.315 81.585 ;
        RECT 13.605 81.415 15.605 81.585 ;
        RECT 15.895 81.415 17.895 81.585 ;
        RECT 18.185 81.415 20.185 81.585 ;
        RECT 20.475 81.415 22.475 81.585 ;
        RECT 22.765 81.415 24.765 81.585 ;
        RECT 25.055 81.415 27.055 81.585 ;
        RECT 27.345 81.415 29.345 81.585 ;
        RECT 11.085 73.160 11.255 81.200 ;
        RECT 13.375 73.160 13.545 81.200 ;
        RECT 15.665 73.160 15.835 81.200 ;
        RECT 17.955 73.160 18.125 81.200 ;
        RECT 20.245 73.160 20.415 81.200 ;
        RECT 22.535 73.160 22.705 81.200 ;
        RECT 24.825 73.160 24.995 81.200 ;
        RECT 27.115 73.160 27.285 81.200 ;
        RECT 29.405 73.160 29.575 81.200 ;
        RECT 11.315 72.775 13.315 72.945 ;
        RECT 13.605 72.775 15.605 72.945 ;
        RECT 15.895 72.775 17.895 72.945 ;
        RECT 18.185 72.775 20.185 72.945 ;
        RECT 20.475 72.775 22.475 72.945 ;
        RECT 22.765 72.775 24.765 72.945 ;
        RECT 25.055 72.775 27.055 72.945 ;
        RECT 27.345 72.775 29.345 72.945 ;
        RECT 30.075 72.255 30.245 82.105 ;
        RECT 30.975 81.415 32.975 81.585 ;
        RECT 33.265 81.415 35.265 81.585 ;
        RECT 35.555 81.415 37.555 81.585 ;
        RECT 37.845 81.415 39.845 81.585 ;
        RECT 40.135 81.415 42.135 81.585 ;
        RECT 42.425 81.415 44.425 81.585 ;
        RECT 44.715 81.415 46.715 81.585 ;
        RECT 47.005 81.415 49.005 81.585 ;
        RECT 30.745 73.160 30.915 81.200 ;
        RECT 33.035 73.160 33.205 81.200 ;
        RECT 35.325 73.160 35.495 81.200 ;
        RECT 37.615 73.160 37.785 81.200 ;
        RECT 39.905 73.160 40.075 81.200 ;
        RECT 42.195 73.160 42.365 81.200 ;
        RECT 44.485 73.160 44.655 81.200 ;
        RECT 46.775 73.160 46.945 81.200 ;
        RECT 49.065 73.160 49.235 81.200 ;
        RECT 30.975 72.775 32.975 72.945 ;
        RECT 33.265 72.775 35.265 72.945 ;
        RECT 35.555 72.775 37.555 72.945 ;
        RECT 37.845 72.775 39.845 72.945 ;
        RECT 40.135 72.775 42.135 72.945 ;
        RECT 42.425 72.775 44.425 72.945 ;
        RECT 44.715 72.775 46.715 72.945 ;
        RECT 47.005 72.775 49.005 72.945 ;
        RECT 49.735 72.255 49.905 82.105 ;
        RECT 50.635 81.415 52.635 81.585 ;
        RECT 52.925 81.415 54.925 81.585 ;
        RECT 55.215 81.415 57.215 81.585 ;
        RECT 57.505 81.415 59.505 81.585 ;
        RECT 59.795 81.415 61.795 81.585 ;
        RECT 62.085 81.415 64.085 81.585 ;
        RECT 64.375 81.415 66.375 81.585 ;
        RECT 66.665 81.415 68.665 81.585 ;
        RECT 50.405 73.160 50.575 81.200 ;
        RECT 52.695 73.160 52.865 81.200 ;
        RECT 54.985 73.160 55.155 81.200 ;
        RECT 57.275 73.160 57.445 81.200 ;
        RECT 59.565 73.160 59.735 81.200 ;
        RECT 61.855 73.160 62.025 81.200 ;
        RECT 64.145 73.160 64.315 81.200 ;
        RECT 66.435 73.160 66.605 81.200 ;
        RECT 68.725 73.160 68.895 81.200 ;
        RECT 50.635 72.775 52.635 72.945 ;
        RECT 52.925 72.775 54.925 72.945 ;
        RECT 55.215 72.775 57.215 72.945 ;
        RECT 57.505 72.775 59.505 72.945 ;
        RECT 59.795 72.775 61.795 72.945 ;
        RECT 62.085 72.775 64.085 72.945 ;
        RECT 64.375 72.775 66.375 72.945 ;
        RECT 66.665 72.775 68.665 72.945 ;
        RECT 69.395 72.255 69.565 82.105 ;
        RECT 70.295 81.415 72.295 81.585 ;
        RECT 72.585 81.415 74.585 81.585 ;
        RECT 74.875 81.415 76.875 81.585 ;
        RECT 77.165 81.415 79.165 81.585 ;
        RECT 79.455 81.415 81.455 81.585 ;
        RECT 81.745 81.415 83.745 81.585 ;
        RECT 84.035 81.415 86.035 81.585 ;
        RECT 86.325 81.415 88.325 81.585 ;
        RECT 70.065 73.160 70.235 81.200 ;
        RECT 72.355 73.160 72.525 81.200 ;
        RECT 74.645 73.160 74.815 81.200 ;
        RECT 76.935 73.160 77.105 81.200 ;
        RECT 79.225 73.160 79.395 81.200 ;
        RECT 81.515 73.160 81.685 81.200 ;
        RECT 83.805 73.160 83.975 81.200 ;
        RECT 86.095 73.160 86.265 81.200 ;
        RECT 88.385 73.160 88.555 81.200 ;
        RECT 70.295 72.775 72.295 72.945 ;
        RECT 72.585 72.775 74.585 72.945 ;
        RECT 74.875 72.775 76.875 72.945 ;
        RECT 77.165 72.775 79.165 72.945 ;
        RECT 79.455 72.775 81.455 72.945 ;
        RECT 81.745 72.775 83.745 72.945 ;
        RECT 84.035 72.775 86.035 72.945 ;
        RECT 86.325 72.775 88.325 72.945 ;
        RECT 89.055 72.255 89.225 82.105 ;
        RECT 89.955 81.415 91.955 81.585 ;
        RECT 92.245 81.415 94.245 81.585 ;
        RECT 94.535 81.415 96.535 81.585 ;
        RECT 96.825 81.415 98.825 81.585 ;
        RECT 99.115 81.415 101.115 81.585 ;
        RECT 101.405 81.415 103.405 81.585 ;
        RECT 103.695 81.415 105.695 81.585 ;
        RECT 105.985 81.415 107.985 81.585 ;
        RECT 89.725 73.160 89.895 81.200 ;
        RECT 92.015 73.160 92.185 81.200 ;
        RECT 94.305 73.160 94.475 81.200 ;
        RECT 96.595 73.160 96.765 81.200 ;
        RECT 98.885 73.160 99.055 81.200 ;
        RECT 101.175 73.160 101.345 81.200 ;
        RECT 103.465 73.160 103.635 81.200 ;
        RECT 105.755 73.160 105.925 81.200 ;
        RECT 108.045 73.160 108.215 81.200 ;
        RECT 89.955 72.775 91.955 72.945 ;
        RECT 92.245 72.775 94.245 72.945 ;
        RECT 94.535 72.775 96.535 72.945 ;
        RECT 96.825 72.775 98.825 72.945 ;
        RECT 99.115 72.775 101.115 72.945 ;
        RECT 101.405 72.775 103.405 72.945 ;
        RECT 103.695 72.775 105.695 72.945 ;
        RECT 105.985 72.775 107.985 72.945 ;
        RECT 108.715 72.255 108.885 82.105 ;
        RECT 109.615 81.415 111.615 81.585 ;
        RECT 111.905 81.415 113.905 81.585 ;
        RECT 114.195 81.415 116.195 81.585 ;
        RECT 116.485 81.415 118.485 81.585 ;
        RECT 118.775 81.415 120.775 81.585 ;
        RECT 121.065 81.415 123.065 81.585 ;
        RECT 123.355 81.415 125.355 81.585 ;
        RECT 125.645 81.415 127.645 81.585 ;
        RECT 109.385 73.160 109.555 81.200 ;
        RECT 111.675 73.160 111.845 81.200 ;
        RECT 113.965 73.160 114.135 81.200 ;
        RECT 116.255 73.160 116.425 81.200 ;
        RECT 118.545 73.160 118.715 81.200 ;
        RECT 120.835 73.160 121.005 81.200 ;
        RECT 123.125 73.160 123.295 81.200 ;
        RECT 125.415 73.160 125.585 81.200 ;
        RECT 127.705 73.160 127.875 81.200 ;
        RECT 109.615 72.775 111.615 72.945 ;
        RECT 111.905 72.775 113.905 72.945 ;
        RECT 114.195 72.775 116.195 72.945 ;
        RECT 116.485 72.775 118.485 72.945 ;
        RECT 118.775 72.775 120.775 72.945 ;
        RECT 121.065 72.775 123.065 72.945 ;
        RECT 123.355 72.775 125.355 72.945 ;
        RECT 125.645 72.775 127.645 72.945 ;
        RECT 128.375 72.255 128.905 82.105 ;
        RECT 10.055 72.085 128.905 72.255 ;
        RECT 10.055 62.235 10.585 72.085 ;
        RECT 11.315 71.395 13.315 71.565 ;
        RECT 13.605 71.395 15.605 71.565 ;
        RECT 15.895 71.395 17.895 71.565 ;
        RECT 18.185 71.395 20.185 71.565 ;
        RECT 20.475 71.395 22.475 71.565 ;
        RECT 22.765 71.395 24.765 71.565 ;
        RECT 25.055 71.395 27.055 71.565 ;
        RECT 27.345 71.395 29.345 71.565 ;
        RECT 11.085 63.140 11.255 71.180 ;
        RECT 13.375 63.140 13.545 71.180 ;
        RECT 15.665 63.140 15.835 71.180 ;
        RECT 17.955 63.140 18.125 71.180 ;
        RECT 20.245 63.140 20.415 71.180 ;
        RECT 22.535 63.140 22.705 71.180 ;
        RECT 24.825 63.140 24.995 71.180 ;
        RECT 27.115 63.140 27.285 71.180 ;
        RECT 29.405 63.140 29.575 71.180 ;
        RECT 11.315 62.755 13.315 62.925 ;
        RECT 13.605 62.755 15.605 62.925 ;
        RECT 15.895 62.755 17.895 62.925 ;
        RECT 18.185 62.755 20.185 62.925 ;
        RECT 20.475 62.755 22.475 62.925 ;
        RECT 22.765 62.755 24.765 62.925 ;
        RECT 25.055 62.755 27.055 62.925 ;
        RECT 27.345 62.755 29.345 62.925 ;
        RECT 30.075 62.235 30.245 72.085 ;
        RECT 30.975 71.395 32.975 71.565 ;
        RECT 33.265 71.395 35.265 71.565 ;
        RECT 35.555 71.395 37.555 71.565 ;
        RECT 37.845 71.395 39.845 71.565 ;
        RECT 40.135 71.395 42.135 71.565 ;
        RECT 42.425 71.395 44.425 71.565 ;
        RECT 44.715 71.395 46.715 71.565 ;
        RECT 47.005 71.395 49.005 71.565 ;
        RECT 30.745 63.140 30.915 71.180 ;
        RECT 33.035 63.140 33.205 71.180 ;
        RECT 35.325 63.140 35.495 71.180 ;
        RECT 37.615 63.140 37.785 71.180 ;
        RECT 39.905 63.140 40.075 71.180 ;
        RECT 42.195 63.140 42.365 71.180 ;
        RECT 44.485 63.140 44.655 71.180 ;
        RECT 46.775 63.140 46.945 71.180 ;
        RECT 49.065 63.140 49.235 71.180 ;
        RECT 30.975 62.755 32.975 62.925 ;
        RECT 33.265 62.755 35.265 62.925 ;
        RECT 35.555 62.755 37.555 62.925 ;
        RECT 37.845 62.755 39.845 62.925 ;
        RECT 40.135 62.755 42.135 62.925 ;
        RECT 42.425 62.755 44.425 62.925 ;
        RECT 44.715 62.755 46.715 62.925 ;
        RECT 47.005 62.755 49.005 62.925 ;
        RECT 49.735 62.235 49.905 72.085 ;
        RECT 50.635 71.395 52.635 71.565 ;
        RECT 52.925 71.395 54.925 71.565 ;
        RECT 55.215 71.395 57.215 71.565 ;
        RECT 57.505 71.395 59.505 71.565 ;
        RECT 59.795 71.395 61.795 71.565 ;
        RECT 62.085 71.395 64.085 71.565 ;
        RECT 64.375 71.395 66.375 71.565 ;
        RECT 66.665 71.395 68.665 71.565 ;
        RECT 50.405 63.140 50.575 71.180 ;
        RECT 52.695 63.140 52.865 71.180 ;
        RECT 54.985 63.140 55.155 71.180 ;
        RECT 57.275 63.140 57.445 71.180 ;
        RECT 59.565 63.140 59.735 71.180 ;
        RECT 61.855 63.140 62.025 71.180 ;
        RECT 64.145 63.140 64.315 71.180 ;
        RECT 66.435 63.140 66.605 71.180 ;
        RECT 68.725 63.140 68.895 71.180 ;
        RECT 50.635 62.755 52.635 62.925 ;
        RECT 52.925 62.755 54.925 62.925 ;
        RECT 55.215 62.755 57.215 62.925 ;
        RECT 57.505 62.755 59.505 62.925 ;
        RECT 59.795 62.755 61.795 62.925 ;
        RECT 62.085 62.755 64.085 62.925 ;
        RECT 64.375 62.755 66.375 62.925 ;
        RECT 66.665 62.755 68.665 62.925 ;
        RECT 69.395 62.235 69.565 72.085 ;
        RECT 70.295 71.395 72.295 71.565 ;
        RECT 72.585 71.395 74.585 71.565 ;
        RECT 74.875 71.395 76.875 71.565 ;
        RECT 77.165 71.395 79.165 71.565 ;
        RECT 79.455 71.395 81.455 71.565 ;
        RECT 81.745 71.395 83.745 71.565 ;
        RECT 84.035 71.395 86.035 71.565 ;
        RECT 86.325 71.395 88.325 71.565 ;
        RECT 70.065 63.140 70.235 71.180 ;
        RECT 72.355 63.140 72.525 71.180 ;
        RECT 74.645 63.140 74.815 71.180 ;
        RECT 76.935 63.140 77.105 71.180 ;
        RECT 79.225 63.140 79.395 71.180 ;
        RECT 81.515 63.140 81.685 71.180 ;
        RECT 83.805 63.140 83.975 71.180 ;
        RECT 86.095 63.140 86.265 71.180 ;
        RECT 88.385 63.140 88.555 71.180 ;
        RECT 70.295 62.755 72.295 62.925 ;
        RECT 72.585 62.755 74.585 62.925 ;
        RECT 74.875 62.755 76.875 62.925 ;
        RECT 77.165 62.755 79.165 62.925 ;
        RECT 79.455 62.755 81.455 62.925 ;
        RECT 81.745 62.755 83.745 62.925 ;
        RECT 84.035 62.755 86.035 62.925 ;
        RECT 86.325 62.755 88.325 62.925 ;
        RECT 89.055 62.235 89.225 72.085 ;
        RECT 89.955 71.395 91.955 71.565 ;
        RECT 92.245 71.395 94.245 71.565 ;
        RECT 94.535 71.395 96.535 71.565 ;
        RECT 96.825 71.395 98.825 71.565 ;
        RECT 99.115 71.395 101.115 71.565 ;
        RECT 101.405 71.395 103.405 71.565 ;
        RECT 103.695 71.395 105.695 71.565 ;
        RECT 105.985 71.395 107.985 71.565 ;
        RECT 89.725 63.140 89.895 71.180 ;
        RECT 92.015 63.140 92.185 71.180 ;
        RECT 94.305 63.140 94.475 71.180 ;
        RECT 96.595 63.140 96.765 71.180 ;
        RECT 98.885 63.140 99.055 71.180 ;
        RECT 101.175 63.140 101.345 71.180 ;
        RECT 103.465 63.140 103.635 71.180 ;
        RECT 105.755 63.140 105.925 71.180 ;
        RECT 108.045 63.140 108.215 71.180 ;
        RECT 89.955 62.755 91.955 62.925 ;
        RECT 92.245 62.755 94.245 62.925 ;
        RECT 94.535 62.755 96.535 62.925 ;
        RECT 96.825 62.755 98.825 62.925 ;
        RECT 99.115 62.755 101.115 62.925 ;
        RECT 101.405 62.755 103.405 62.925 ;
        RECT 103.695 62.755 105.695 62.925 ;
        RECT 105.985 62.755 107.985 62.925 ;
        RECT 108.715 62.235 108.885 72.085 ;
        RECT 109.615 71.395 111.615 71.565 ;
        RECT 111.905 71.395 113.905 71.565 ;
        RECT 114.195 71.395 116.195 71.565 ;
        RECT 116.485 71.395 118.485 71.565 ;
        RECT 118.775 71.395 120.775 71.565 ;
        RECT 121.065 71.395 123.065 71.565 ;
        RECT 123.355 71.395 125.355 71.565 ;
        RECT 125.645 71.395 127.645 71.565 ;
        RECT 109.385 63.140 109.555 71.180 ;
        RECT 111.675 63.140 111.845 71.180 ;
        RECT 113.965 63.140 114.135 71.180 ;
        RECT 116.255 63.140 116.425 71.180 ;
        RECT 118.545 63.140 118.715 71.180 ;
        RECT 120.835 63.140 121.005 71.180 ;
        RECT 123.125 63.140 123.295 71.180 ;
        RECT 125.415 63.140 125.585 71.180 ;
        RECT 127.705 63.140 127.875 71.180 ;
        RECT 109.615 62.755 111.615 62.925 ;
        RECT 111.905 62.755 113.905 62.925 ;
        RECT 114.195 62.755 116.195 62.925 ;
        RECT 116.485 62.755 118.485 62.925 ;
        RECT 118.775 62.755 120.775 62.925 ;
        RECT 121.065 62.755 123.065 62.925 ;
        RECT 123.355 62.755 125.355 62.925 ;
        RECT 125.645 62.755 127.645 62.925 ;
        RECT 128.375 62.235 128.905 72.085 ;
        RECT 10.055 62.065 128.905 62.235 ;
        RECT 10.055 52.215 10.585 62.065 ;
        RECT 11.315 61.375 13.315 61.545 ;
        RECT 13.605 61.375 15.605 61.545 ;
        RECT 15.895 61.375 17.895 61.545 ;
        RECT 18.185 61.375 20.185 61.545 ;
        RECT 20.475 61.375 22.475 61.545 ;
        RECT 22.765 61.375 24.765 61.545 ;
        RECT 25.055 61.375 27.055 61.545 ;
        RECT 27.345 61.375 29.345 61.545 ;
        RECT 11.085 53.120 11.255 61.160 ;
        RECT 13.375 53.120 13.545 61.160 ;
        RECT 15.665 53.120 15.835 61.160 ;
        RECT 17.955 53.120 18.125 61.160 ;
        RECT 20.245 53.120 20.415 61.160 ;
        RECT 22.535 53.120 22.705 61.160 ;
        RECT 24.825 53.120 24.995 61.160 ;
        RECT 27.115 53.120 27.285 61.160 ;
        RECT 29.405 53.120 29.575 61.160 ;
        RECT 11.315 52.735 13.315 52.905 ;
        RECT 13.605 52.735 15.605 52.905 ;
        RECT 15.895 52.735 17.895 52.905 ;
        RECT 18.185 52.735 20.185 52.905 ;
        RECT 20.475 52.735 22.475 52.905 ;
        RECT 22.765 52.735 24.765 52.905 ;
        RECT 25.055 52.735 27.055 52.905 ;
        RECT 27.345 52.735 29.345 52.905 ;
        RECT 30.075 52.215 30.245 62.065 ;
        RECT 30.975 61.375 32.975 61.545 ;
        RECT 33.265 61.375 35.265 61.545 ;
        RECT 35.555 61.375 37.555 61.545 ;
        RECT 37.845 61.375 39.845 61.545 ;
        RECT 40.135 61.375 42.135 61.545 ;
        RECT 42.425 61.375 44.425 61.545 ;
        RECT 44.715 61.375 46.715 61.545 ;
        RECT 47.005 61.375 49.005 61.545 ;
        RECT 30.745 53.120 30.915 61.160 ;
        RECT 33.035 53.120 33.205 61.160 ;
        RECT 35.325 53.120 35.495 61.160 ;
        RECT 37.615 53.120 37.785 61.160 ;
        RECT 39.905 53.120 40.075 61.160 ;
        RECT 42.195 53.120 42.365 61.160 ;
        RECT 44.485 53.120 44.655 61.160 ;
        RECT 46.775 53.120 46.945 61.160 ;
        RECT 49.065 53.120 49.235 61.160 ;
        RECT 30.975 52.735 32.975 52.905 ;
        RECT 33.265 52.735 35.265 52.905 ;
        RECT 35.555 52.735 37.555 52.905 ;
        RECT 37.845 52.735 39.845 52.905 ;
        RECT 40.135 52.735 42.135 52.905 ;
        RECT 42.425 52.735 44.425 52.905 ;
        RECT 44.715 52.735 46.715 52.905 ;
        RECT 47.005 52.735 49.005 52.905 ;
        RECT 49.735 52.215 49.905 62.065 ;
        RECT 50.635 61.375 52.635 61.545 ;
        RECT 52.925 61.375 54.925 61.545 ;
        RECT 55.215 61.375 57.215 61.545 ;
        RECT 57.505 61.375 59.505 61.545 ;
        RECT 59.795 61.375 61.795 61.545 ;
        RECT 62.085 61.375 64.085 61.545 ;
        RECT 64.375 61.375 66.375 61.545 ;
        RECT 66.665 61.375 68.665 61.545 ;
        RECT 50.405 53.120 50.575 61.160 ;
        RECT 52.695 53.120 52.865 61.160 ;
        RECT 54.985 53.120 55.155 61.160 ;
        RECT 57.275 53.120 57.445 61.160 ;
        RECT 59.565 53.120 59.735 61.160 ;
        RECT 61.855 53.120 62.025 61.160 ;
        RECT 64.145 53.120 64.315 61.160 ;
        RECT 66.435 53.120 66.605 61.160 ;
        RECT 68.725 53.120 68.895 61.160 ;
        RECT 50.635 52.735 52.635 52.905 ;
        RECT 52.925 52.735 54.925 52.905 ;
        RECT 55.215 52.735 57.215 52.905 ;
        RECT 57.505 52.735 59.505 52.905 ;
        RECT 59.795 52.735 61.795 52.905 ;
        RECT 62.085 52.735 64.085 52.905 ;
        RECT 64.375 52.735 66.375 52.905 ;
        RECT 66.665 52.735 68.665 52.905 ;
        RECT 69.395 52.215 69.565 62.065 ;
        RECT 70.295 61.375 72.295 61.545 ;
        RECT 72.585 61.375 74.585 61.545 ;
        RECT 74.875 61.375 76.875 61.545 ;
        RECT 77.165 61.375 79.165 61.545 ;
        RECT 79.455 61.375 81.455 61.545 ;
        RECT 81.745 61.375 83.745 61.545 ;
        RECT 84.035 61.375 86.035 61.545 ;
        RECT 86.325 61.375 88.325 61.545 ;
        RECT 70.065 53.120 70.235 61.160 ;
        RECT 72.355 53.120 72.525 61.160 ;
        RECT 74.645 53.120 74.815 61.160 ;
        RECT 76.935 53.120 77.105 61.160 ;
        RECT 79.225 53.120 79.395 61.160 ;
        RECT 81.515 53.120 81.685 61.160 ;
        RECT 83.805 53.120 83.975 61.160 ;
        RECT 86.095 53.120 86.265 61.160 ;
        RECT 88.385 53.120 88.555 61.160 ;
        RECT 70.295 52.735 72.295 52.905 ;
        RECT 72.585 52.735 74.585 52.905 ;
        RECT 74.875 52.735 76.875 52.905 ;
        RECT 77.165 52.735 79.165 52.905 ;
        RECT 79.455 52.735 81.455 52.905 ;
        RECT 81.745 52.735 83.745 52.905 ;
        RECT 84.035 52.735 86.035 52.905 ;
        RECT 86.325 52.735 88.325 52.905 ;
        RECT 89.055 52.215 89.225 62.065 ;
        RECT 89.955 61.375 91.955 61.545 ;
        RECT 92.245 61.375 94.245 61.545 ;
        RECT 94.535 61.375 96.535 61.545 ;
        RECT 96.825 61.375 98.825 61.545 ;
        RECT 99.115 61.375 101.115 61.545 ;
        RECT 101.405 61.375 103.405 61.545 ;
        RECT 103.695 61.375 105.695 61.545 ;
        RECT 105.985 61.375 107.985 61.545 ;
        RECT 89.725 53.120 89.895 61.160 ;
        RECT 92.015 53.120 92.185 61.160 ;
        RECT 94.305 53.120 94.475 61.160 ;
        RECT 96.595 53.120 96.765 61.160 ;
        RECT 98.885 53.120 99.055 61.160 ;
        RECT 101.175 53.120 101.345 61.160 ;
        RECT 103.465 53.120 103.635 61.160 ;
        RECT 105.755 53.120 105.925 61.160 ;
        RECT 108.045 53.120 108.215 61.160 ;
        RECT 89.955 52.735 91.955 52.905 ;
        RECT 92.245 52.735 94.245 52.905 ;
        RECT 94.535 52.735 96.535 52.905 ;
        RECT 96.825 52.735 98.825 52.905 ;
        RECT 99.115 52.735 101.115 52.905 ;
        RECT 101.405 52.735 103.405 52.905 ;
        RECT 103.695 52.735 105.695 52.905 ;
        RECT 105.985 52.735 107.985 52.905 ;
        RECT 108.715 52.215 108.885 62.065 ;
        RECT 109.615 61.375 111.615 61.545 ;
        RECT 111.905 61.375 113.905 61.545 ;
        RECT 114.195 61.375 116.195 61.545 ;
        RECT 116.485 61.375 118.485 61.545 ;
        RECT 118.775 61.375 120.775 61.545 ;
        RECT 121.065 61.375 123.065 61.545 ;
        RECT 123.355 61.375 125.355 61.545 ;
        RECT 125.645 61.375 127.645 61.545 ;
        RECT 109.385 53.120 109.555 61.160 ;
        RECT 111.675 53.120 111.845 61.160 ;
        RECT 113.965 53.120 114.135 61.160 ;
        RECT 116.255 53.120 116.425 61.160 ;
        RECT 118.545 53.120 118.715 61.160 ;
        RECT 120.835 53.120 121.005 61.160 ;
        RECT 123.125 53.120 123.295 61.160 ;
        RECT 125.415 53.120 125.585 61.160 ;
        RECT 127.705 53.120 127.875 61.160 ;
        RECT 109.615 52.735 111.615 52.905 ;
        RECT 111.905 52.735 113.905 52.905 ;
        RECT 114.195 52.735 116.195 52.905 ;
        RECT 116.485 52.735 118.485 52.905 ;
        RECT 118.775 52.735 120.775 52.905 ;
        RECT 121.065 52.735 123.065 52.905 ;
        RECT 123.355 52.735 125.355 52.905 ;
        RECT 125.645 52.735 127.645 52.905 ;
        RECT 128.375 52.215 128.905 62.065 ;
        RECT 10.055 52.045 128.905 52.215 ;
        RECT 10.055 42.195 10.585 52.045 ;
        RECT 11.315 51.355 13.315 51.525 ;
        RECT 13.605 51.355 15.605 51.525 ;
        RECT 15.895 51.355 17.895 51.525 ;
        RECT 18.185 51.355 20.185 51.525 ;
        RECT 20.475 51.355 22.475 51.525 ;
        RECT 22.765 51.355 24.765 51.525 ;
        RECT 25.055 51.355 27.055 51.525 ;
        RECT 27.345 51.355 29.345 51.525 ;
        RECT 11.085 43.100 11.255 51.140 ;
        RECT 13.375 43.100 13.545 51.140 ;
        RECT 15.665 43.100 15.835 51.140 ;
        RECT 17.955 43.100 18.125 51.140 ;
        RECT 20.245 43.100 20.415 51.140 ;
        RECT 22.535 43.100 22.705 51.140 ;
        RECT 24.825 43.100 24.995 51.140 ;
        RECT 27.115 43.100 27.285 51.140 ;
        RECT 29.405 43.100 29.575 51.140 ;
        RECT 11.315 42.715 13.315 42.885 ;
        RECT 13.605 42.715 15.605 42.885 ;
        RECT 15.895 42.715 17.895 42.885 ;
        RECT 18.185 42.715 20.185 42.885 ;
        RECT 20.475 42.715 22.475 42.885 ;
        RECT 22.765 42.715 24.765 42.885 ;
        RECT 25.055 42.715 27.055 42.885 ;
        RECT 27.345 42.715 29.345 42.885 ;
        RECT 30.075 42.195 30.245 52.045 ;
        RECT 30.975 51.355 32.975 51.525 ;
        RECT 33.265 51.355 35.265 51.525 ;
        RECT 35.555 51.355 37.555 51.525 ;
        RECT 37.845 51.355 39.845 51.525 ;
        RECT 40.135 51.355 42.135 51.525 ;
        RECT 42.425 51.355 44.425 51.525 ;
        RECT 44.715 51.355 46.715 51.525 ;
        RECT 47.005 51.355 49.005 51.525 ;
        RECT 30.745 43.100 30.915 51.140 ;
        RECT 33.035 43.100 33.205 51.140 ;
        RECT 35.325 43.100 35.495 51.140 ;
        RECT 37.615 43.100 37.785 51.140 ;
        RECT 39.905 43.100 40.075 51.140 ;
        RECT 42.195 43.100 42.365 51.140 ;
        RECT 44.485 43.100 44.655 51.140 ;
        RECT 46.775 43.100 46.945 51.140 ;
        RECT 49.065 43.100 49.235 51.140 ;
        RECT 30.975 42.715 32.975 42.885 ;
        RECT 33.265 42.715 35.265 42.885 ;
        RECT 35.555 42.715 37.555 42.885 ;
        RECT 37.845 42.715 39.845 42.885 ;
        RECT 40.135 42.715 42.135 42.885 ;
        RECT 42.425 42.715 44.425 42.885 ;
        RECT 44.715 42.715 46.715 42.885 ;
        RECT 47.005 42.715 49.005 42.885 ;
        RECT 49.735 42.195 49.905 52.045 ;
        RECT 50.635 51.355 52.635 51.525 ;
        RECT 52.925 51.355 54.925 51.525 ;
        RECT 55.215 51.355 57.215 51.525 ;
        RECT 57.505 51.355 59.505 51.525 ;
        RECT 59.795 51.355 61.795 51.525 ;
        RECT 62.085 51.355 64.085 51.525 ;
        RECT 64.375 51.355 66.375 51.525 ;
        RECT 66.665 51.355 68.665 51.525 ;
        RECT 50.405 43.100 50.575 51.140 ;
        RECT 52.695 43.100 52.865 51.140 ;
        RECT 54.985 43.100 55.155 51.140 ;
        RECT 57.275 43.100 57.445 51.140 ;
        RECT 59.565 43.100 59.735 51.140 ;
        RECT 61.855 43.100 62.025 51.140 ;
        RECT 64.145 43.100 64.315 51.140 ;
        RECT 66.435 43.100 66.605 51.140 ;
        RECT 68.725 43.100 68.895 51.140 ;
        RECT 50.635 42.715 52.635 42.885 ;
        RECT 52.925 42.715 54.925 42.885 ;
        RECT 55.215 42.715 57.215 42.885 ;
        RECT 57.505 42.715 59.505 42.885 ;
        RECT 59.795 42.715 61.795 42.885 ;
        RECT 62.085 42.715 64.085 42.885 ;
        RECT 64.375 42.715 66.375 42.885 ;
        RECT 66.665 42.715 68.665 42.885 ;
        RECT 69.395 42.195 69.565 52.045 ;
        RECT 70.295 51.355 72.295 51.525 ;
        RECT 72.585 51.355 74.585 51.525 ;
        RECT 74.875 51.355 76.875 51.525 ;
        RECT 77.165 51.355 79.165 51.525 ;
        RECT 79.455 51.355 81.455 51.525 ;
        RECT 81.745 51.355 83.745 51.525 ;
        RECT 84.035 51.355 86.035 51.525 ;
        RECT 86.325 51.355 88.325 51.525 ;
        RECT 70.065 43.100 70.235 51.140 ;
        RECT 72.355 43.100 72.525 51.140 ;
        RECT 74.645 43.100 74.815 51.140 ;
        RECT 76.935 43.100 77.105 51.140 ;
        RECT 79.225 43.100 79.395 51.140 ;
        RECT 81.515 43.100 81.685 51.140 ;
        RECT 83.805 43.100 83.975 51.140 ;
        RECT 86.095 43.100 86.265 51.140 ;
        RECT 88.385 43.100 88.555 51.140 ;
        RECT 70.295 42.715 72.295 42.885 ;
        RECT 72.585 42.715 74.585 42.885 ;
        RECT 74.875 42.715 76.875 42.885 ;
        RECT 77.165 42.715 79.165 42.885 ;
        RECT 79.455 42.715 81.455 42.885 ;
        RECT 81.745 42.715 83.745 42.885 ;
        RECT 84.035 42.715 86.035 42.885 ;
        RECT 86.325 42.715 88.325 42.885 ;
        RECT 89.055 42.195 89.225 52.045 ;
        RECT 89.955 51.355 91.955 51.525 ;
        RECT 92.245 51.355 94.245 51.525 ;
        RECT 94.535 51.355 96.535 51.525 ;
        RECT 96.825 51.355 98.825 51.525 ;
        RECT 99.115 51.355 101.115 51.525 ;
        RECT 101.405 51.355 103.405 51.525 ;
        RECT 103.695 51.355 105.695 51.525 ;
        RECT 105.985 51.355 107.985 51.525 ;
        RECT 89.725 43.100 89.895 51.140 ;
        RECT 92.015 43.100 92.185 51.140 ;
        RECT 94.305 43.100 94.475 51.140 ;
        RECT 96.595 43.100 96.765 51.140 ;
        RECT 98.885 43.100 99.055 51.140 ;
        RECT 101.175 43.100 101.345 51.140 ;
        RECT 103.465 43.100 103.635 51.140 ;
        RECT 105.755 43.100 105.925 51.140 ;
        RECT 108.045 43.100 108.215 51.140 ;
        RECT 89.955 42.715 91.955 42.885 ;
        RECT 92.245 42.715 94.245 42.885 ;
        RECT 94.535 42.715 96.535 42.885 ;
        RECT 96.825 42.715 98.825 42.885 ;
        RECT 99.115 42.715 101.115 42.885 ;
        RECT 101.405 42.715 103.405 42.885 ;
        RECT 103.695 42.715 105.695 42.885 ;
        RECT 105.985 42.715 107.985 42.885 ;
        RECT 108.715 42.195 108.885 52.045 ;
        RECT 109.615 51.355 111.615 51.525 ;
        RECT 111.905 51.355 113.905 51.525 ;
        RECT 114.195 51.355 116.195 51.525 ;
        RECT 116.485 51.355 118.485 51.525 ;
        RECT 118.775 51.355 120.775 51.525 ;
        RECT 121.065 51.355 123.065 51.525 ;
        RECT 123.355 51.355 125.355 51.525 ;
        RECT 125.645 51.355 127.645 51.525 ;
        RECT 109.385 43.100 109.555 51.140 ;
        RECT 111.675 43.100 111.845 51.140 ;
        RECT 113.965 43.100 114.135 51.140 ;
        RECT 116.255 43.100 116.425 51.140 ;
        RECT 118.545 43.100 118.715 51.140 ;
        RECT 120.835 43.100 121.005 51.140 ;
        RECT 123.125 43.100 123.295 51.140 ;
        RECT 125.415 43.100 125.585 51.140 ;
        RECT 127.705 43.100 127.875 51.140 ;
        RECT 109.615 42.715 111.615 42.885 ;
        RECT 111.905 42.715 113.905 42.885 ;
        RECT 114.195 42.715 116.195 42.885 ;
        RECT 116.485 42.715 118.485 42.885 ;
        RECT 118.775 42.715 120.775 42.885 ;
        RECT 121.065 42.715 123.065 42.885 ;
        RECT 123.355 42.715 125.355 42.885 ;
        RECT 125.645 42.715 127.645 42.885 ;
        RECT 128.375 42.195 128.905 52.045 ;
        RECT 10.055 41.665 128.905 42.195 ;
        RECT 10.055 39.070 74.665 39.600 ;
        RECT 10.055 29.310 10.585 39.070 ;
        RECT 11.375 38.380 13.375 38.550 ;
        RECT 13.665 38.380 15.665 38.550 ;
        RECT 15.955 38.380 17.955 38.550 ;
        RECT 18.245 38.380 20.245 38.550 ;
        RECT 11.145 30.170 11.315 38.210 ;
        RECT 13.435 30.170 13.605 38.210 ;
        RECT 15.725 30.170 15.895 38.210 ;
        RECT 18.015 30.170 18.185 38.210 ;
        RECT 20.305 30.170 20.475 38.210 ;
        RECT 11.375 29.830 13.375 30.000 ;
        RECT 13.665 29.830 15.665 30.000 ;
        RECT 15.955 29.830 17.955 30.000 ;
        RECT 18.245 29.830 20.245 30.000 ;
        RECT 21.035 29.310 21.205 39.070 ;
        RECT 21.995 38.380 23.995 38.550 ;
        RECT 24.285 38.380 26.285 38.550 ;
        RECT 26.575 38.380 28.575 38.550 ;
        RECT 28.865 38.380 30.865 38.550 ;
        RECT 21.765 30.170 21.935 38.210 ;
        RECT 24.055 30.170 24.225 38.210 ;
        RECT 26.345 30.170 26.515 38.210 ;
        RECT 28.635 30.170 28.805 38.210 ;
        RECT 30.925 30.170 31.095 38.210 ;
        RECT 21.995 29.830 23.995 30.000 ;
        RECT 24.285 29.830 26.285 30.000 ;
        RECT 26.575 29.830 28.575 30.000 ;
        RECT 28.865 29.830 30.865 30.000 ;
        RECT 31.655 29.310 31.825 39.070 ;
        RECT 32.615 38.380 34.615 38.550 ;
        RECT 34.905 38.380 36.905 38.550 ;
        RECT 37.195 38.380 39.195 38.550 ;
        RECT 39.485 38.380 41.485 38.550 ;
        RECT 32.385 30.170 32.555 38.210 ;
        RECT 34.675 30.170 34.845 38.210 ;
        RECT 36.965 30.170 37.135 38.210 ;
        RECT 39.255 30.170 39.425 38.210 ;
        RECT 41.545 30.170 41.715 38.210 ;
        RECT 32.615 29.830 34.615 30.000 ;
        RECT 34.905 29.830 36.905 30.000 ;
        RECT 37.195 29.830 39.195 30.000 ;
        RECT 39.485 29.830 41.485 30.000 ;
        RECT 42.275 29.310 42.445 39.070 ;
        RECT 43.235 38.380 45.235 38.550 ;
        RECT 45.525 38.380 47.525 38.550 ;
        RECT 47.815 38.380 49.815 38.550 ;
        RECT 50.105 38.380 52.105 38.550 ;
        RECT 43.005 30.170 43.175 38.210 ;
        RECT 45.295 30.170 45.465 38.210 ;
        RECT 47.585 30.170 47.755 38.210 ;
        RECT 49.875 30.170 50.045 38.210 ;
        RECT 52.165 30.170 52.335 38.210 ;
        RECT 43.235 29.830 45.235 30.000 ;
        RECT 45.525 29.830 47.525 30.000 ;
        RECT 47.815 29.830 49.815 30.000 ;
        RECT 50.105 29.830 52.105 30.000 ;
        RECT 52.895 29.310 53.065 39.070 ;
        RECT 53.855 38.380 55.855 38.550 ;
        RECT 56.145 38.380 58.145 38.550 ;
        RECT 58.435 38.380 60.435 38.550 ;
        RECT 60.725 38.380 62.725 38.550 ;
        RECT 53.625 30.170 53.795 38.210 ;
        RECT 55.915 30.170 56.085 38.210 ;
        RECT 58.205 30.170 58.375 38.210 ;
        RECT 60.495 30.170 60.665 38.210 ;
        RECT 62.785 30.170 62.955 38.210 ;
        RECT 53.855 29.830 55.855 30.000 ;
        RECT 56.145 29.830 58.145 30.000 ;
        RECT 58.435 29.830 60.435 30.000 ;
        RECT 60.725 29.830 62.725 30.000 ;
        RECT 63.515 29.310 63.685 39.070 ;
        RECT 64.475 38.380 66.475 38.550 ;
        RECT 66.765 38.380 68.765 38.550 ;
        RECT 69.055 38.380 71.055 38.550 ;
        RECT 71.345 38.380 73.345 38.550 ;
        RECT 64.245 30.170 64.415 38.210 ;
        RECT 66.535 30.170 66.705 38.210 ;
        RECT 68.825 30.170 68.995 38.210 ;
        RECT 71.115 30.170 71.285 38.210 ;
        RECT 73.405 30.170 73.575 38.210 ;
        RECT 64.475 29.830 66.475 30.000 ;
        RECT 66.765 29.830 68.765 30.000 ;
        RECT 69.055 29.830 71.055 30.000 ;
        RECT 71.345 29.830 73.345 30.000 ;
        RECT 74.135 29.310 74.665 39.070 ;
        RECT 10.055 29.140 74.665 29.310 ;
        RECT 10.055 19.380 10.585 29.140 ;
        RECT 11.375 28.450 13.375 28.620 ;
        RECT 13.665 28.450 15.665 28.620 ;
        RECT 15.955 28.450 17.955 28.620 ;
        RECT 18.245 28.450 20.245 28.620 ;
        RECT 11.145 20.240 11.315 28.280 ;
        RECT 13.435 20.240 13.605 28.280 ;
        RECT 15.725 20.240 15.895 28.280 ;
        RECT 18.015 20.240 18.185 28.280 ;
        RECT 20.305 20.240 20.475 28.280 ;
        RECT 11.375 19.900 13.375 20.070 ;
        RECT 13.665 19.900 15.665 20.070 ;
        RECT 15.955 19.900 17.955 20.070 ;
        RECT 18.245 19.900 20.245 20.070 ;
        RECT 21.035 19.380 21.205 29.140 ;
        RECT 21.995 28.450 23.995 28.620 ;
        RECT 24.285 28.450 26.285 28.620 ;
        RECT 26.575 28.450 28.575 28.620 ;
        RECT 28.865 28.450 30.865 28.620 ;
        RECT 21.765 20.240 21.935 28.280 ;
        RECT 24.055 20.240 24.225 28.280 ;
        RECT 26.345 20.240 26.515 28.280 ;
        RECT 28.635 20.240 28.805 28.280 ;
        RECT 30.925 20.240 31.095 28.280 ;
        RECT 21.995 19.900 23.995 20.070 ;
        RECT 24.285 19.900 26.285 20.070 ;
        RECT 26.575 19.900 28.575 20.070 ;
        RECT 28.865 19.900 30.865 20.070 ;
        RECT 31.655 19.380 31.825 29.140 ;
        RECT 32.615 28.450 34.615 28.620 ;
        RECT 34.905 28.450 36.905 28.620 ;
        RECT 37.195 28.450 39.195 28.620 ;
        RECT 39.485 28.450 41.485 28.620 ;
        RECT 32.385 20.240 32.555 28.280 ;
        RECT 34.675 20.240 34.845 28.280 ;
        RECT 36.965 20.240 37.135 28.280 ;
        RECT 39.255 20.240 39.425 28.280 ;
        RECT 41.545 20.240 41.715 28.280 ;
        RECT 32.615 19.900 34.615 20.070 ;
        RECT 34.905 19.900 36.905 20.070 ;
        RECT 37.195 19.900 39.195 20.070 ;
        RECT 39.485 19.900 41.485 20.070 ;
        RECT 42.275 19.380 42.445 29.140 ;
        RECT 43.235 28.450 45.235 28.620 ;
        RECT 45.525 28.450 47.525 28.620 ;
        RECT 47.815 28.450 49.815 28.620 ;
        RECT 50.105 28.450 52.105 28.620 ;
        RECT 43.005 20.240 43.175 28.280 ;
        RECT 45.295 20.240 45.465 28.280 ;
        RECT 47.585 20.240 47.755 28.280 ;
        RECT 49.875 20.240 50.045 28.280 ;
        RECT 52.165 20.240 52.335 28.280 ;
        RECT 43.235 19.900 45.235 20.070 ;
        RECT 45.525 19.900 47.525 20.070 ;
        RECT 47.815 19.900 49.815 20.070 ;
        RECT 50.105 19.900 52.105 20.070 ;
        RECT 52.895 19.380 53.065 29.140 ;
        RECT 53.855 28.450 55.855 28.620 ;
        RECT 56.145 28.450 58.145 28.620 ;
        RECT 58.435 28.450 60.435 28.620 ;
        RECT 60.725 28.450 62.725 28.620 ;
        RECT 53.625 20.240 53.795 28.280 ;
        RECT 55.915 20.240 56.085 28.280 ;
        RECT 58.205 20.240 58.375 28.280 ;
        RECT 60.495 20.240 60.665 28.280 ;
        RECT 62.785 20.240 62.955 28.280 ;
        RECT 53.855 19.900 55.855 20.070 ;
        RECT 56.145 19.900 58.145 20.070 ;
        RECT 58.435 19.900 60.435 20.070 ;
        RECT 60.725 19.900 62.725 20.070 ;
        RECT 63.515 19.380 63.685 29.140 ;
        RECT 64.475 28.450 66.475 28.620 ;
        RECT 66.765 28.450 68.765 28.620 ;
        RECT 69.055 28.450 71.055 28.620 ;
        RECT 71.345 28.450 73.345 28.620 ;
        RECT 64.245 20.240 64.415 28.280 ;
        RECT 66.535 20.240 66.705 28.280 ;
        RECT 68.825 20.240 68.995 28.280 ;
        RECT 71.115 20.240 71.285 28.280 ;
        RECT 73.405 20.240 73.575 28.280 ;
        RECT 64.475 19.900 66.475 20.070 ;
        RECT 66.765 19.900 68.765 20.070 ;
        RECT 69.055 19.900 71.055 20.070 ;
        RECT 71.345 19.900 73.345 20.070 ;
        RECT 74.135 19.380 74.665 29.140 ;
        RECT 10.055 19.210 74.665 19.380 ;
        RECT 10.055 9.450 10.585 19.210 ;
        RECT 11.375 18.520 13.375 18.690 ;
        RECT 13.665 18.520 15.665 18.690 ;
        RECT 15.955 18.520 17.955 18.690 ;
        RECT 18.245 18.520 20.245 18.690 ;
        RECT 11.145 10.310 11.315 18.350 ;
        RECT 13.435 10.310 13.605 18.350 ;
        RECT 15.725 10.310 15.895 18.350 ;
        RECT 18.015 10.310 18.185 18.350 ;
        RECT 20.305 10.310 20.475 18.350 ;
        RECT 11.375 9.970 13.375 10.140 ;
        RECT 13.665 9.970 15.665 10.140 ;
        RECT 15.955 9.970 17.955 10.140 ;
        RECT 18.245 9.970 20.245 10.140 ;
        RECT 21.035 9.450 21.205 19.210 ;
        RECT 21.995 18.520 23.995 18.690 ;
        RECT 24.285 18.520 26.285 18.690 ;
        RECT 26.575 18.520 28.575 18.690 ;
        RECT 28.865 18.520 30.865 18.690 ;
        RECT 21.765 10.310 21.935 18.350 ;
        RECT 24.055 10.310 24.225 18.350 ;
        RECT 26.345 10.310 26.515 18.350 ;
        RECT 28.635 10.310 28.805 18.350 ;
        RECT 30.925 10.310 31.095 18.350 ;
        RECT 21.995 9.970 23.995 10.140 ;
        RECT 24.285 9.970 26.285 10.140 ;
        RECT 26.575 9.970 28.575 10.140 ;
        RECT 28.865 9.970 30.865 10.140 ;
        RECT 31.655 9.450 31.825 19.210 ;
        RECT 32.615 18.520 34.615 18.690 ;
        RECT 34.905 18.520 36.905 18.690 ;
        RECT 37.195 18.520 39.195 18.690 ;
        RECT 39.485 18.520 41.485 18.690 ;
        RECT 32.385 10.310 32.555 18.350 ;
        RECT 34.675 10.310 34.845 18.350 ;
        RECT 36.965 10.310 37.135 18.350 ;
        RECT 39.255 10.310 39.425 18.350 ;
        RECT 41.545 10.310 41.715 18.350 ;
        RECT 32.615 9.970 34.615 10.140 ;
        RECT 34.905 9.970 36.905 10.140 ;
        RECT 37.195 9.970 39.195 10.140 ;
        RECT 39.485 9.970 41.485 10.140 ;
        RECT 42.275 9.450 42.445 19.210 ;
        RECT 43.235 18.520 45.235 18.690 ;
        RECT 45.525 18.520 47.525 18.690 ;
        RECT 47.815 18.520 49.815 18.690 ;
        RECT 50.105 18.520 52.105 18.690 ;
        RECT 43.005 10.310 43.175 18.350 ;
        RECT 45.295 10.310 45.465 18.350 ;
        RECT 47.585 10.310 47.755 18.350 ;
        RECT 49.875 10.310 50.045 18.350 ;
        RECT 52.165 10.310 52.335 18.350 ;
        RECT 43.235 9.970 45.235 10.140 ;
        RECT 45.525 9.970 47.525 10.140 ;
        RECT 47.815 9.970 49.815 10.140 ;
        RECT 50.105 9.970 52.105 10.140 ;
        RECT 52.895 9.450 53.065 19.210 ;
        RECT 53.855 18.520 55.855 18.690 ;
        RECT 56.145 18.520 58.145 18.690 ;
        RECT 58.435 18.520 60.435 18.690 ;
        RECT 60.725 18.520 62.725 18.690 ;
        RECT 53.625 10.310 53.795 18.350 ;
        RECT 55.915 10.310 56.085 18.350 ;
        RECT 58.205 10.310 58.375 18.350 ;
        RECT 60.495 10.310 60.665 18.350 ;
        RECT 62.785 10.310 62.955 18.350 ;
        RECT 53.855 9.970 55.855 10.140 ;
        RECT 56.145 9.970 58.145 10.140 ;
        RECT 58.435 9.970 60.435 10.140 ;
        RECT 60.725 9.970 62.725 10.140 ;
        RECT 63.515 9.450 63.685 19.210 ;
        RECT 64.475 18.520 66.475 18.690 ;
        RECT 66.765 18.520 68.765 18.690 ;
        RECT 69.055 18.520 71.055 18.690 ;
        RECT 71.345 18.520 73.345 18.690 ;
        RECT 64.245 10.310 64.415 18.350 ;
        RECT 66.535 10.310 66.705 18.350 ;
        RECT 68.825 10.310 68.995 18.350 ;
        RECT 71.115 10.310 71.285 18.350 ;
        RECT 73.405 10.310 73.575 18.350 ;
        RECT 64.475 9.970 66.475 10.140 ;
        RECT 66.765 9.970 68.765 10.140 ;
        RECT 69.055 9.970 71.055 10.140 ;
        RECT 71.345 9.970 73.345 10.140 ;
        RECT 74.135 9.450 74.665 19.210 ;
        RECT 10.055 8.920 74.665 9.450 ;
        RECT 79.695 39.070 128.905 39.600 ;
        RECT 79.695 29.310 80.225 39.070 ;
        RECT 80.785 38.210 85.535 39.070 ;
        RECT 80.785 30.170 80.955 38.210 ;
        RECT 83.075 30.170 83.245 38.210 ;
        RECT 85.365 30.170 85.535 38.210 ;
        RECT 81.015 29.830 83.015 30.000 ;
        RECT 83.305 29.830 85.305 30.000 ;
        RECT 86.095 29.310 86.265 39.070 ;
        RECT 87.055 38.380 89.055 38.550 ;
        RECT 89.345 38.380 91.345 38.550 ;
        RECT 86.825 30.170 86.995 38.210 ;
        RECT 89.115 30.170 89.285 38.210 ;
        RECT 91.405 30.170 91.575 38.210 ;
        RECT 87.055 29.830 89.055 30.000 ;
        RECT 89.345 29.830 91.345 30.000 ;
        RECT 92.135 29.310 92.305 39.070 ;
        RECT 93.095 38.380 95.095 38.550 ;
        RECT 95.385 38.380 97.385 38.550 ;
        RECT 92.865 30.170 93.035 38.210 ;
        RECT 95.155 30.170 95.325 38.210 ;
        RECT 97.445 30.170 97.615 38.210 ;
        RECT 93.095 29.830 95.095 30.000 ;
        RECT 95.385 29.830 97.385 30.000 ;
        RECT 98.175 29.310 98.345 39.070 ;
        RECT 99.135 38.380 101.135 38.550 ;
        RECT 101.425 38.380 103.425 38.550 ;
        RECT 98.905 30.170 99.075 38.210 ;
        RECT 101.195 30.170 101.365 38.210 ;
        RECT 103.485 30.170 103.655 38.210 ;
        RECT 99.135 29.830 101.135 30.000 ;
        RECT 101.425 29.830 103.425 30.000 ;
        RECT 104.215 29.310 104.385 39.070 ;
        RECT 105.175 38.380 107.175 38.550 ;
        RECT 107.465 38.380 109.465 38.550 ;
        RECT 104.945 30.170 105.115 38.210 ;
        RECT 107.235 30.170 107.405 38.210 ;
        RECT 109.525 30.170 109.695 38.210 ;
        RECT 105.175 29.830 107.175 30.000 ;
        RECT 107.465 29.830 109.465 30.000 ;
        RECT 110.255 29.310 110.425 39.070 ;
        RECT 111.215 38.380 113.215 38.550 ;
        RECT 113.505 38.380 115.505 38.550 ;
        RECT 110.985 30.170 111.155 38.210 ;
        RECT 113.275 30.170 113.445 38.210 ;
        RECT 115.565 30.170 115.735 38.210 ;
        RECT 111.215 29.830 113.215 30.000 ;
        RECT 113.505 29.830 115.505 30.000 ;
        RECT 116.295 29.310 116.465 39.070 ;
        RECT 117.255 38.380 119.255 38.550 ;
        RECT 119.545 38.380 121.545 38.550 ;
        RECT 117.025 30.170 117.195 38.210 ;
        RECT 119.315 30.170 119.485 38.210 ;
        RECT 121.605 30.170 121.775 38.210 ;
        RECT 117.255 29.830 119.255 30.000 ;
        RECT 119.545 29.830 121.545 30.000 ;
        RECT 122.335 29.310 122.505 39.070 ;
        RECT 123.065 38.210 127.815 39.070 ;
        RECT 123.065 30.170 123.235 38.210 ;
        RECT 125.355 30.170 125.525 38.210 ;
        RECT 127.645 30.170 127.815 38.210 ;
        RECT 123.295 29.830 125.295 30.000 ;
        RECT 125.585 29.830 127.585 30.000 ;
        RECT 128.375 29.310 128.905 39.070 ;
        RECT 79.695 29.140 128.905 29.310 ;
        RECT 79.695 19.380 80.225 29.140 ;
        RECT 81.015 28.450 83.015 28.620 ;
        RECT 83.305 28.450 85.305 28.620 ;
        RECT 80.785 20.240 80.955 28.280 ;
        RECT 83.075 20.240 83.245 28.280 ;
        RECT 85.365 20.240 85.535 28.280 ;
        RECT 80.785 19.380 85.535 20.240 ;
        RECT 86.095 19.380 86.265 29.140 ;
        RECT 87.055 28.450 89.055 28.620 ;
        RECT 89.345 28.450 91.345 28.620 ;
        RECT 86.825 20.240 86.995 28.280 ;
        RECT 89.115 20.240 89.285 28.280 ;
        RECT 91.405 20.240 91.575 28.280 ;
        RECT 87.055 19.900 89.055 20.070 ;
        RECT 89.345 19.900 91.345 20.070 ;
        RECT 92.135 19.380 92.305 29.140 ;
        RECT 93.095 28.450 95.095 28.620 ;
        RECT 95.385 28.450 97.385 28.620 ;
        RECT 92.865 20.240 93.035 28.280 ;
        RECT 95.155 20.240 95.325 28.280 ;
        RECT 97.445 20.240 97.615 28.280 ;
        RECT 93.095 19.900 95.095 20.070 ;
        RECT 95.385 19.900 97.385 20.070 ;
        RECT 98.175 19.380 98.345 29.140 ;
        RECT 99.135 28.450 101.135 28.620 ;
        RECT 101.425 28.450 103.425 28.620 ;
        RECT 98.905 20.240 99.075 28.280 ;
        RECT 101.195 20.240 101.365 28.280 ;
        RECT 103.485 20.240 103.655 28.280 ;
        RECT 99.135 19.900 101.135 20.070 ;
        RECT 101.425 19.900 103.425 20.070 ;
        RECT 104.215 19.380 104.385 29.140 ;
        RECT 105.175 28.450 107.175 28.620 ;
        RECT 107.465 28.450 109.465 28.620 ;
        RECT 104.945 20.240 105.115 28.280 ;
        RECT 107.235 20.240 107.405 28.280 ;
        RECT 109.525 20.240 109.695 28.280 ;
        RECT 105.175 19.900 107.175 20.070 ;
        RECT 107.465 19.900 109.465 20.070 ;
        RECT 110.255 19.380 110.425 29.140 ;
        RECT 111.215 28.450 113.215 28.620 ;
        RECT 113.505 28.450 115.505 28.620 ;
        RECT 110.985 20.240 111.155 28.280 ;
        RECT 113.275 20.240 113.445 28.280 ;
        RECT 115.565 20.240 115.735 28.280 ;
        RECT 111.215 19.900 113.215 20.070 ;
        RECT 113.505 19.900 115.505 20.070 ;
        RECT 116.295 19.380 116.465 29.140 ;
        RECT 117.255 28.450 119.255 28.620 ;
        RECT 119.545 28.450 121.545 28.620 ;
        RECT 117.025 20.240 117.195 28.280 ;
        RECT 119.315 20.240 119.485 28.280 ;
        RECT 121.605 20.240 121.775 28.280 ;
        RECT 117.255 19.900 119.255 20.070 ;
        RECT 119.545 19.900 121.545 20.070 ;
        RECT 122.335 19.380 122.505 29.140 ;
        RECT 123.295 28.450 125.295 28.620 ;
        RECT 125.585 28.450 127.585 28.620 ;
        RECT 123.065 20.240 123.235 28.280 ;
        RECT 125.355 20.240 125.525 28.280 ;
        RECT 127.645 20.240 127.815 28.280 ;
        RECT 123.065 19.380 127.815 20.240 ;
        RECT 128.375 19.380 128.905 29.140 ;
        RECT 79.695 19.210 128.905 19.380 ;
        RECT 79.695 9.450 80.225 19.210 ;
        RECT 81.015 18.520 83.015 18.690 ;
        RECT 83.305 18.520 85.305 18.690 ;
        RECT 80.785 10.310 80.955 18.350 ;
        RECT 83.075 10.310 83.245 18.350 ;
        RECT 85.365 10.310 85.535 18.350 ;
        RECT 80.785 9.450 85.535 10.310 ;
        RECT 86.095 9.450 86.265 19.210 ;
        RECT 87.055 18.520 89.055 18.690 ;
        RECT 89.345 18.520 91.345 18.690 ;
        RECT 86.825 10.310 86.995 18.350 ;
        RECT 89.115 10.310 89.285 18.350 ;
        RECT 91.405 10.310 91.575 18.350 ;
        RECT 86.825 9.450 91.575 10.310 ;
        RECT 92.135 9.450 92.305 19.210 ;
        RECT 93.095 18.520 95.095 18.690 ;
        RECT 95.385 18.520 97.385 18.690 ;
        RECT 92.865 10.310 93.035 18.350 ;
        RECT 95.155 10.310 95.325 18.350 ;
        RECT 97.445 10.310 97.615 18.350 ;
        RECT 92.865 9.450 97.615 10.310 ;
        RECT 98.175 9.450 98.345 19.210 ;
        RECT 99.135 18.520 101.135 18.690 ;
        RECT 101.425 18.520 103.425 18.690 ;
        RECT 98.905 10.310 99.075 18.350 ;
        RECT 101.195 10.310 101.365 18.350 ;
        RECT 103.485 10.310 103.655 18.350 ;
        RECT 98.905 9.450 103.655 10.310 ;
        RECT 104.215 9.450 104.385 19.210 ;
        RECT 105.175 18.520 107.175 18.690 ;
        RECT 107.465 18.520 109.465 18.690 ;
        RECT 104.945 10.310 105.115 18.350 ;
        RECT 107.235 10.310 107.405 18.350 ;
        RECT 109.525 10.310 109.695 18.350 ;
        RECT 104.945 9.450 109.695 10.310 ;
        RECT 110.255 9.450 110.425 19.210 ;
        RECT 111.215 18.520 113.215 18.690 ;
        RECT 113.505 18.520 115.505 18.690 ;
        RECT 110.985 10.310 111.155 18.350 ;
        RECT 113.275 10.310 113.445 18.350 ;
        RECT 115.565 10.310 115.735 18.350 ;
        RECT 110.985 9.450 115.735 10.310 ;
        RECT 116.295 9.450 116.465 19.210 ;
        RECT 117.255 18.520 119.255 18.690 ;
        RECT 119.545 18.520 121.545 18.690 ;
        RECT 117.025 10.310 117.195 18.350 ;
        RECT 119.315 10.310 119.485 18.350 ;
        RECT 121.605 10.310 121.775 18.350 ;
        RECT 117.025 9.450 121.775 10.310 ;
        RECT 122.335 9.450 122.505 19.210 ;
        RECT 123.295 18.520 125.295 18.690 ;
        RECT 125.585 18.520 127.585 18.690 ;
        RECT 123.065 10.310 123.235 18.350 ;
        RECT 125.355 10.310 125.525 18.350 ;
        RECT 127.645 10.310 127.815 18.350 ;
        RECT 123.065 9.450 127.815 10.310 ;
        RECT 128.375 9.450 128.905 19.210 ;
        RECT 135.150 18.895 135.680 104.785 ;
        RECT 136.265 103.615 138.425 104.305 ;
        RECT 136.265 102.445 138.425 103.135 ;
        RECT 136.265 101.275 138.425 101.965 ;
        RECT 136.265 100.105 138.425 100.795 ;
        RECT 136.265 98.935 138.425 99.625 ;
        RECT 136.265 97.765 138.425 98.455 ;
        RECT 136.265 96.595 138.425 97.285 ;
        RECT 136.265 95.425 138.425 96.115 ;
        RECT 136.265 94.255 138.425 94.945 ;
        RECT 136.265 93.085 138.425 93.775 ;
        RECT 136.265 91.915 138.425 92.605 ;
        RECT 136.265 90.745 138.425 91.435 ;
        RECT 136.265 89.575 138.425 90.265 ;
        RECT 136.265 88.405 138.425 89.095 ;
        RECT 136.265 87.235 138.425 87.925 ;
        RECT 136.265 86.065 138.425 86.755 ;
        RECT 136.265 84.895 138.425 85.585 ;
        RECT 136.265 83.725 138.425 84.415 ;
        RECT 136.265 82.555 138.425 83.245 ;
        RECT 136.265 81.385 138.425 82.075 ;
        RECT 136.265 80.215 138.425 80.905 ;
        RECT 136.265 79.045 138.425 79.735 ;
        RECT 136.265 77.875 138.425 78.565 ;
        RECT 136.265 76.705 138.425 77.395 ;
        RECT 136.265 75.535 138.425 76.225 ;
        RECT 136.265 74.365 138.425 75.055 ;
        RECT 136.265 73.195 138.425 73.885 ;
        RECT 136.265 72.025 138.425 72.715 ;
        RECT 136.265 70.855 138.425 71.545 ;
        RECT 136.265 69.685 138.425 70.375 ;
        RECT 136.265 68.515 138.425 69.205 ;
        RECT 136.265 67.345 138.425 68.035 ;
        RECT 136.265 66.175 138.425 66.865 ;
        RECT 136.265 65.005 138.425 65.695 ;
        RECT 136.265 63.835 138.425 64.525 ;
        RECT 136.265 62.665 138.425 63.355 ;
        RECT 136.265 61.495 138.425 62.185 ;
        RECT 136.265 60.325 138.425 61.015 ;
        RECT 136.265 59.155 138.425 59.845 ;
        RECT 136.265 57.985 138.425 58.675 ;
        RECT 136.265 56.815 138.425 57.505 ;
        RECT 136.265 55.645 138.425 56.335 ;
        RECT 136.265 54.475 138.425 55.165 ;
        RECT 136.265 53.305 138.425 53.995 ;
        RECT 136.265 52.135 138.425 52.825 ;
        RECT 136.265 50.965 138.425 51.655 ;
        RECT 136.265 49.795 138.425 50.485 ;
        RECT 136.265 48.625 138.425 49.315 ;
        RECT 136.265 47.455 138.425 48.145 ;
        RECT 136.265 46.285 138.425 46.975 ;
        RECT 136.265 45.115 138.425 45.805 ;
        RECT 136.265 43.945 138.425 44.635 ;
        RECT 136.265 42.775 138.425 43.465 ;
        RECT 136.265 41.605 138.425 42.295 ;
        RECT 136.265 40.435 138.425 41.125 ;
        RECT 136.265 39.265 138.425 39.955 ;
        RECT 136.265 38.095 138.425 38.785 ;
        RECT 136.265 36.925 138.425 37.615 ;
        RECT 136.265 35.755 138.425 36.445 ;
        RECT 136.265 34.585 138.425 35.275 ;
        RECT 136.265 33.415 138.425 34.105 ;
        RECT 136.265 32.245 138.425 32.935 ;
        RECT 136.265 31.075 138.425 31.765 ;
        RECT 136.265 29.905 138.425 30.595 ;
        RECT 136.265 28.735 138.425 29.425 ;
        RECT 136.265 27.565 138.425 28.255 ;
        RECT 136.265 26.395 138.425 27.085 ;
        RECT 136.265 25.225 138.425 25.915 ;
        RECT 136.265 24.055 138.425 24.745 ;
        RECT 136.265 22.885 138.425 23.575 ;
        RECT 136.265 21.715 138.425 22.405 ;
        RECT 136.265 20.545 138.425 21.235 ;
        RECT 136.265 19.375 138.425 20.065 ;
        RECT 139.150 18.895 145.540 104.785 ;
        RECT 146.265 103.615 148.425 104.305 ;
        RECT 146.265 102.445 148.425 103.135 ;
        RECT 146.265 101.275 148.425 101.965 ;
        RECT 146.265 100.105 148.425 100.795 ;
        RECT 146.265 98.935 148.425 99.625 ;
        RECT 146.265 97.765 148.425 98.455 ;
        RECT 146.265 96.595 148.425 97.285 ;
        RECT 146.265 95.425 148.425 96.115 ;
        RECT 146.265 94.255 148.425 94.945 ;
        RECT 146.265 93.085 148.425 93.775 ;
        RECT 146.265 91.915 148.425 92.605 ;
        RECT 146.265 90.745 148.425 91.435 ;
        RECT 146.265 89.575 148.425 90.265 ;
        RECT 146.265 88.405 148.425 89.095 ;
        RECT 146.265 87.235 148.425 87.925 ;
        RECT 146.265 86.065 148.425 86.755 ;
        RECT 146.265 84.895 148.425 85.585 ;
        RECT 146.265 83.725 148.425 84.415 ;
        RECT 146.265 82.555 148.425 83.245 ;
        RECT 146.265 81.385 148.425 82.075 ;
        RECT 146.265 80.215 148.425 80.905 ;
        RECT 146.265 79.045 148.425 79.735 ;
        RECT 146.265 77.875 148.425 78.565 ;
        RECT 146.265 76.705 148.425 77.395 ;
        RECT 146.265 75.535 148.425 76.225 ;
        RECT 146.265 74.365 148.425 75.055 ;
        RECT 146.265 73.195 148.425 73.885 ;
        RECT 146.265 72.025 148.425 72.715 ;
        RECT 146.265 70.855 148.425 71.545 ;
        RECT 146.265 69.685 148.425 70.375 ;
        RECT 146.265 68.515 148.425 69.205 ;
        RECT 146.265 67.345 148.425 68.035 ;
        RECT 146.265 66.175 148.425 66.865 ;
        RECT 146.265 65.005 148.425 65.695 ;
        RECT 146.265 63.835 148.425 64.525 ;
        RECT 146.265 62.665 148.425 63.355 ;
        RECT 146.265 61.495 148.425 62.185 ;
        RECT 146.265 60.325 148.425 61.015 ;
        RECT 146.265 59.155 148.425 59.845 ;
        RECT 146.265 57.985 148.425 58.675 ;
        RECT 146.265 56.815 148.425 57.505 ;
        RECT 146.265 55.645 148.425 56.335 ;
        RECT 146.265 54.475 148.425 55.165 ;
        RECT 146.265 53.305 148.425 53.995 ;
        RECT 146.265 52.135 148.425 52.825 ;
        RECT 146.265 50.965 148.425 51.655 ;
        RECT 146.265 49.795 148.425 50.485 ;
        RECT 146.265 48.625 148.425 49.315 ;
        RECT 146.265 47.455 148.425 48.145 ;
        RECT 146.265 46.285 148.425 46.975 ;
        RECT 146.265 45.115 148.425 45.805 ;
        RECT 146.265 43.945 148.425 44.635 ;
        RECT 146.265 42.775 148.425 43.465 ;
        RECT 146.265 41.605 148.425 42.295 ;
        RECT 146.265 40.435 148.425 41.125 ;
        RECT 146.265 39.265 148.425 39.955 ;
        RECT 146.265 38.095 148.425 38.785 ;
        RECT 146.265 36.925 148.425 37.615 ;
        RECT 146.265 35.755 148.425 36.445 ;
        RECT 146.265 34.585 148.425 35.275 ;
        RECT 146.265 33.415 148.425 34.105 ;
        RECT 146.265 32.245 148.425 32.935 ;
        RECT 146.265 31.075 148.425 31.765 ;
        RECT 146.265 29.905 148.425 30.595 ;
        RECT 146.265 28.735 148.425 29.425 ;
        RECT 146.265 27.565 148.425 28.255 ;
        RECT 146.265 26.395 148.425 27.085 ;
        RECT 146.265 25.225 148.425 25.915 ;
        RECT 146.265 24.055 148.425 24.745 ;
        RECT 146.265 22.885 148.425 23.575 ;
        RECT 146.265 21.715 148.425 22.405 ;
        RECT 146.265 20.545 148.425 21.235 ;
        RECT 146.265 19.375 148.425 20.065 ;
        RECT 149.010 18.895 149.540 104.785 ;
        RECT 135.150 13.490 149.540 18.895 ;
        RECT 79.695 8.920 128.905 9.450 ;
        RECT 155.300 4.700 155.700 180.620 ;
        RECT 165.235 179.815 166.445 180.905 ;
        RECT 166.615 180.955 166.785 181.865 ;
        RECT 167.570 181.795 167.775 182.195 ;
        RECT 167.945 181.965 168.280 182.365 ;
        RECT 168.545 181.815 168.715 182.195 ;
        RECT 168.895 181.985 169.225 182.365 ;
        RECT 166.955 181.125 167.315 181.705 ;
        RECT 167.570 181.625 168.255 181.795 ;
        RECT 168.545 181.645 169.210 181.815 ;
        RECT 169.405 181.690 169.665 182.195 ;
        RECT 167.495 180.955 167.745 181.455 ;
        RECT 166.615 180.785 167.745 180.955 ;
        RECT 166.615 180.015 166.885 180.785 ;
        RECT 167.915 180.595 168.255 181.625 ;
        RECT 168.475 181.095 168.805 181.465 ;
        RECT 169.040 181.390 169.210 181.645 ;
        RECT 169.040 181.060 169.325 181.390 ;
        RECT 169.040 180.915 169.210 181.060 ;
        RECT 167.055 179.815 167.385 180.595 ;
        RECT 167.590 180.420 168.255 180.595 ;
        RECT 168.545 180.745 169.210 180.915 ;
        RECT 169.495 180.890 169.665 181.690 ;
        RECT 169.835 181.595 171.505 182.365 ;
        RECT 171.830 181.715 172.160 182.180 ;
        RECT 172.330 181.895 172.500 182.365 ;
        RECT 172.670 181.715 173.000 182.195 ;
        RECT 169.835 181.075 170.585 181.595 ;
        RECT 171.830 181.545 173.000 181.715 ;
        RECT 170.755 180.905 171.505 181.425 ;
        RECT 171.675 181.165 172.320 181.375 ;
        RECT 172.490 181.165 173.060 181.375 ;
        RECT 173.230 180.995 173.400 182.195 ;
        RECT 173.940 181.795 174.110 182.000 ;
        RECT 167.590 180.015 167.775 180.420 ;
        RECT 167.945 179.815 168.280 180.240 ;
        RECT 168.545 179.985 168.715 180.745 ;
        RECT 168.895 179.815 169.225 180.575 ;
        RECT 169.395 179.985 169.665 180.890 ;
        RECT 169.835 179.815 171.505 180.905 ;
        RECT 171.890 179.815 172.220 180.915 ;
        RECT 172.695 180.585 173.400 180.995 ;
        RECT 173.570 181.625 174.110 181.795 ;
        RECT 174.390 181.625 174.560 182.365 ;
        RECT 174.955 182.000 175.125 182.025 ;
        RECT 174.825 181.625 175.185 182.000 ;
        RECT 173.570 180.925 173.740 181.625 ;
        RECT 173.910 181.125 174.240 181.455 ;
        RECT 174.410 181.125 174.760 181.455 ;
        RECT 173.570 180.755 174.195 180.925 ;
        RECT 174.410 180.585 174.675 181.125 ;
        RECT 174.930 180.970 175.185 181.625 ;
        RECT 175.510 181.715 175.840 182.180 ;
        RECT 176.010 181.895 176.180 182.365 ;
        RECT 176.350 181.715 176.680 182.195 ;
        RECT 175.510 181.545 176.680 181.715 ;
        RECT 175.355 181.165 176.000 181.375 ;
        RECT 176.170 181.165 176.740 181.375 ;
        RECT 176.910 180.995 177.080 182.195 ;
        RECT 177.620 181.795 177.790 182.000 ;
        RECT 172.695 180.415 174.675 180.585 ;
        RECT 172.695 179.985 173.020 180.415 ;
        RECT 173.190 179.815 173.520 180.235 ;
        RECT 174.265 179.815 174.675 180.245 ;
        RECT 174.845 179.985 175.185 180.970 ;
        RECT 175.570 179.815 175.900 180.915 ;
        RECT 176.375 180.585 177.080 180.995 ;
        RECT 177.250 181.625 177.790 181.795 ;
        RECT 178.070 181.625 178.240 182.365 ;
        RECT 178.505 181.625 178.865 182.000 ;
        RECT 177.250 180.925 177.420 181.625 ;
        RECT 177.590 181.125 177.920 181.455 ;
        RECT 178.090 181.125 178.440 181.455 ;
        RECT 177.250 180.755 177.875 180.925 ;
        RECT 178.090 180.585 178.355 181.125 ;
        RECT 178.610 180.970 178.865 181.625 ;
        RECT 176.375 180.415 178.355 180.585 ;
        RECT 176.375 179.985 176.700 180.415 ;
        RECT 176.870 179.815 177.200 180.235 ;
        RECT 177.945 179.815 178.355 180.245 ;
        RECT 178.525 179.985 178.865 180.970 ;
        RECT 179.035 181.690 179.305 182.035 ;
        RECT 179.495 181.965 179.875 182.365 ;
        RECT 180.045 181.795 180.215 182.145 ;
        RECT 180.385 181.885 181.120 182.365 ;
        RECT 179.035 180.955 179.205 181.690 ;
        RECT 179.475 181.625 180.215 181.795 ;
        RECT 181.290 181.715 181.600 182.185 ;
        RECT 179.475 181.455 179.645 181.625 ;
        RECT 180.865 181.545 181.600 181.715 ;
        RECT 182.720 181.625 182.975 182.195 ;
        RECT 183.145 181.965 183.475 182.365 ;
        RECT 183.900 181.830 184.430 182.195 ;
        RECT 184.620 182.025 184.895 182.195 ;
        RECT 184.615 181.855 184.895 182.025 ;
        RECT 183.900 181.795 184.075 181.830 ;
        RECT 183.145 181.625 184.075 181.795 ;
        RECT 180.865 181.455 181.115 181.545 ;
        RECT 179.415 181.125 179.645 181.455 ;
        RECT 180.375 181.125 181.115 181.455 ;
        RECT 181.285 181.125 181.620 181.375 ;
        RECT 179.475 180.955 179.645 181.125 ;
        RECT 179.035 179.985 179.305 180.955 ;
        RECT 179.475 180.785 180.720 180.955 ;
        RECT 179.515 179.815 179.795 180.615 ;
        RECT 180.300 180.535 180.720 180.785 ;
        RECT 180.945 180.565 181.115 181.125 ;
        RECT 182.720 180.955 182.890 181.625 ;
        RECT 183.145 181.455 183.315 181.625 ;
        RECT 183.060 181.125 183.315 181.455 ;
        RECT 183.540 181.125 183.735 181.455 ;
        RECT 179.975 180.035 181.170 180.365 ;
        RECT 181.365 179.815 181.620 180.955 ;
        RECT 182.720 179.985 183.055 180.955 ;
        RECT 183.225 179.815 183.395 180.955 ;
        RECT 183.565 180.155 183.735 181.125 ;
        RECT 183.905 180.495 184.075 181.625 ;
        RECT 184.245 180.835 184.415 181.635 ;
        RECT 184.620 181.035 184.895 181.855 ;
        RECT 185.065 180.835 185.255 182.195 ;
        RECT 185.435 181.830 185.945 182.365 ;
        RECT 186.165 181.555 186.410 182.160 ;
        RECT 186.860 181.625 187.115 182.195 ;
        RECT 187.285 181.965 187.615 182.365 ;
        RECT 188.040 181.830 188.570 182.195 ;
        RECT 188.040 181.795 188.215 181.830 ;
        RECT 187.285 181.625 188.215 181.795 ;
        RECT 188.760 181.685 189.035 182.195 ;
        RECT 185.455 181.385 186.685 181.555 ;
        RECT 184.245 180.665 185.255 180.835 ;
        RECT 185.425 180.820 186.175 181.010 ;
        RECT 183.905 180.325 185.030 180.495 ;
        RECT 185.425 180.155 185.595 180.820 ;
        RECT 186.345 180.575 186.685 181.385 ;
        RECT 183.565 179.985 185.595 180.155 ;
        RECT 185.765 179.815 185.935 180.575 ;
        RECT 186.170 180.165 186.685 180.575 ;
        RECT 186.860 180.955 187.030 181.625 ;
        RECT 187.285 181.455 187.455 181.625 ;
        RECT 187.200 181.125 187.455 181.455 ;
        RECT 187.680 181.125 187.875 181.455 ;
        RECT 186.860 179.985 187.195 180.955 ;
        RECT 187.365 179.815 187.535 180.955 ;
        RECT 187.705 180.155 187.875 181.125 ;
        RECT 188.045 180.495 188.215 181.625 ;
        RECT 188.385 180.835 188.555 181.635 ;
        RECT 188.755 181.515 189.035 181.685 ;
        RECT 188.760 181.035 189.035 181.515 ;
        RECT 189.205 180.835 189.395 182.195 ;
        RECT 189.575 181.830 190.085 182.365 ;
        RECT 190.305 181.555 190.550 182.160 ;
        RECT 190.995 181.640 191.285 182.365 ;
        RECT 192.650 181.555 192.895 182.160 ;
        RECT 193.115 181.830 193.625 182.365 ;
        RECT 189.595 181.385 190.825 181.555 ;
        RECT 188.385 180.665 189.395 180.835 ;
        RECT 189.565 180.820 190.315 181.010 ;
        RECT 188.045 180.325 189.170 180.495 ;
        RECT 189.565 180.155 189.735 180.820 ;
        RECT 190.485 180.575 190.825 181.385 ;
        RECT 192.375 181.385 193.605 181.555 ;
        RECT 187.705 179.985 189.735 180.155 ;
        RECT 189.905 179.815 190.075 180.575 ;
        RECT 190.310 180.165 190.825 180.575 ;
        RECT 190.995 179.815 191.285 180.980 ;
        RECT 192.375 180.575 192.715 181.385 ;
        RECT 192.885 180.820 193.635 181.010 ;
        RECT 192.375 180.165 192.890 180.575 ;
        RECT 193.125 179.815 193.295 180.575 ;
        RECT 193.465 180.155 193.635 180.820 ;
        RECT 193.805 180.835 193.995 182.195 ;
        RECT 194.165 182.025 194.440 182.195 ;
        RECT 194.165 181.855 194.445 182.025 ;
        RECT 194.165 181.035 194.440 181.855 ;
        RECT 194.630 181.830 195.160 182.195 ;
        RECT 195.585 181.965 195.915 182.365 ;
        RECT 194.985 181.795 195.160 181.830 ;
        RECT 194.645 180.835 194.815 181.635 ;
        RECT 193.805 180.665 194.815 180.835 ;
        RECT 194.985 181.625 195.915 181.795 ;
        RECT 196.085 181.625 196.340 182.195 ;
        RECT 194.985 180.495 195.155 181.625 ;
        RECT 195.745 181.455 195.915 181.625 ;
        RECT 194.030 180.325 195.155 180.495 ;
        RECT 195.325 181.125 195.520 181.455 ;
        RECT 195.745 181.125 196.000 181.455 ;
        RECT 195.325 180.155 195.495 181.125 ;
        RECT 196.170 180.955 196.340 181.625 ;
        RECT 193.465 179.985 195.495 180.155 ;
        RECT 195.665 179.815 195.835 180.955 ;
        RECT 196.005 179.985 196.340 180.955 ;
        RECT 196.520 181.625 196.775 182.195 ;
        RECT 196.945 181.965 197.275 182.365 ;
        RECT 197.700 181.830 198.230 182.195 ;
        RECT 197.700 181.795 197.875 181.830 ;
        RECT 196.945 181.625 197.875 181.795 ;
        RECT 196.520 180.955 196.690 181.625 ;
        RECT 196.945 181.455 197.115 181.625 ;
        RECT 196.860 181.125 197.115 181.455 ;
        RECT 197.340 181.125 197.535 181.455 ;
        RECT 196.520 179.985 196.855 180.955 ;
        RECT 197.025 179.815 197.195 180.955 ;
        RECT 197.365 180.155 197.535 181.125 ;
        RECT 197.705 180.495 197.875 181.625 ;
        RECT 198.045 180.835 198.215 181.635 ;
        RECT 198.420 181.345 198.695 182.195 ;
        RECT 198.415 181.175 198.695 181.345 ;
        RECT 198.420 181.035 198.695 181.175 ;
        RECT 198.865 180.835 199.055 182.195 ;
        RECT 199.235 181.830 199.745 182.365 ;
        RECT 199.965 181.555 200.210 182.160 ;
        RECT 200.660 181.625 200.915 182.195 ;
        RECT 201.085 181.965 201.415 182.365 ;
        RECT 201.840 181.830 202.370 182.195 ;
        RECT 201.840 181.795 202.015 181.830 ;
        RECT 201.085 181.625 202.015 181.795 ;
        RECT 199.255 181.385 200.485 181.555 ;
        RECT 198.045 180.665 199.055 180.835 ;
        RECT 199.225 180.820 199.975 181.010 ;
        RECT 197.705 180.325 198.830 180.495 ;
        RECT 199.225 180.155 199.395 180.820 ;
        RECT 200.145 180.575 200.485 181.385 ;
        RECT 197.365 179.985 199.395 180.155 ;
        RECT 199.565 179.815 199.735 180.575 ;
        RECT 199.970 180.165 200.485 180.575 ;
        RECT 200.660 180.955 200.830 181.625 ;
        RECT 201.085 181.455 201.255 181.625 ;
        RECT 201.000 181.125 201.255 181.455 ;
        RECT 201.480 181.125 201.675 181.455 ;
        RECT 200.660 179.985 200.995 180.955 ;
        RECT 201.165 179.815 201.335 180.955 ;
        RECT 201.505 180.155 201.675 181.125 ;
        RECT 201.845 180.495 202.015 181.625 ;
        RECT 202.185 180.835 202.355 181.635 ;
        RECT 202.560 181.345 202.835 182.195 ;
        RECT 202.555 181.175 202.835 181.345 ;
        RECT 202.560 181.035 202.835 181.175 ;
        RECT 203.005 180.835 203.195 182.195 ;
        RECT 203.375 181.830 203.885 182.365 ;
        RECT 204.105 181.555 204.350 182.160 ;
        RECT 205.805 181.815 205.975 182.195 ;
        RECT 206.155 181.985 206.485 182.365 ;
        RECT 205.805 181.645 206.470 181.815 ;
        RECT 206.665 181.690 206.925 182.195 ;
        RECT 203.395 181.385 204.625 181.555 ;
        RECT 202.185 180.665 203.195 180.835 ;
        RECT 203.365 180.820 204.115 181.010 ;
        RECT 201.845 180.325 202.970 180.495 ;
        RECT 203.365 180.155 203.535 180.820 ;
        RECT 204.285 180.575 204.625 181.385 ;
        RECT 205.735 181.095 206.065 181.465 ;
        RECT 206.300 181.390 206.470 181.645 ;
        RECT 206.300 181.060 206.585 181.390 ;
        RECT 206.300 180.915 206.470 181.060 ;
        RECT 201.505 179.985 203.535 180.155 ;
        RECT 203.705 179.815 203.875 180.575 ;
        RECT 204.110 180.165 204.625 180.575 ;
        RECT 205.805 180.745 206.470 180.915 ;
        RECT 206.755 180.890 206.925 181.690 ;
        RECT 205.805 179.985 205.975 180.745 ;
        RECT 206.155 179.815 206.485 180.575 ;
        RECT 206.655 179.985 206.925 180.890 ;
        RECT 207.095 179.985 207.355 182.195 ;
        RECT 207.605 181.905 207.775 182.365 ;
        RECT 207.945 182.025 208.940 182.195 ;
        RECT 209.470 182.035 209.640 182.195 ;
        RECT 207.945 181.735 208.115 182.025 ;
        RECT 208.770 181.865 208.940 182.025 ;
        RECT 209.110 181.865 209.640 182.035 ;
        RECT 207.545 181.565 208.115 181.735 ;
        RECT 208.285 181.685 208.460 181.855 ;
        RECT 207.545 180.785 207.715 181.565 ;
        RECT 208.285 181.525 208.700 181.685 ;
        RECT 208.290 181.515 208.700 181.525 ;
        RECT 208.025 181.175 208.480 181.345 ;
        RECT 207.545 180.615 208.195 180.785 ;
        RECT 209.110 180.695 209.280 181.865 ;
        RECT 209.985 181.795 210.160 182.125 ;
        RECT 210.330 181.985 210.660 182.365 ;
        RECT 209.450 181.515 209.690 181.685 ;
        RECT 207.525 179.815 207.855 180.195 ;
        RECT 208.025 180.155 208.195 180.615 ;
        RECT 208.495 180.465 209.280 180.695 ;
        RECT 208.495 180.325 208.825 180.465 ;
        RECT 209.520 180.315 209.690 181.515 ;
        RECT 209.985 181.345 210.155 181.795 ;
        RECT 210.930 181.735 211.175 182.155 ;
        RECT 211.350 181.905 211.520 182.365 ;
        RECT 211.690 182.025 213.290 182.195 ;
        RECT 211.690 181.985 212.045 182.025 ;
        RECT 212.280 181.735 212.450 181.855 ;
        RECT 210.930 181.565 212.450 181.735 ;
        RECT 212.280 181.525 212.450 181.565 ;
        RECT 212.620 181.605 212.950 181.855 ;
        RECT 213.120 181.655 213.290 182.025 ;
        RECT 213.580 181.645 213.870 182.365 ;
        RECT 214.580 182.025 215.655 182.195 ;
        RECT 212.620 181.530 212.935 181.605 ;
        RECT 209.865 181.175 210.155 181.345 ;
        RECT 208.980 180.155 209.310 180.195 ;
        RECT 208.025 179.985 209.310 180.155 ;
        RECT 209.480 179.985 209.690 180.315 ;
        RECT 209.985 180.315 210.155 181.175 ;
        RECT 210.325 180.775 210.615 181.455 ;
        RECT 211.090 181.345 211.420 181.395 ;
        RECT 211.065 181.175 211.420 181.345 ;
        RECT 211.090 180.775 211.420 181.175 ;
        RECT 211.625 181.345 211.870 181.395 ;
        RECT 212.265 181.345 212.595 181.355 ;
        RECT 211.625 181.175 211.925 181.345 ;
        RECT 212.210 181.185 212.595 181.345 ;
        RECT 212.210 181.175 212.380 181.185 ;
        RECT 211.625 180.775 211.870 181.175 ;
        RECT 212.765 181.005 212.935 181.530 ;
        RECT 212.175 180.835 212.935 181.005 ;
        RECT 210.940 180.365 212.005 180.535 ;
        RECT 209.985 179.985 210.170 180.315 ;
        RECT 210.340 179.815 210.690 180.195 ;
        RECT 210.940 179.985 211.110 180.365 ;
        RECT 211.280 179.815 211.610 180.195 ;
        RECT 211.835 180.155 212.005 180.365 ;
        RECT 212.175 180.325 212.505 180.835 ;
        RECT 212.675 180.155 212.845 180.665 ;
        RECT 213.105 180.455 213.405 181.455 ;
        RECT 214.050 181.345 214.410 182.020 ;
        RECT 214.580 181.690 214.750 182.025 ;
        RECT 214.920 181.685 215.260 181.855 ;
        RECT 214.970 181.515 215.260 181.685 ;
        RECT 215.485 181.815 215.655 182.025 ;
        RECT 215.825 181.985 216.155 182.365 ;
        RECT 216.325 181.815 216.495 182.190 ;
        RECT 215.485 181.645 216.495 181.815 ;
        RECT 216.755 181.640 217.045 182.365 ;
        RECT 217.220 181.565 217.475 182.365 ;
        RECT 217.645 181.725 217.975 182.185 ;
        RECT 214.050 181.165 214.590 181.345 ;
        RECT 214.050 181.055 214.410 181.165 ;
        RECT 213.605 180.825 214.410 181.055 ;
        RECT 215.090 180.995 215.260 181.515 ;
        RECT 214.625 180.825 215.260 180.995 ;
        RECT 215.430 180.835 215.865 181.455 ;
        RECT 216.175 181.345 216.520 181.455 ;
        RECT 216.175 181.175 216.525 181.345 ;
        RECT 216.175 180.835 216.520 181.175 ;
        RECT 211.835 179.985 212.845 180.155 ;
        RECT 213.105 179.815 213.435 180.195 ;
        RECT 213.605 179.985 213.955 180.825 ;
        RECT 214.125 180.155 214.295 180.655 ;
        RECT 214.625 180.495 214.795 180.825 ;
        RECT 214.465 180.325 214.795 180.495 ;
        RECT 214.965 180.485 216.495 180.655 ;
        RECT 214.965 180.325 215.135 180.485 ;
        RECT 215.485 180.155 215.655 180.315 ;
        RECT 214.125 179.985 215.655 180.155 ;
        RECT 215.825 179.815 216.155 180.195 ;
        RECT 216.325 179.985 216.495 180.485 ;
        RECT 216.755 179.815 217.045 180.980 ;
        RECT 217.645 180.955 217.815 181.725 ;
        RECT 218.145 181.635 218.395 182.365 ;
        RECT 218.565 181.455 218.875 182.075 ;
        RECT 219.190 181.985 220.085 182.155 ;
        RECT 217.985 181.125 218.295 181.455 ;
        RECT 218.465 181.375 218.875 181.455 ;
        RECT 219.125 181.415 219.745 181.745 ;
        RECT 218.465 181.125 218.775 181.375 ;
        RECT 218.125 180.955 218.295 181.125 ;
        RECT 217.225 179.815 217.475 180.955 ;
        RECT 217.645 180.615 217.955 180.955 ;
        RECT 218.125 180.785 218.735 180.955 ;
        RECT 218.945 180.805 219.285 181.205 ;
        RECT 217.645 179.995 218.055 180.615 ;
        RECT 218.225 179.815 218.395 180.615 ;
        RECT 218.565 180.325 218.735 180.785 ;
        RECT 219.455 180.465 219.745 181.415 ;
        RECT 219.915 180.885 220.085 181.985 ;
        RECT 220.285 181.905 220.615 182.365 ;
        RECT 220.810 181.865 221.015 182.195 ;
        RECT 220.295 181.055 220.665 181.735 ;
        RECT 220.845 180.885 221.015 181.865 ;
        RECT 219.915 180.715 221.015 180.885 ;
        RECT 218.565 180.155 218.885 180.325 ;
        RECT 219.915 180.295 220.085 180.715 ;
        RECT 220.825 180.555 221.015 180.715 ;
        RECT 219.135 180.125 220.085 180.295 ;
        RECT 220.310 179.815 220.655 180.445 ;
        RECT 221.230 180.325 221.420 182.105 ;
        RECT 220.895 180.155 221.420 180.325 ;
        RECT 221.590 181.775 221.825 182.105 ;
        RECT 221.995 181.985 222.425 182.155 ;
        RECT 221.590 180.640 221.760 181.775 ;
        RECT 221.995 181.390 222.165 181.985 ;
        RECT 222.630 181.905 222.960 182.365 ;
        RECT 223.340 181.915 223.940 182.085 ;
        RECT 221.930 181.060 222.165 181.390 ;
        RECT 222.335 181.130 222.625 181.735 ;
        RECT 222.795 181.435 223.170 181.735 ;
        RECT 222.795 181.130 223.000 181.435 ;
        RECT 223.340 181.215 223.510 181.915 ;
        RECT 221.995 180.960 222.165 181.060 ;
        RECT 223.170 181.045 223.510 181.215 ;
        RECT 223.680 181.415 224.005 181.745 ;
        RECT 224.175 181.685 224.390 182.055 ;
        RECT 224.565 181.985 224.895 182.365 ;
        RECT 225.065 181.815 225.240 182.105 ;
        RECT 221.995 180.790 222.265 180.960 ;
        RECT 222.095 180.665 222.265 180.790 ;
        RECT 221.590 180.325 221.845 180.640 ;
        RECT 222.095 180.495 222.440 180.665 ;
        RECT 221.590 180.155 222.105 180.325 ;
        RECT 222.585 179.815 222.815 180.395 ;
        RECT 223.170 180.325 223.340 181.045 ;
        RECT 223.680 180.875 223.850 181.415 ;
        RECT 224.175 181.355 224.575 181.685 ;
        RECT 224.745 181.645 225.240 181.815 ;
        RECT 223.510 180.665 223.850 180.875 ;
        RECT 224.020 181.005 224.190 181.165 ;
        RECT 224.020 180.835 224.405 181.005 ;
        RECT 224.745 180.665 224.915 181.645 ;
        RECT 225.495 181.615 226.705 182.365 ;
        RECT 226.965 181.815 227.135 182.190 ;
        RECT 227.305 181.985 227.635 182.365 ;
        RECT 227.805 182.025 228.880 182.195 ;
        RECT 227.805 181.815 227.975 182.025 ;
        RECT 226.965 181.645 227.975 181.815 ;
        RECT 228.200 181.685 228.540 181.855 ;
        RECT 228.710 181.690 228.880 182.025 ;
        RECT 225.085 180.705 225.265 181.475 ;
        RECT 225.495 181.075 226.015 181.615 ;
        RECT 228.200 181.515 228.490 181.685 ;
        RECT 226.185 180.905 226.705 181.445 ;
        RECT 226.940 181.345 227.285 181.455 ;
        RECT 226.935 181.175 227.285 181.345 ;
        RECT 223.510 180.535 224.915 180.665 ;
        RECT 223.510 180.495 225.235 180.535 ;
        RECT 224.745 180.365 225.235 180.495 ;
        RECT 223.170 180.155 224.000 180.325 ;
        RECT 224.565 179.815 224.895 180.195 ;
        RECT 225.065 180.075 225.235 180.365 ;
        RECT 225.495 179.815 226.705 180.905 ;
        RECT 226.940 180.835 227.285 181.175 ;
        RECT 227.595 180.835 228.030 181.455 ;
        RECT 228.200 180.995 228.370 181.515 ;
        RECT 229.050 181.345 229.410 182.020 ;
        RECT 229.590 181.645 229.880 182.365 ;
        RECT 230.170 182.025 231.770 182.195 ;
        RECT 230.170 181.655 230.340 182.025 ;
        RECT 231.415 181.985 231.770 182.025 ;
        RECT 231.940 181.905 232.110 182.365 ;
        RECT 230.510 181.605 230.840 181.855 ;
        RECT 230.525 181.530 230.840 181.605 ;
        RECT 231.010 181.735 231.180 181.855 ;
        RECT 232.285 181.735 232.530 182.155 ;
        RECT 232.800 181.985 233.130 182.365 ;
        RECT 233.300 181.795 233.475 182.125 ;
        RECT 233.820 182.035 233.990 182.195 ;
        RECT 233.820 181.865 234.350 182.035 ;
        RECT 234.520 182.025 235.515 182.195 ;
        RECT 234.520 181.865 234.690 182.025 ;
        RECT 231.010 181.565 232.530 181.735 ;
        RECT 228.870 181.165 229.410 181.345 ;
        RECT 229.050 181.055 229.410 181.165 ;
        RECT 228.200 180.825 228.835 180.995 ;
        RECT 229.050 180.825 229.855 181.055 ;
        RECT 226.965 180.485 228.495 180.655 ;
        RECT 226.965 179.985 227.135 180.485 ;
        RECT 228.325 180.325 228.495 180.485 ;
        RECT 228.665 180.495 228.835 180.825 ;
        RECT 228.665 180.325 228.995 180.495 ;
        RECT 227.305 179.815 227.635 180.195 ;
        RECT 227.805 180.155 227.975 180.315 ;
        RECT 229.165 180.155 229.335 180.655 ;
        RECT 227.805 179.985 229.335 180.155 ;
        RECT 229.505 179.985 229.855 180.825 ;
        RECT 230.055 180.455 230.355 181.455 ;
        RECT 230.525 181.005 230.695 181.530 ;
        RECT 231.010 181.525 231.180 181.565 ;
        RECT 230.865 181.345 231.195 181.355 ;
        RECT 231.590 181.345 231.835 181.395 ;
        RECT 230.865 181.185 231.250 181.345 ;
        RECT 231.080 181.175 231.250 181.185 ;
        RECT 231.535 181.175 231.835 181.345 ;
        RECT 230.525 180.835 231.285 181.005 ;
        RECT 230.025 179.815 230.355 180.195 ;
        RECT 230.615 180.155 230.785 180.665 ;
        RECT 230.955 180.325 231.285 180.835 ;
        RECT 231.590 180.775 231.835 181.175 ;
        RECT 232.040 180.775 232.370 181.395 ;
        RECT 232.845 180.775 233.135 181.455 ;
        RECT 233.305 181.345 233.475 181.795 ;
        RECT 233.770 181.515 234.010 181.685 ;
        RECT 233.305 181.175 233.595 181.345 ;
        RECT 231.455 180.365 232.520 180.535 ;
        RECT 231.455 180.155 231.625 180.365 ;
        RECT 230.615 179.985 231.625 180.155 ;
        RECT 231.850 179.815 232.180 180.195 ;
        RECT 232.350 179.985 232.520 180.365 ;
        RECT 233.305 180.315 233.475 181.175 ;
        RECT 232.770 179.815 233.120 180.195 ;
        RECT 233.290 179.985 233.475 180.315 ;
        RECT 233.770 180.315 233.940 181.515 ;
        RECT 234.180 180.695 234.350 181.865 ;
        RECT 235.000 181.685 235.175 181.855 ;
        RECT 234.760 181.525 235.175 181.685 ;
        RECT 235.345 181.735 235.515 182.025 ;
        RECT 235.685 181.905 235.855 182.365 ;
        RECT 235.345 181.565 235.915 181.735 ;
        RECT 234.760 181.515 235.170 181.525 ;
        RECT 234.980 181.175 235.435 181.345 ;
        RECT 235.745 180.785 235.915 181.565 ;
        RECT 234.180 180.465 234.965 180.695 ;
        RECT 234.635 180.325 234.965 180.465 ;
        RECT 235.265 180.615 235.915 180.785 ;
        RECT 233.770 179.985 233.980 180.315 ;
        RECT 234.150 180.155 234.480 180.195 ;
        RECT 235.265 180.155 235.435 180.615 ;
        RECT 234.150 179.985 235.435 180.155 ;
        RECT 235.605 179.815 235.935 180.195 ;
        RECT 236.105 179.985 236.365 182.195 ;
        RECT 236.535 181.690 236.795 182.195 ;
        RECT 236.975 181.985 237.305 182.365 ;
        RECT 237.485 181.815 237.655 182.195 ;
        RECT 236.535 180.890 236.705 181.690 ;
        RECT 236.990 181.645 237.655 181.815 ;
        RECT 236.990 181.390 237.160 181.645 ;
        RECT 237.915 181.615 239.125 182.365 ;
        RECT 236.875 181.060 237.160 181.390 ;
        RECT 237.395 181.095 237.725 181.465 ;
        RECT 236.990 180.915 237.160 181.060 ;
        RECT 236.535 179.985 236.805 180.890 ;
        RECT 236.990 180.745 237.655 180.915 ;
        RECT 236.975 179.815 237.305 180.575 ;
        RECT 237.485 179.985 237.655 180.745 ;
        RECT 237.915 180.905 238.435 181.445 ;
        RECT 238.605 181.075 239.125 181.615 ;
        RECT 237.915 179.815 239.125 180.905 ;
        RECT 165.150 179.645 239.210 179.815 ;
        RECT 165.235 178.555 166.445 179.645 ;
        RECT 165.235 177.845 165.755 178.385 ;
        RECT 165.925 178.015 166.445 178.555 ;
        RECT 167.625 178.715 167.795 179.475 ;
        RECT 167.975 178.885 168.305 179.645 ;
        RECT 167.625 178.545 168.290 178.715 ;
        RECT 168.475 178.570 168.745 179.475 ;
        RECT 168.120 178.400 168.290 178.545 ;
        RECT 167.555 177.995 167.885 178.365 ;
        RECT 168.120 178.070 168.405 178.400 ;
        RECT 165.235 177.095 166.445 177.845 ;
        RECT 168.120 177.815 168.290 178.070 ;
        RECT 167.625 177.645 168.290 177.815 ;
        RECT 168.575 177.770 168.745 178.570 ;
        RECT 167.625 177.265 167.795 177.645 ;
        RECT 167.975 177.095 168.305 177.475 ;
        RECT 168.485 177.265 168.745 177.770 ;
        RECT 168.915 178.675 169.185 179.445 ;
        RECT 169.355 178.865 169.685 179.645 ;
        RECT 169.890 179.040 170.075 179.445 ;
        RECT 170.245 179.220 170.580 179.645 ;
        RECT 169.890 178.865 170.555 179.040 ;
        RECT 168.915 178.505 170.045 178.675 ;
        RECT 168.915 177.595 169.085 178.505 ;
        RECT 169.255 177.755 169.615 178.335 ;
        RECT 169.795 178.005 170.045 178.505 ;
        RECT 170.215 177.835 170.555 178.865 ;
        RECT 170.970 178.545 171.300 179.645 ;
        RECT 171.775 179.045 172.100 179.475 ;
        RECT 172.270 179.225 172.600 179.645 ;
        RECT 173.345 179.215 173.755 179.645 ;
        RECT 171.775 178.875 173.755 179.045 ;
        RECT 171.775 178.465 172.480 178.875 ;
        RECT 170.755 178.085 171.400 178.295 ;
        RECT 171.570 178.085 172.140 178.295 ;
        RECT 169.870 177.665 170.555 177.835 ;
        RECT 170.910 177.745 172.080 177.915 ;
        RECT 168.915 177.265 169.175 177.595 ;
        RECT 169.385 177.095 169.660 177.575 ;
        RECT 169.870 177.265 170.075 177.665 ;
        RECT 170.245 177.095 170.580 177.495 ;
        RECT 170.910 177.280 171.240 177.745 ;
        RECT 171.410 177.095 171.580 177.565 ;
        RECT 171.750 177.265 172.080 177.745 ;
        RECT 172.310 177.265 172.480 178.465 ;
        RECT 172.650 178.535 173.275 178.705 ;
        RECT 172.650 177.835 172.820 178.535 ;
        RECT 173.490 178.335 173.755 178.875 ;
        RECT 173.925 178.490 174.265 179.475 ;
        RECT 174.490 178.775 174.775 179.645 ;
        RECT 174.945 179.015 175.205 179.475 ;
        RECT 175.380 179.185 175.635 179.645 ;
        RECT 175.805 179.015 176.065 179.475 ;
        RECT 174.945 178.845 176.065 179.015 ;
        RECT 176.235 178.845 176.545 179.645 ;
        RECT 174.945 178.595 175.205 178.845 ;
        RECT 176.715 178.675 177.025 179.475 ;
        RECT 172.990 178.005 173.320 178.335 ;
        RECT 173.490 178.005 173.840 178.335 ;
        RECT 174.010 177.835 174.265 178.490 ;
        RECT 172.650 177.665 173.190 177.835 ;
        RECT 173.020 177.460 173.190 177.665 ;
        RECT 173.470 177.095 173.640 177.835 ;
        RECT 173.905 177.460 174.265 177.835 ;
        RECT 174.450 178.425 175.205 178.595 ;
        RECT 175.995 178.505 177.025 178.675 ;
        RECT 174.450 177.915 174.855 178.425 ;
        RECT 175.995 178.255 176.165 178.505 ;
        RECT 175.025 178.085 176.165 178.255 ;
        RECT 174.450 177.745 176.100 177.915 ;
        RECT 176.335 177.765 176.685 178.335 ;
        RECT 174.495 177.095 174.775 177.575 ;
        RECT 174.945 177.355 175.205 177.745 ;
        RECT 175.380 177.095 175.635 177.575 ;
        RECT 175.805 177.355 176.100 177.745 ;
        RECT 176.855 177.595 177.025 178.505 ;
        RECT 178.115 178.480 178.405 179.645 ;
        RECT 178.575 178.505 178.845 179.475 ;
        RECT 179.055 178.845 179.335 179.645 ;
        RECT 179.515 179.095 180.710 179.425 ;
        RECT 179.840 178.675 180.260 178.925 ;
        RECT 179.015 178.505 180.260 178.675 ;
        RECT 176.280 177.095 176.555 177.575 ;
        RECT 176.725 177.265 177.025 177.595 ;
        RECT 178.115 177.095 178.405 177.820 ;
        RECT 178.575 177.770 178.745 178.505 ;
        RECT 179.015 178.335 179.185 178.505 ;
        RECT 180.485 178.335 180.655 178.895 ;
        RECT 180.905 178.505 181.160 179.645 ;
        RECT 181.425 178.715 181.595 179.475 ;
        RECT 181.775 178.885 182.105 179.645 ;
        RECT 181.425 178.545 182.090 178.715 ;
        RECT 182.275 178.570 182.545 179.475 ;
        RECT 181.920 178.400 182.090 178.545 ;
        RECT 178.955 178.005 179.185 178.335 ;
        RECT 179.915 178.005 180.655 178.335 ;
        RECT 180.825 178.085 181.160 178.335 ;
        RECT 179.015 177.835 179.185 178.005 ;
        RECT 180.405 177.915 180.655 178.005 ;
        RECT 181.355 177.995 181.685 178.365 ;
        RECT 181.920 178.070 182.205 178.400 ;
        RECT 178.575 177.425 178.845 177.770 ;
        RECT 179.015 177.665 179.755 177.835 ;
        RECT 180.405 177.745 181.140 177.915 ;
        RECT 181.920 177.815 182.090 178.070 ;
        RECT 179.035 177.095 179.415 177.495 ;
        RECT 179.585 177.315 179.755 177.665 ;
        RECT 179.925 177.095 180.660 177.575 ;
        RECT 180.830 177.275 181.140 177.745 ;
        RECT 181.425 177.645 182.090 177.815 ;
        RECT 182.375 177.770 182.545 178.570 ;
        RECT 181.425 177.265 181.595 177.645 ;
        RECT 181.775 177.095 182.105 177.475 ;
        RECT 182.285 177.265 182.545 177.770 ;
        RECT 182.720 178.505 183.055 179.475 ;
        RECT 183.225 178.505 183.395 179.645 ;
        RECT 183.565 179.305 185.595 179.475 ;
        RECT 182.720 177.835 182.890 178.505 ;
        RECT 183.565 178.335 183.735 179.305 ;
        RECT 183.060 178.005 183.315 178.335 ;
        RECT 183.540 178.005 183.735 178.335 ;
        RECT 183.905 178.965 185.030 179.135 ;
        RECT 183.145 177.835 183.315 178.005 ;
        RECT 183.905 177.835 184.075 178.965 ;
        RECT 182.720 177.265 182.975 177.835 ;
        RECT 183.145 177.665 184.075 177.835 ;
        RECT 184.245 178.625 185.255 178.795 ;
        RECT 184.245 177.825 184.415 178.625 ;
        RECT 183.900 177.630 184.075 177.665 ;
        RECT 183.145 177.095 183.475 177.495 ;
        RECT 183.900 177.265 184.430 177.630 ;
        RECT 184.620 177.605 184.895 178.425 ;
        RECT 184.615 177.435 184.895 177.605 ;
        RECT 184.620 177.265 184.895 177.435 ;
        RECT 185.065 177.265 185.255 178.625 ;
        RECT 185.425 178.640 185.595 179.305 ;
        RECT 185.765 178.885 185.935 179.645 ;
        RECT 186.170 178.885 186.685 179.295 ;
        RECT 185.425 178.450 186.175 178.640 ;
        RECT 186.345 178.075 186.685 178.885 ;
        RECT 185.455 177.905 186.685 178.075 ;
        RECT 186.855 178.570 187.125 179.475 ;
        RECT 187.295 178.885 187.625 179.645 ;
        RECT 187.805 178.715 187.975 179.475 ;
        RECT 185.435 177.095 185.945 177.630 ;
        RECT 186.165 177.300 186.410 177.905 ;
        RECT 186.855 177.770 187.025 178.570 ;
        RECT 187.310 178.545 187.975 178.715 ;
        RECT 188.235 178.570 188.505 179.475 ;
        RECT 188.675 178.885 189.005 179.645 ;
        RECT 189.185 178.715 189.355 179.475 ;
        RECT 187.310 178.400 187.480 178.545 ;
        RECT 187.195 178.070 187.480 178.400 ;
        RECT 187.310 177.815 187.480 178.070 ;
        RECT 187.715 177.995 188.045 178.365 ;
        RECT 186.855 177.265 187.115 177.770 ;
        RECT 187.310 177.645 187.975 177.815 ;
        RECT 187.295 177.095 187.625 177.475 ;
        RECT 187.805 177.265 187.975 177.645 ;
        RECT 188.235 177.770 188.405 178.570 ;
        RECT 188.690 178.545 189.355 178.715 ;
        RECT 189.705 178.715 189.875 179.475 ;
        RECT 190.055 178.885 190.385 179.645 ;
        RECT 189.705 178.545 190.370 178.715 ;
        RECT 190.555 178.570 190.825 179.475 ;
        RECT 188.690 178.400 188.860 178.545 ;
        RECT 188.575 178.070 188.860 178.400 ;
        RECT 190.200 178.400 190.370 178.545 ;
        RECT 188.690 177.815 188.860 178.070 ;
        RECT 189.095 177.995 189.425 178.365 ;
        RECT 189.635 177.995 189.965 178.365 ;
        RECT 190.200 178.070 190.485 178.400 ;
        RECT 190.200 177.815 190.370 178.070 ;
        RECT 188.235 177.265 188.495 177.770 ;
        RECT 188.690 177.645 189.355 177.815 ;
        RECT 188.675 177.095 189.005 177.475 ;
        RECT 189.185 177.265 189.355 177.645 ;
        RECT 189.705 177.645 190.370 177.815 ;
        RECT 190.655 177.770 190.825 178.570 ;
        RECT 190.995 178.480 191.285 179.645 ;
        RECT 192.005 178.715 192.175 179.475 ;
        RECT 192.355 178.885 192.685 179.645 ;
        RECT 192.005 178.545 192.670 178.715 ;
        RECT 192.855 178.570 193.125 179.475 ;
        RECT 192.500 178.400 192.670 178.545 ;
        RECT 191.935 177.995 192.265 178.365 ;
        RECT 192.500 178.070 192.785 178.400 ;
        RECT 189.705 177.265 189.875 177.645 ;
        RECT 190.055 177.095 190.385 177.475 ;
        RECT 190.565 177.265 190.825 177.770 ;
        RECT 190.995 177.095 191.285 177.820 ;
        RECT 192.500 177.815 192.670 178.070 ;
        RECT 192.005 177.645 192.670 177.815 ;
        RECT 192.955 177.770 193.125 178.570 ;
        RECT 192.005 177.265 192.175 177.645 ;
        RECT 192.355 177.095 192.685 177.475 ;
        RECT 192.865 177.265 193.125 177.770 ;
        RECT 193.295 178.570 193.565 179.475 ;
        RECT 193.735 178.885 194.065 179.645 ;
        RECT 194.245 178.715 194.415 179.475 ;
        RECT 193.295 177.770 193.465 178.570 ;
        RECT 193.750 178.545 194.415 178.715 ;
        RECT 194.765 178.715 194.935 179.475 ;
        RECT 195.115 178.885 195.445 179.645 ;
        RECT 194.765 178.545 195.430 178.715 ;
        RECT 195.615 178.570 195.885 179.475 ;
        RECT 193.750 178.400 193.920 178.545 ;
        RECT 193.635 178.070 193.920 178.400 ;
        RECT 195.260 178.400 195.430 178.545 ;
        RECT 193.750 177.815 193.920 178.070 ;
        RECT 194.155 177.995 194.485 178.365 ;
        RECT 194.695 177.995 195.025 178.365 ;
        RECT 195.260 178.070 195.545 178.400 ;
        RECT 195.260 177.815 195.430 178.070 ;
        RECT 193.295 177.265 193.555 177.770 ;
        RECT 193.750 177.645 194.415 177.815 ;
        RECT 193.735 177.095 194.065 177.475 ;
        RECT 194.245 177.265 194.415 177.645 ;
        RECT 194.765 177.645 195.430 177.815 ;
        RECT 195.715 177.770 195.885 178.570 ;
        RECT 194.765 177.265 194.935 177.645 ;
        RECT 195.115 177.095 195.445 177.475 ;
        RECT 195.625 177.265 195.885 177.770 ;
        RECT 196.060 178.505 196.395 179.475 ;
        RECT 196.565 178.505 196.735 179.645 ;
        RECT 196.905 179.305 198.935 179.475 ;
        RECT 196.060 177.835 196.230 178.505 ;
        RECT 196.905 178.335 197.075 179.305 ;
        RECT 196.400 178.005 196.655 178.335 ;
        RECT 196.880 178.005 197.075 178.335 ;
        RECT 197.245 178.965 198.370 179.135 ;
        RECT 196.485 177.835 196.655 178.005 ;
        RECT 197.245 177.835 197.415 178.965 ;
        RECT 196.060 177.265 196.315 177.835 ;
        RECT 196.485 177.665 197.415 177.835 ;
        RECT 197.585 178.625 198.595 178.795 ;
        RECT 197.585 177.825 197.755 178.625 ;
        RECT 197.240 177.630 197.415 177.665 ;
        RECT 196.485 177.095 196.815 177.495 ;
        RECT 197.240 177.265 197.770 177.630 ;
        RECT 197.960 177.605 198.235 178.425 ;
        RECT 197.955 177.435 198.235 177.605 ;
        RECT 197.960 177.265 198.235 177.435 ;
        RECT 198.405 177.265 198.595 178.625 ;
        RECT 198.765 178.640 198.935 179.305 ;
        RECT 199.105 178.885 199.275 179.645 ;
        RECT 199.510 178.885 200.025 179.295 ;
        RECT 198.765 178.450 199.515 178.640 ;
        RECT 199.685 178.075 200.025 178.885 ;
        RECT 201.205 178.715 201.375 179.475 ;
        RECT 201.555 178.885 201.885 179.645 ;
        RECT 201.205 178.545 201.870 178.715 ;
        RECT 202.055 178.570 202.325 179.475 ;
        RECT 201.700 178.400 201.870 178.545 ;
        RECT 198.795 177.905 200.025 178.075 ;
        RECT 201.135 177.995 201.465 178.365 ;
        RECT 201.700 178.070 201.985 178.400 ;
        RECT 198.775 177.095 199.285 177.630 ;
        RECT 199.505 177.300 199.750 177.905 ;
        RECT 201.700 177.815 201.870 178.070 ;
        RECT 201.205 177.645 201.870 177.815 ;
        RECT 202.155 177.770 202.325 178.570 ;
        RECT 202.585 178.715 202.755 179.475 ;
        RECT 202.935 178.885 203.265 179.645 ;
        RECT 202.585 178.545 203.250 178.715 ;
        RECT 203.435 178.570 203.705 179.475 ;
        RECT 203.080 178.400 203.250 178.545 ;
        RECT 202.515 177.995 202.845 178.365 ;
        RECT 203.080 178.070 203.365 178.400 ;
        RECT 203.080 177.815 203.250 178.070 ;
        RECT 201.205 177.265 201.375 177.645 ;
        RECT 201.555 177.095 201.885 177.475 ;
        RECT 202.065 177.265 202.325 177.770 ;
        RECT 202.585 177.645 203.250 177.815 ;
        RECT 203.535 177.770 203.705 178.570 ;
        RECT 203.875 178.480 204.165 179.645 ;
        RECT 204.885 178.715 205.055 179.475 ;
        RECT 205.235 178.885 205.565 179.645 ;
        RECT 204.885 178.545 205.550 178.715 ;
        RECT 205.735 178.570 206.005 179.475 ;
        RECT 205.380 178.400 205.550 178.545 ;
        RECT 204.815 177.995 205.145 178.365 ;
        RECT 205.380 178.070 205.665 178.400 ;
        RECT 202.585 177.265 202.755 177.645 ;
        RECT 202.935 177.095 203.265 177.475 ;
        RECT 203.445 177.265 203.705 177.770 ;
        RECT 203.875 177.095 204.165 177.820 ;
        RECT 205.380 177.815 205.550 178.070 ;
        RECT 204.885 177.645 205.550 177.815 ;
        RECT 205.835 177.770 206.005 178.570 ;
        RECT 204.885 177.265 205.055 177.645 ;
        RECT 205.235 177.095 205.565 177.475 ;
        RECT 205.745 177.265 206.005 177.770 ;
        RECT 207.095 177.265 207.355 179.475 ;
        RECT 207.525 179.265 207.855 179.645 ;
        RECT 208.025 179.305 209.310 179.475 ;
        RECT 208.025 178.845 208.195 179.305 ;
        RECT 208.980 179.265 209.310 179.305 ;
        RECT 209.480 179.145 209.690 179.475 ;
        RECT 207.545 178.675 208.195 178.845 ;
        RECT 208.495 178.995 208.825 179.135 ;
        RECT 208.495 178.765 209.280 178.995 ;
        RECT 207.545 177.895 207.715 178.675 ;
        RECT 208.025 178.115 208.480 178.285 ;
        RECT 208.290 177.935 208.700 177.945 ;
        RECT 207.545 177.725 208.115 177.895 ;
        RECT 207.605 177.095 207.775 177.555 ;
        RECT 207.945 177.435 208.115 177.725 ;
        RECT 208.285 177.775 208.700 177.935 ;
        RECT 208.285 177.605 208.460 177.775 ;
        RECT 209.110 177.595 209.280 178.765 ;
        RECT 209.520 177.945 209.690 179.145 ;
        RECT 209.985 179.145 210.170 179.475 ;
        RECT 210.340 179.265 210.690 179.645 ;
        RECT 209.985 178.285 210.155 179.145 ;
        RECT 210.940 179.095 211.110 179.475 ;
        RECT 211.280 179.265 211.610 179.645 ;
        RECT 211.835 179.305 212.845 179.475 ;
        RECT 211.835 179.095 212.005 179.305 ;
        RECT 210.940 178.925 212.005 179.095 ;
        RECT 209.865 178.115 210.155 178.285 ;
        RECT 209.450 177.775 209.690 177.945 ;
        RECT 209.985 177.665 210.155 178.115 ;
        RECT 210.325 178.005 210.615 178.685 ;
        RECT 211.090 178.065 211.420 178.685 ;
        RECT 211.625 178.285 211.870 178.685 ;
        RECT 212.175 178.625 212.505 179.135 ;
        RECT 212.675 178.795 212.845 179.305 ;
        RECT 213.105 179.265 213.435 179.645 ;
        RECT 212.175 178.455 212.935 178.625 ;
        RECT 211.625 178.115 211.925 178.285 ;
        RECT 212.210 178.275 212.380 178.285 ;
        RECT 212.210 178.115 212.595 178.275 ;
        RECT 211.625 178.065 211.870 178.115 ;
        RECT 212.265 178.105 212.595 178.115 ;
        RECT 212.280 177.895 212.450 177.935 ;
        RECT 212.765 177.930 212.935 178.455 ;
        RECT 213.105 178.005 213.405 179.005 ;
        RECT 213.605 178.635 213.955 179.475 ;
        RECT 214.125 179.305 215.655 179.475 ;
        RECT 214.125 178.805 214.295 179.305 ;
        RECT 215.485 179.145 215.655 179.305 ;
        RECT 215.825 179.265 216.155 179.645 ;
        RECT 214.465 178.965 214.795 179.135 ;
        RECT 214.625 178.635 214.795 178.965 ;
        RECT 214.965 178.975 215.135 179.135 ;
        RECT 216.325 178.975 216.495 179.475 ;
        RECT 214.965 178.805 216.495 178.975 ;
        RECT 213.605 178.405 214.410 178.635 ;
        RECT 214.625 178.465 215.260 178.635 ;
        RECT 214.050 178.295 214.410 178.405 ;
        RECT 214.050 178.115 214.590 178.295 ;
        RECT 210.930 177.725 212.450 177.895 ;
        RECT 208.770 177.435 208.940 177.595 ;
        RECT 207.945 177.265 208.940 177.435 ;
        RECT 209.110 177.425 209.640 177.595 ;
        RECT 209.470 177.265 209.640 177.425 ;
        RECT 209.985 177.335 210.160 177.665 ;
        RECT 210.330 177.095 210.660 177.475 ;
        RECT 210.930 177.305 211.175 177.725 ;
        RECT 212.280 177.605 212.450 177.725 ;
        RECT 212.620 177.855 212.935 177.930 ;
        RECT 212.620 177.605 212.950 177.855 ;
        RECT 211.350 177.095 211.520 177.555 ;
        RECT 211.690 177.435 212.045 177.475 ;
        RECT 213.120 177.435 213.290 177.805 ;
        RECT 211.690 177.265 213.290 177.435 ;
        RECT 213.580 177.095 213.870 177.815 ;
        RECT 214.050 177.440 214.410 178.115 ;
        RECT 215.090 177.945 215.260 178.465 ;
        RECT 215.430 178.005 215.865 178.625 ;
        RECT 216.175 178.285 216.520 178.625 ;
        RECT 216.755 178.480 217.045 179.645 ;
        RECT 217.305 178.715 217.475 179.475 ;
        RECT 217.655 178.885 217.985 179.645 ;
        RECT 217.305 178.545 217.970 178.715 ;
        RECT 218.155 178.570 218.425 179.475 ;
        RECT 217.800 178.400 217.970 178.545 ;
        RECT 216.175 178.115 216.525 178.285 ;
        RECT 216.175 178.005 216.520 178.115 ;
        RECT 217.235 177.995 217.565 178.365 ;
        RECT 217.800 178.070 218.085 178.400 ;
        RECT 214.970 177.775 215.260 177.945 ;
        RECT 214.580 177.435 214.750 177.770 ;
        RECT 214.920 177.605 215.260 177.775 ;
        RECT 215.485 177.645 216.495 177.815 ;
        RECT 215.485 177.435 215.655 177.645 ;
        RECT 214.580 177.265 215.655 177.435 ;
        RECT 215.825 177.095 216.155 177.475 ;
        RECT 216.325 177.270 216.495 177.645 ;
        RECT 216.755 177.095 217.045 177.820 ;
        RECT 217.800 177.815 217.970 178.070 ;
        RECT 217.305 177.645 217.970 177.815 ;
        RECT 218.255 177.770 218.425 178.570 ;
        RECT 218.685 178.715 218.855 179.475 ;
        RECT 219.035 178.885 219.365 179.645 ;
        RECT 218.685 178.545 219.350 178.715 ;
        RECT 219.535 178.570 219.805 179.475 ;
        RECT 220.065 178.975 220.235 179.475 ;
        RECT 220.405 179.265 220.735 179.645 ;
        RECT 220.905 179.305 222.435 179.475 ;
        RECT 220.905 179.145 221.075 179.305 ;
        RECT 221.425 178.975 221.595 179.135 ;
        RECT 220.065 178.805 221.595 178.975 ;
        RECT 221.765 178.965 222.095 179.135 ;
        RECT 221.765 178.635 221.935 178.965 ;
        RECT 222.265 178.805 222.435 179.305 ;
        RECT 222.605 178.635 222.955 179.475 ;
        RECT 223.125 179.265 223.455 179.645 ;
        RECT 223.715 179.305 224.725 179.475 ;
        RECT 219.180 178.400 219.350 178.545 ;
        RECT 218.615 177.995 218.945 178.365 ;
        RECT 219.180 178.070 219.465 178.400 ;
        RECT 219.180 177.815 219.350 178.070 ;
        RECT 217.305 177.265 217.475 177.645 ;
        RECT 217.655 177.095 217.985 177.475 ;
        RECT 218.165 177.265 218.425 177.770 ;
        RECT 218.685 177.645 219.350 177.815 ;
        RECT 219.635 177.770 219.805 178.570 ;
        RECT 220.040 178.285 220.385 178.625 ;
        RECT 220.035 178.115 220.385 178.285 ;
        RECT 220.040 178.005 220.385 178.115 ;
        RECT 220.695 178.005 221.130 178.625 ;
        RECT 221.300 178.465 221.935 178.635 ;
        RECT 221.300 177.945 221.470 178.465 ;
        RECT 222.150 178.405 222.955 178.635 ;
        RECT 222.150 178.295 222.510 178.405 ;
        RECT 221.970 178.115 222.510 178.295 ;
        RECT 218.685 177.265 218.855 177.645 ;
        RECT 219.035 177.095 219.365 177.475 ;
        RECT 219.545 177.265 219.805 177.770 ;
        RECT 220.065 177.645 221.075 177.815 ;
        RECT 220.065 177.270 220.235 177.645 ;
        RECT 220.405 177.095 220.735 177.475 ;
        RECT 220.905 177.435 221.075 177.645 ;
        RECT 221.300 177.775 221.590 177.945 ;
        RECT 221.300 177.605 221.640 177.775 ;
        RECT 221.810 177.435 221.980 177.770 ;
        RECT 222.150 177.440 222.510 178.115 ;
        RECT 223.155 178.005 223.455 179.005 ;
        RECT 223.715 178.795 223.885 179.305 ;
        RECT 224.055 178.625 224.385 179.135 ;
        RECT 224.555 179.095 224.725 179.305 ;
        RECT 224.950 179.265 225.280 179.645 ;
        RECT 225.450 179.095 225.620 179.475 ;
        RECT 225.870 179.265 226.220 179.645 ;
        RECT 226.390 179.145 226.575 179.475 ;
        RECT 224.555 178.925 225.620 179.095 ;
        RECT 223.625 178.455 224.385 178.625 ;
        RECT 223.625 177.930 223.795 178.455 ;
        RECT 224.690 178.285 224.935 178.685 ;
        RECT 224.180 178.275 224.350 178.285 ;
        RECT 223.965 178.115 224.350 178.275 ;
        RECT 224.635 178.115 224.935 178.285 ;
        RECT 223.965 178.105 224.295 178.115 ;
        RECT 224.690 178.065 224.935 178.115 ;
        RECT 225.140 178.625 225.470 178.685 ;
        RECT 225.140 178.455 225.495 178.625 ;
        RECT 225.140 178.065 225.470 178.455 ;
        RECT 225.945 178.005 226.235 178.685 ;
        RECT 226.405 178.285 226.575 179.145 ;
        RECT 226.870 179.145 227.080 179.475 ;
        RECT 227.250 179.305 228.535 179.475 ;
        RECT 227.250 179.265 227.580 179.305 ;
        RECT 226.405 178.115 226.695 178.285 ;
        RECT 223.625 177.855 223.940 177.930 ;
        RECT 220.905 177.265 221.980 177.435 ;
        RECT 222.690 177.095 222.980 177.815 ;
        RECT 223.270 177.435 223.440 177.805 ;
        RECT 223.610 177.605 223.940 177.855 ;
        RECT 224.110 177.895 224.280 177.935 ;
        RECT 224.110 177.725 225.630 177.895 ;
        RECT 224.110 177.605 224.280 177.725 ;
        RECT 224.515 177.435 224.870 177.475 ;
        RECT 223.270 177.265 224.870 177.435 ;
        RECT 225.040 177.095 225.210 177.555 ;
        RECT 225.385 177.305 225.630 177.725 ;
        RECT 226.405 177.665 226.575 178.115 ;
        RECT 226.870 177.945 227.040 179.145 ;
        RECT 227.735 178.995 228.065 179.135 ;
        RECT 227.280 178.765 228.065 178.995 ;
        RECT 228.365 178.845 228.535 179.305 ;
        RECT 228.705 179.265 229.035 179.645 ;
        RECT 226.870 177.775 227.110 177.945 ;
        RECT 225.900 177.095 226.230 177.475 ;
        RECT 226.400 177.335 226.575 177.665 ;
        RECT 227.280 177.595 227.450 178.765 ;
        RECT 228.365 178.675 229.015 178.845 ;
        RECT 228.080 178.115 228.535 178.285 ;
        RECT 227.860 177.935 228.270 177.945 ;
        RECT 227.860 177.775 228.275 177.935 ;
        RECT 228.845 177.895 229.015 178.675 ;
        RECT 228.100 177.605 228.275 177.775 ;
        RECT 228.445 177.725 229.015 177.895 ;
        RECT 226.920 177.425 227.450 177.595 ;
        RECT 227.620 177.435 227.790 177.595 ;
        RECT 228.445 177.435 228.615 177.725 ;
        RECT 226.920 177.265 227.090 177.425 ;
        RECT 227.620 177.265 228.615 177.435 ;
        RECT 228.785 177.095 228.955 177.555 ;
        RECT 229.205 177.265 229.465 179.475 ;
        RECT 229.635 178.480 229.925 179.645 ;
        RECT 230.095 178.570 230.365 179.475 ;
        RECT 230.535 178.885 230.865 179.645 ;
        RECT 231.045 178.715 231.215 179.475 ;
        RECT 229.635 177.095 229.925 177.820 ;
        RECT 230.095 177.770 230.265 178.570 ;
        RECT 230.550 178.545 231.215 178.715 ;
        RECT 231.475 178.570 231.745 179.475 ;
        RECT 231.915 178.885 232.245 179.645 ;
        RECT 232.425 178.715 232.595 179.475 ;
        RECT 230.550 178.400 230.720 178.545 ;
        RECT 230.435 178.070 230.720 178.400 ;
        RECT 230.550 177.815 230.720 178.070 ;
        RECT 230.955 177.995 231.285 178.365 ;
        RECT 230.095 177.265 230.355 177.770 ;
        RECT 230.550 177.645 231.215 177.815 ;
        RECT 230.535 177.095 230.865 177.475 ;
        RECT 231.045 177.265 231.215 177.645 ;
        RECT 231.475 177.770 231.645 178.570 ;
        RECT 231.930 178.545 232.595 178.715 ;
        RECT 232.855 178.570 233.125 179.475 ;
        RECT 233.295 178.885 233.625 179.645 ;
        RECT 233.805 178.715 233.975 179.475 ;
        RECT 231.930 178.400 232.100 178.545 ;
        RECT 231.815 178.070 232.100 178.400 ;
        RECT 231.930 177.815 232.100 178.070 ;
        RECT 232.335 177.995 232.665 178.365 ;
        RECT 231.475 177.265 231.735 177.770 ;
        RECT 231.930 177.645 232.595 177.815 ;
        RECT 231.915 177.095 232.245 177.475 ;
        RECT 232.425 177.265 232.595 177.645 ;
        RECT 232.855 177.770 233.025 178.570 ;
        RECT 233.310 178.545 233.975 178.715 ;
        RECT 234.235 178.570 234.505 179.475 ;
        RECT 234.675 178.885 235.005 179.645 ;
        RECT 235.185 178.715 235.355 179.475 ;
        RECT 233.310 178.400 233.480 178.545 ;
        RECT 233.195 178.070 233.480 178.400 ;
        RECT 233.310 177.815 233.480 178.070 ;
        RECT 233.715 177.995 234.045 178.365 ;
        RECT 232.855 177.265 233.115 177.770 ;
        RECT 233.310 177.645 233.975 177.815 ;
        RECT 233.295 177.095 233.625 177.475 ;
        RECT 233.805 177.265 233.975 177.645 ;
        RECT 234.235 177.770 234.405 178.570 ;
        RECT 234.690 178.545 235.355 178.715 ;
        RECT 235.615 178.570 235.885 179.475 ;
        RECT 236.055 178.885 236.385 179.645 ;
        RECT 236.565 178.715 236.735 179.475 ;
        RECT 234.690 178.400 234.860 178.545 ;
        RECT 234.575 178.070 234.860 178.400 ;
        RECT 234.690 177.815 234.860 178.070 ;
        RECT 235.095 177.995 235.425 178.365 ;
        RECT 234.235 177.265 234.495 177.770 ;
        RECT 234.690 177.645 235.355 177.815 ;
        RECT 234.675 177.095 235.005 177.475 ;
        RECT 235.185 177.265 235.355 177.645 ;
        RECT 235.615 177.770 235.785 178.570 ;
        RECT 236.070 178.545 236.735 178.715 ;
        RECT 237.915 178.555 239.125 179.645 ;
        RECT 236.070 178.400 236.240 178.545 ;
        RECT 235.955 178.070 236.240 178.400 ;
        RECT 236.070 177.815 236.240 178.070 ;
        RECT 236.475 177.995 236.805 178.365 ;
        RECT 237.915 178.015 238.435 178.555 ;
        RECT 238.605 177.845 239.125 178.385 ;
        RECT 235.615 177.265 235.875 177.770 ;
        RECT 236.070 177.645 236.735 177.815 ;
        RECT 236.055 177.095 236.385 177.475 ;
        RECT 236.565 177.265 236.735 177.645 ;
        RECT 237.915 177.095 239.125 177.845 ;
        RECT 165.150 176.925 239.210 177.095 ;
        RECT 162.095 106.340 311.135 106.510 ;
        RECT 162.180 105.590 163.390 106.340 ;
        RECT 162.180 105.050 162.700 105.590 ;
        RECT 164.025 105.500 164.285 106.340 ;
        RECT 164.460 105.595 164.715 106.170 ;
        RECT 164.885 105.960 165.215 106.340 ;
        RECT 165.430 105.790 165.600 106.170 ;
        RECT 164.885 105.620 165.600 105.790 ;
        RECT 162.870 104.880 163.390 105.420 ;
        RECT 162.180 103.790 163.390 104.880 ;
        RECT 164.025 103.790 164.285 104.940 ;
        RECT 164.460 104.865 164.630 105.595 ;
        RECT 164.885 105.430 165.055 105.620 ;
        RECT 164.800 105.100 165.055 105.430 ;
        RECT 164.885 104.890 165.055 105.100 ;
        RECT 165.335 105.070 165.690 105.440 ;
        RECT 164.460 103.960 164.715 104.865 ;
        RECT 164.885 104.720 165.600 104.890 ;
        RECT 164.885 103.790 165.215 104.550 ;
        RECT 165.430 103.960 165.600 104.720 ;
        RECT 166.780 103.960 167.530 106.170 ;
        RECT 167.760 105.860 168.040 106.340 ;
        RECT 168.210 105.690 168.470 106.080 ;
        RECT 168.645 105.860 168.900 106.340 ;
        RECT 169.070 105.690 169.365 106.080 ;
        RECT 169.545 105.860 169.820 106.340 ;
        RECT 169.990 105.840 170.290 106.170 ;
        RECT 167.715 105.520 169.365 105.690 ;
        RECT 167.715 105.010 168.120 105.520 ;
        RECT 168.290 105.180 169.430 105.350 ;
        RECT 167.715 104.840 168.470 105.010 ;
        RECT 167.755 103.790 168.040 104.660 ;
        RECT 168.210 104.590 168.470 104.840 ;
        RECT 169.260 104.930 169.430 105.180 ;
        RECT 169.600 105.100 169.950 105.670 ;
        RECT 170.120 104.930 170.290 105.840 ;
        RECT 170.465 105.500 170.725 106.340 ;
        RECT 170.900 105.595 171.155 106.170 ;
        RECT 171.325 105.960 171.655 106.340 ;
        RECT 171.870 105.790 172.040 106.170 ;
        RECT 172.360 105.860 172.640 106.340 ;
        RECT 171.325 105.620 172.040 105.790 ;
        RECT 172.810 105.690 173.070 106.080 ;
        RECT 173.245 105.860 173.500 106.340 ;
        RECT 173.670 105.690 173.965 106.080 ;
        RECT 174.145 105.860 174.420 106.340 ;
        RECT 174.590 105.840 174.890 106.170 ;
        RECT 169.260 104.760 170.290 104.930 ;
        RECT 168.210 104.420 169.330 104.590 ;
        RECT 168.210 103.960 168.470 104.420 ;
        RECT 168.645 103.790 168.900 104.250 ;
        RECT 169.070 103.960 169.330 104.420 ;
        RECT 169.500 103.790 169.810 104.590 ;
        RECT 169.980 103.960 170.290 104.760 ;
        RECT 170.465 103.790 170.725 104.940 ;
        RECT 170.900 104.865 171.070 105.595 ;
        RECT 171.325 105.430 171.495 105.620 ;
        RECT 172.315 105.520 173.965 105.690 ;
        RECT 171.240 105.100 171.495 105.430 ;
        RECT 171.325 104.890 171.495 105.100 ;
        RECT 171.775 105.070 172.130 105.440 ;
        RECT 172.315 105.010 172.720 105.520 ;
        RECT 172.890 105.180 174.030 105.350 ;
        RECT 170.900 103.960 171.155 104.865 ;
        RECT 171.325 104.720 172.040 104.890 ;
        RECT 172.315 104.840 173.070 105.010 ;
        RECT 171.325 103.790 171.655 104.550 ;
        RECT 171.870 103.960 172.040 104.720 ;
        RECT 172.355 103.790 172.640 104.660 ;
        RECT 172.810 104.590 173.070 104.840 ;
        RECT 173.860 104.930 174.030 105.180 ;
        RECT 174.200 105.100 174.550 105.670 ;
        RECT 174.720 104.930 174.890 105.840 ;
        RECT 175.060 105.615 175.350 106.340 ;
        RECT 176.070 105.790 176.240 106.170 ;
        RECT 176.455 105.960 176.785 106.340 ;
        RECT 176.070 105.620 176.785 105.790 ;
        RECT 175.980 105.070 176.335 105.440 ;
        RECT 176.615 105.430 176.785 105.620 ;
        RECT 176.955 105.595 177.210 106.170 ;
        RECT 176.615 105.100 176.870 105.430 ;
        RECT 173.860 104.760 174.890 104.930 ;
        RECT 172.810 104.420 173.930 104.590 ;
        RECT 172.810 103.960 173.070 104.420 ;
        RECT 173.245 103.790 173.500 104.250 ;
        RECT 173.670 103.960 173.930 104.420 ;
        RECT 174.100 103.790 174.410 104.590 ;
        RECT 174.580 103.960 174.890 104.760 ;
        RECT 175.060 103.790 175.350 104.955 ;
        RECT 176.615 104.890 176.785 105.100 ;
        RECT 176.070 104.720 176.785 104.890 ;
        RECT 177.040 104.865 177.210 105.595 ;
        RECT 177.385 105.500 177.645 106.340 ;
        RECT 177.910 105.790 178.080 106.170 ;
        RECT 178.295 105.960 178.625 106.340 ;
        RECT 177.910 105.620 178.625 105.790 ;
        RECT 177.820 105.070 178.175 105.440 ;
        RECT 178.455 105.430 178.625 105.620 ;
        RECT 178.795 105.595 179.050 106.170 ;
        RECT 178.455 105.100 178.710 105.430 ;
        RECT 176.070 103.960 176.240 104.720 ;
        RECT 176.455 103.790 176.785 104.550 ;
        RECT 176.955 103.960 177.210 104.865 ;
        RECT 177.385 103.790 177.645 104.940 ;
        RECT 178.455 104.890 178.625 105.100 ;
        RECT 177.910 104.720 178.625 104.890 ;
        RECT 178.880 104.865 179.050 105.595 ;
        RECT 179.225 105.500 179.485 106.340 ;
        RECT 179.720 105.860 180.000 106.340 ;
        RECT 180.170 105.690 180.430 106.080 ;
        RECT 180.605 105.860 180.860 106.340 ;
        RECT 181.030 105.690 181.325 106.080 ;
        RECT 181.505 105.860 181.780 106.340 ;
        RECT 181.950 105.840 182.250 106.170 ;
        RECT 179.675 105.520 181.325 105.690 ;
        RECT 179.675 105.010 180.080 105.520 ;
        RECT 180.250 105.180 181.390 105.350 ;
        RECT 177.910 103.960 178.080 104.720 ;
        RECT 178.295 103.790 178.625 104.550 ;
        RECT 178.795 103.960 179.050 104.865 ;
        RECT 179.225 103.790 179.485 104.940 ;
        RECT 179.675 104.840 180.430 105.010 ;
        RECT 179.715 103.790 180.000 104.660 ;
        RECT 180.170 104.590 180.430 104.840 ;
        RECT 181.220 104.930 181.390 105.180 ;
        RECT 181.560 105.100 181.910 105.670 ;
        RECT 182.080 104.930 182.250 105.840 ;
        RECT 182.510 105.790 182.680 106.170 ;
        RECT 182.895 105.960 183.225 106.340 ;
        RECT 182.510 105.620 183.225 105.790 ;
        RECT 182.420 105.070 182.775 105.440 ;
        RECT 183.055 105.430 183.225 105.620 ;
        RECT 183.395 105.595 183.650 106.170 ;
        RECT 183.055 105.100 183.310 105.430 ;
        RECT 181.220 104.760 182.250 104.930 ;
        RECT 183.055 104.890 183.225 105.100 ;
        RECT 180.170 104.420 181.290 104.590 ;
        RECT 180.170 103.960 180.430 104.420 ;
        RECT 180.605 103.790 180.860 104.250 ;
        RECT 181.030 103.960 181.290 104.420 ;
        RECT 181.460 103.790 181.770 104.590 ;
        RECT 181.940 103.960 182.250 104.760 ;
        RECT 182.510 104.720 183.225 104.890 ;
        RECT 183.480 104.865 183.650 105.595 ;
        RECT 183.825 105.500 184.085 106.340 ;
        RECT 184.265 105.500 184.525 106.340 ;
        RECT 184.700 105.595 184.955 106.170 ;
        RECT 185.125 105.960 185.455 106.340 ;
        RECT 185.670 105.790 185.840 106.170 ;
        RECT 185.125 105.620 185.840 105.790 ;
        RECT 186.190 105.790 186.360 106.170 ;
        RECT 186.575 105.960 186.905 106.340 ;
        RECT 186.190 105.620 186.905 105.790 ;
        RECT 182.510 103.960 182.680 104.720 ;
        RECT 182.895 103.790 183.225 104.550 ;
        RECT 183.395 103.960 183.650 104.865 ;
        RECT 183.825 103.790 184.085 104.940 ;
        RECT 184.265 103.790 184.525 104.940 ;
        RECT 184.700 104.865 184.870 105.595 ;
        RECT 185.125 105.430 185.295 105.620 ;
        RECT 185.040 105.100 185.295 105.430 ;
        RECT 185.125 104.890 185.295 105.100 ;
        RECT 185.575 105.070 185.930 105.440 ;
        RECT 186.100 105.070 186.455 105.440 ;
        RECT 186.735 105.430 186.905 105.620 ;
        RECT 187.075 105.595 187.330 106.170 ;
        RECT 186.735 105.100 186.990 105.430 ;
        RECT 186.735 104.890 186.905 105.100 ;
        RECT 184.700 103.960 184.955 104.865 ;
        RECT 185.125 104.720 185.840 104.890 ;
        RECT 185.125 103.790 185.455 104.550 ;
        RECT 185.670 103.960 185.840 104.720 ;
        RECT 186.190 104.720 186.905 104.890 ;
        RECT 187.160 104.865 187.330 105.595 ;
        RECT 187.505 105.500 187.765 106.340 ;
        RECT 187.940 105.615 188.230 106.340 ;
        RECT 188.460 105.860 188.740 106.340 ;
        RECT 188.910 105.690 189.170 106.080 ;
        RECT 189.345 105.860 189.600 106.340 ;
        RECT 189.770 105.690 190.065 106.080 ;
        RECT 190.245 105.860 190.520 106.340 ;
        RECT 190.690 105.840 190.990 106.170 ;
        RECT 188.415 105.520 190.065 105.690 ;
        RECT 188.415 105.010 188.820 105.520 ;
        RECT 188.990 105.180 190.130 105.350 ;
        RECT 186.190 103.960 186.360 104.720 ;
        RECT 186.575 103.790 186.905 104.550 ;
        RECT 187.075 103.960 187.330 104.865 ;
        RECT 187.505 103.790 187.765 104.940 ;
        RECT 187.940 103.790 188.230 104.955 ;
        RECT 188.415 104.840 189.170 105.010 ;
        RECT 188.455 103.790 188.740 104.660 ;
        RECT 188.910 104.590 189.170 104.840 ;
        RECT 189.960 104.930 190.130 105.180 ;
        RECT 190.300 105.100 190.650 105.670 ;
        RECT 190.820 104.930 190.990 105.840 ;
        RECT 191.160 105.590 192.370 106.340 ;
        RECT 192.600 105.860 192.880 106.340 ;
        RECT 193.050 105.690 193.310 106.080 ;
        RECT 193.485 105.860 193.740 106.340 ;
        RECT 193.910 105.690 194.205 106.080 ;
        RECT 194.385 105.860 194.660 106.340 ;
        RECT 194.830 105.840 195.130 106.170 ;
        RECT 191.160 105.050 191.680 105.590 ;
        RECT 192.555 105.520 194.205 105.690 ;
        RECT 189.960 104.760 190.990 104.930 ;
        RECT 191.850 104.880 192.370 105.420 ;
        RECT 188.910 104.420 190.030 104.590 ;
        RECT 188.910 103.960 189.170 104.420 ;
        RECT 189.345 103.790 189.600 104.250 ;
        RECT 189.770 103.960 190.030 104.420 ;
        RECT 190.200 103.790 190.510 104.590 ;
        RECT 190.680 103.960 190.990 104.760 ;
        RECT 191.160 103.790 192.370 104.880 ;
        RECT 192.555 105.010 192.960 105.520 ;
        RECT 193.130 105.180 194.270 105.350 ;
        RECT 192.555 104.840 193.310 105.010 ;
        RECT 192.595 103.790 192.880 104.660 ;
        RECT 193.050 104.590 193.310 104.840 ;
        RECT 194.100 104.930 194.270 105.180 ;
        RECT 194.440 105.100 194.790 105.670 ;
        RECT 194.960 104.930 195.130 105.840 ;
        RECT 195.390 105.790 195.560 106.170 ;
        RECT 195.775 105.960 196.105 106.340 ;
        RECT 195.390 105.620 196.105 105.790 ;
        RECT 195.300 105.070 195.655 105.440 ;
        RECT 195.935 105.430 196.105 105.620 ;
        RECT 196.275 105.595 196.530 106.170 ;
        RECT 195.935 105.100 196.190 105.430 ;
        RECT 194.100 104.760 195.130 104.930 ;
        RECT 195.935 104.890 196.105 105.100 ;
        RECT 193.050 104.420 194.170 104.590 ;
        RECT 193.050 103.960 193.310 104.420 ;
        RECT 193.485 103.790 193.740 104.250 ;
        RECT 193.910 103.960 194.170 104.420 ;
        RECT 194.340 103.790 194.650 104.590 ;
        RECT 194.820 103.960 195.130 104.760 ;
        RECT 195.390 104.720 196.105 104.890 ;
        RECT 196.360 104.865 196.530 105.595 ;
        RECT 196.705 105.500 196.965 106.340 ;
        RECT 197.145 105.500 197.405 106.340 ;
        RECT 197.580 105.595 197.835 106.170 ;
        RECT 198.005 105.960 198.335 106.340 ;
        RECT 198.550 105.790 198.720 106.170 ;
        RECT 198.005 105.620 198.720 105.790 ;
        RECT 199.070 105.790 199.240 106.170 ;
        RECT 199.455 105.960 199.785 106.340 ;
        RECT 199.070 105.620 199.785 105.790 ;
        RECT 195.390 103.960 195.560 104.720 ;
        RECT 195.775 103.790 196.105 104.550 ;
        RECT 196.275 103.960 196.530 104.865 ;
        RECT 196.705 103.790 196.965 104.940 ;
        RECT 197.145 103.790 197.405 104.940 ;
        RECT 197.580 104.865 197.750 105.595 ;
        RECT 198.005 105.430 198.175 105.620 ;
        RECT 197.920 105.100 198.175 105.430 ;
        RECT 198.005 104.890 198.175 105.100 ;
        RECT 198.455 105.070 198.810 105.440 ;
        RECT 198.980 105.070 199.335 105.440 ;
        RECT 199.615 105.430 199.785 105.620 ;
        RECT 199.955 105.595 200.210 106.170 ;
        RECT 199.615 105.100 199.870 105.430 ;
        RECT 199.615 104.890 199.785 105.100 ;
        RECT 197.580 103.960 197.835 104.865 ;
        RECT 198.005 104.720 198.720 104.890 ;
        RECT 198.005 103.790 198.335 104.550 ;
        RECT 198.550 103.960 198.720 104.720 ;
        RECT 199.070 104.720 199.785 104.890 ;
        RECT 200.040 104.865 200.210 105.595 ;
        RECT 200.385 105.500 200.645 106.340 ;
        RECT 200.820 105.615 201.110 106.340 ;
        RECT 201.340 105.860 201.620 106.340 ;
        RECT 201.790 105.690 202.050 106.080 ;
        RECT 202.225 105.860 202.480 106.340 ;
        RECT 202.650 105.690 202.945 106.080 ;
        RECT 203.125 105.860 203.400 106.340 ;
        RECT 203.570 105.840 203.870 106.170 ;
        RECT 201.295 105.520 202.945 105.690 ;
        RECT 201.295 105.010 201.700 105.520 ;
        RECT 201.870 105.180 203.010 105.350 ;
        RECT 199.070 103.960 199.240 104.720 ;
        RECT 199.455 103.790 199.785 104.550 ;
        RECT 199.955 103.960 200.210 104.865 ;
        RECT 200.385 103.790 200.645 104.940 ;
        RECT 200.820 103.790 201.110 104.955 ;
        RECT 201.295 104.840 202.050 105.010 ;
        RECT 201.335 103.790 201.620 104.660 ;
        RECT 201.790 104.590 202.050 104.840 ;
        RECT 202.840 104.930 203.010 105.180 ;
        RECT 203.180 105.100 203.530 105.670 ;
        RECT 203.700 104.930 203.870 105.840 ;
        RECT 202.840 104.760 203.870 104.930 ;
        RECT 201.790 104.420 202.910 104.590 ;
        RECT 201.790 103.960 202.050 104.420 ;
        RECT 202.225 103.790 202.480 104.250 ;
        RECT 202.650 103.960 202.910 104.420 ;
        RECT 203.080 103.790 203.390 104.590 ;
        RECT 203.560 103.960 203.870 104.760 ;
        RECT 204.040 105.840 204.340 106.170 ;
        RECT 204.510 105.860 204.785 106.340 ;
        RECT 204.040 104.930 204.210 105.840 ;
        RECT 204.965 105.690 205.260 106.080 ;
        RECT 205.430 105.860 205.685 106.340 ;
        RECT 205.860 105.690 206.120 106.080 ;
        RECT 206.290 105.860 206.570 106.340 ;
        RECT 204.380 105.100 204.730 105.670 ;
        RECT 204.965 105.520 206.615 105.690 ;
        RECT 204.900 105.180 206.040 105.350 ;
        RECT 204.900 104.930 205.070 105.180 ;
        RECT 206.210 105.010 206.615 105.520 ;
        RECT 204.040 104.760 205.070 104.930 ;
        RECT 205.860 104.840 206.615 105.010 ;
        RECT 206.805 105.600 207.060 106.170 ;
        RECT 207.230 105.940 207.560 106.340 ;
        RECT 207.985 105.805 208.515 106.170 ;
        RECT 207.985 105.770 208.160 105.805 ;
        RECT 207.230 105.600 208.160 105.770 ;
        RECT 206.805 104.930 206.975 105.600 ;
        RECT 207.230 105.430 207.400 105.600 ;
        RECT 207.145 105.100 207.400 105.430 ;
        RECT 207.625 105.100 207.820 105.430 ;
        RECT 204.040 103.960 204.350 104.760 ;
        RECT 205.860 104.590 206.120 104.840 ;
        RECT 204.520 103.790 204.830 104.590 ;
        RECT 205.000 104.420 206.120 104.590 ;
        RECT 205.000 103.960 205.260 104.420 ;
        RECT 205.430 103.790 205.685 104.250 ;
        RECT 205.860 103.960 206.120 104.420 ;
        RECT 206.290 103.790 206.575 104.660 ;
        RECT 206.805 103.960 207.140 104.930 ;
        RECT 207.310 103.790 207.480 104.930 ;
        RECT 207.650 104.130 207.820 105.100 ;
        RECT 207.990 104.470 208.160 105.600 ;
        RECT 208.330 104.810 208.500 105.610 ;
        RECT 208.705 105.320 208.980 106.170 ;
        RECT 208.700 105.150 208.980 105.320 ;
        RECT 208.705 105.010 208.980 105.150 ;
        RECT 209.150 104.810 209.340 106.170 ;
        RECT 209.520 105.805 210.030 106.340 ;
        RECT 210.250 105.530 210.495 106.135 ;
        RECT 209.540 105.360 210.770 105.530 ;
        RECT 211.865 105.500 212.125 106.340 ;
        RECT 212.300 105.595 212.555 106.170 ;
        RECT 212.725 105.960 213.055 106.340 ;
        RECT 213.270 105.790 213.440 106.170 ;
        RECT 212.725 105.620 213.440 105.790 ;
        RECT 208.330 104.640 209.340 104.810 ;
        RECT 209.510 104.795 210.260 104.985 ;
        RECT 207.990 104.300 209.115 104.470 ;
        RECT 209.510 104.130 209.680 104.795 ;
        RECT 210.430 104.550 210.770 105.360 ;
        RECT 207.650 103.960 209.680 104.130 ;
        RECT 209.850 103.790 210.020 104.550 ;
        RECT 210.255 104.140 210.770 104.550 ;
        RECT 211.865 103.790 212.125 104.940 ;
        RECT 212.300 104.865 212.470 105.595 ;
        RECT 212.725 105.430 212.895 105.620 ;
        RECT 213.700 105.615 213.990 106.340 ;
        RECT 214.220 105.860 214.500 106.340 ;
        RECT 214.670 105.690 214.930 106.080 ;
        RECT 215.105 105.860 215.360 106.340 ;
        RECT 215.530 105.690 215.825 106.080 ;
        RECT 216.005 105.860 216.280 106.340 ;
        RECT 216.450 105.840 216.750 106.170 ;
        RECT 214.175 105.520 215.825 105.690 ;
        RECT 212.640 105.100 212.895 105.430 ;
        RECT 212.725 104.890 212.895 105.100 ;
        RECT 213.175 105.070 213.530 105.440 ;
        RECT 214.175 105.010 214.580 105.520 ;
        RECT 214.750 105.180 215.890 105.350 ;
        RECT 212.300 103.960 212.555 104.865 ;
        RECT 212.725 104.720 213.440 104.890 ;
        RECT 212.725 103.790 213.055 104.550 ;
        RECT 213.270 103.960 213.440 104.720 ;
        RECT 213.700 103.790 213.990 104.955 ;
        RECT 214.175 104.840 214.930 105.010 ;
        RECT 214.215 103.790 214.500 104.660 ;
        RECT 214.670 104.590 214.930 104.840 ;
        RECT 215.720 104.930 215.890 105.180 ;
        RECT 216.060 105.100 216.410 105.670 ;
        RECT 216.580 104.930 216.750 105.840 ;
        RECT 216.920 105.590 218.130 106.340 ;
        RECT 218.390 105.790 218.560 106.170 ;
        RECT 218.775 105.960 219.105 106.340 ;
        RECT 218.390 105.620 219.105 105.790 ;
        RECT 216.920 105.050 217.440 105.590 ;
        RECT 215.720 104.760 216.750 104.930 ;
        RECT 217.610 104.880 218.130 105.420 ;
        RECT 218.300 105.070 218.655 105.440 ;
        RECT 218.935 105.430 219.105 105.620 ;
        RECT 219.275 105.595 219.530 106.170 ;
        RECT 218.935 105.100 219.190 105.430 ;
        RECT 218.935 104.890 219.105 105.100 ;
        RECT 214.670 104.420 215.790 104.590 ;
        RECT 214.670 103.960 214.930 104.420 ;
        RECT 215.105 103.790 215.360 104.250 ;
        RECT 215.530 103.960 215.790 104.420 ;
        RECT 215.960 103.790 216.270 104.590 ;
        RECT 216.440 103.960 216.750 104.760 ;
        RECT 216.920 103.790 218.130 104.880 ;
        RECT 218.390 104.720 219.105 104.890 ;
        RECT 219.360 104.865 219.530 105.595 ;
        RECT 219.705 105.500 219.965 106.340 ;
        RECT 220.140 105.840 220.440 106.170 ;
        RECT 220.610 105.860 220.885 106.340 ;
        RECT 218.390 103.960 218.560 104.720 ;
        RECT 218.775 103.790 219.105 104.550 ;
        RECT 219.275 103.960 219.530 104.865 ;
        RECT 219.705 103.790 219.965 104.940 ;
        RECT 220.140 104.930 220.310 105.840 ;
        RECT 221.065 105.690 221.360 106.080 ;
        RECT 221.530 105.860 221.785 106.340 ;
        RECT 221.960 105.690 222.220 106.080 ;
        RECT 222.390 105.860 222.670 106.340 ;
        RECT 222.990 105.790 223.160 106.170 ;
        RECT 223.375 105.960 223.705 106.340 ;
        RECT 220.480 105.100 220.830 105.670 ;
        RECT 221.065 105.520 222.715 105.690 ;
        RECT 222.990 105.620 223.705 105.790 ;
        RECT 221.000 105.180 222.140 105.350 ;
        RECT 221.000 104.930 221.170 105.180 ;
        RECT 222.310 105.010 222.715 105.520 ;
        RECT 222.900 105.070 223.255 105.440 ;
        RECT 223.535 105.430 223.705 105.620 ;
        RECT 223.875 105.595 224.130 106.170 ;
        RECT 223.535 105.100 223.790 105.430 ;
        RECT 220.140 104.760 221.170 104.930 ;
        RECT 221.960 104.840 222.715 105.010 ;
        RECT 223.535 104.890 223.705 105.100 ;
        RECT 220.140 103.960 220.450 104.760 ;
        RECT 221.960 104.590 222.220 104.840 ;
        RECT 222.990 104.720 223.705 104.890 ;
        RECT 223.960 104.865 224.130 105.595 ;
        RECT 224.305 105.500 224.565 106.340 ;
        RECT 224.830 105.790 225.000 106.170 ;
        RECT 225.215 105.960 225.545 106.340 ;
        RECT 224.830 105.620 225.545 105.790 ;
        RECT 224.740 105.070 225.095 105.440 ;
        RECT 225.375 105.430 225.545 105.620 ;
        RECT 225.715 105.595 225.970 106.170 ;
        RECT 225.375 105.100 225.630 105.430 ;
        RECT 220.620 103.790 220.930 104.590 ;
        RECT 221.100 104.420 222.220 104.590 ;
        RECT 221.100 103.960 221.360 104.420 ;
        RECT 221.530 103.790 221.785 104.250 ;
        RECT 221.960 103.960 222.220 104.420 ;
        RECT 222.390 103.790 222.675 104.660 ;
        RECT 222.990 103.960 223.160 104.720 ;
        RECT 223.375 103.790 223.705 104.550 ;
        RECT 223.875 103.960 224.130 104.865 ;
        RECT 224.305 103.790 224.565 104.940 ;
        RECT 225.375 104.890 225.545 105.100 ;
        RECT 224.830 104.720 225.545 104.890 ;
        RECT 225.800 104.865 225.970 105.595 ;
        RECT 226.145 105.500 226.405 106.340 ;
        RECT 226.580 105.615 226.870 106.340 ;
        RECT 227.560 105.860 227.840 106.340 ;
        RECT 228.010 105.690 228.270 106.080 ;
        RECT 228.445 105.860 228.700 106.340 ;
        RECT 228.870 105.690 229.165 106.080 ;
        RECT 229.345 105.860 229.620 106.340 ;
        RECT 229.790 105.840 230.090 106.170 ;
        RECT 227.515 105.520 229.165 105.690 ;
        RECT 227.515 105.010 227.920 105.520 ;
        RECT 228.090 105.180 229.230 105.350 ;
        RECT 224.830 103.960 225.000 104.720 ;
        RECT 225.215 103.790 225.545 104.550 ;
        RECT 225.715 103.960 225.970 104.865 ;
        RECT 226.145 103.790 226.405 104.940 ;
        RECT 226.580 103.790 226.870 104.955 ;
        RECT 227.515 104.840 228.270 105.010 ;
        RECT 227.555 103.790 227.840 104.660 ;
        RECT 228.010 104.590 228.270 104.840 ;
        RECT 229.060 104.930 229.230 105.180 ;
        RECT 229.400 105.100 229.750 105.670 ;
        RECT 229.920 104.930 230.090 105.840 ;
        RECT 230.350 105.790 230.520 106.170 ;
        RECT 230.735 105.960 231.065 106.340 ;
        RECT 230.350 105.620 231.065 105.790 ;
        RECT 230.260 105.070 230.615 105.440 ;
        RECT 230.895 105.430 231.065 105.620 ;
        RECT 231.235 105.595 231.490 106.170 ;
        RECT 230.895 105.100 231.150 105.430 ;
        RECT 229.060 104.760 230.090 104.930 ;
        RECT 230.895 104.890 231.065 105.100 ;
        RECT 228.010 104.420 229.130 104.590 ;
        RECT 228.010 103.960 228.270 104.420 ;
        RECT 228.445 103.790 228.700 104.250 ;
        RECT 228.870 103.960 229.130 104.420 ;
        RECT 229.300 103.790 229.610 104.590 ;
        RECT 229.780 103.960 230.090 104.760 ;
        RECT 230.350 104.720 231.065 104.890 ;
        RECT 231.320 104.865 231.490 105.595 ;
        RECT 231.665 105.500 231.925 106.340 ;
        RECT 232.190 105.790 232.360 106.170 ;
        RECT 232.575 105.960 232.905 106.340 ;
        RECT 232.190 105.620 232.905 105.790 ;
        RECT 232.100 105.070 232.455 105.440 ;
        RECT 232.735 105.430 232.905 105.620 ;
        RECT 233.075 105.595 233.330 106.170 ;
        RECT 232.735 105.100 232.990 105.430 ;
        RECT 230.350 103.960 230.520 104.720 ;
        RECT 230.735 103.790 231.065 104.550 ;
        RECT 231.235 103.960 231.490 104.865 ;
        RECT 231.665 103.790 231.925 104.940 ;
        RECT 232.735 104.890 232.905 105.100 ;
        RECT 232.190 104.720 232.905 104.890 ;
        RECT 233.160 104.865 233.330 105.595 ;
        RECT 233.505 105.500 233.765 106.340 ;
        RECT 233.940 105.840 234.240 106.170 ;
        RECT 234.410 105.860 234.685 106.340 ;
        RECT 232.190 103.960 232.360 104.720 ;
        RECT 232.575 103.790 232.905 104.550 ;
        RECT 233.075 103.960 233.330 104.865 ;
        RECT 233.505 103.790 233.765 104.940 ;
        RECT 233.940 104.930 234.110 105.840 ;
        RECT 234.865 105.690 235.160 106.080 ;
        RECT 235.330 105.860 235.585 106.340 ;
        RECT 235.760 105.690 236.020 106.080 ;
        RECT 236.190 105.860 236.470 106.340 ;
        RECT 237.710 105.790 237.880 106.170 ;
        RECT 238.095 105.960 238.425 106.340 ;
        RECT 234.280 105.100 234.630 105.670 ;
        RECT 234.865 105.520 236.515 105.690 ;
        RECT 237.710 105.620 238.425 105.790 ;
        RECT 234.800 105.180 235.940 105.350 ;
        RECT 234.800 104.930 234.970 105.180 ;
        RECT 236.110 105.010 236.515 105.520 ;
        RECT 237.620 105.070 237.975 105.440 ;
        RECT 238.255 105.430 238.425 105.620 ;
        RECT 238.595 105.595 238.850 106.170 ;
        RECT 238.255 105.100 238.510 105.430 ;
        RECT 233.940 104.760 234.970 104.930 ;
        RECT 235.760 104.840 236.515 105.010 ;
        RECT 238.255 104.890 238.425 105.100 ;
        RECT 233.940 103.960 234.250 104.760 ;
        RECT 235.760 104.590 236.020 104.840 ;
        RECT 237.710 104.720 238.425 104.890 ;
        RECT 238.680 104.865 238.850 105.595 ;
        RECT 239.025 105.500 239.285 106.340 ;
        RECT 239.460 105.615 239.750 106.340 ;
        RECT 239.925 105.600 240.180 106.170 ;
        RECT 240.350 105.940 240.680 106.340 ;
        RECT 241.105 105.805 241.635 106.170 ;
        RECT 241.105 105.770 241.280 105.805 ;
        RECT 240.350 105.600 241.280 105.770 ;
        RECT 234.420 103.790 234.730 104.590 ;
        RECT 234.900 104.420 236.020 104.590 ;
        RECT 234.900 103.960 235.160 104.420 ;
        RECT 235.330 103.790 235.585 104.250 ;
        RECT 235.760 103.960 236.020 104.420 ;
        RECT 236.190 103.790 236.475 104.660 ;
        RECT 237.710 103.960 237.880 104.720 ;
        RECT 238.095 103.790 238.425 104.550 ;
        RECT 238.595 103.960 238.850 104.865 ;
        RECT 239.025 103.790 239.285 104.940 ;
        RECT 239.460 103.790 239.750 104.955 ;
        RECT 239.925 104.930 240.095 105.600 ;
        RECT 240.350 105.430 240.520 105.600 ;
        RECT 240.265 105.100 240.520 105.430 ;
        RECT 240.745 105.100 240.940 105.430 ;
        RECT 239.925 103.960 240.260 104.930 ;
        RECT 240.430 103.790 240.600 104.930 ;
        RECT 240.770 104.130 240.940 105.100 ;
        RECT 241.110 104.470 241.280 105.600 ;
        RECT 241.450 104.810 241.620 105.610 ;
        RECT 241.825 105.320 242.100 106.170 ;
        RECT 241.820 105.150 242.100 105.320 ;
        RECT 241.825 105.010 242.100 105.150 ;
        RECT 242.270 104.810 242.460 106.170 ;
        RECT 242.640 105.805 243.150 106.340 ;
        RECT 243.370 105.530 243.615 106.135 ;
        RECT 244.335 105.530 244.580 106.135 ;
        RECT 244.800 105.805 245.310 106.340 ;
        RECT 242.660 105.360 243.890 105.530 ;
        RECT 241.450 104.640 242.460 104.810 ;
        RECT 242.630 104.795 243.380 104.985 ;
        RECT 241.110 104.300 242.235 104.470 ;
        RECT 242.630 104.130 242.800 104.795 ;
        RECT 243.550 104.550 243.890 105.360 ;
        RECT 240.770 103.960 242.800 104.130 ;
        RECT 242.970 103.790 243.140 104.550 ;
        RECT 243.375 104.140 243.890 104.550 ;
        RECT 244.060 105.360 245.290 105.530 ;
        RECT 244.060 104.550 244.400 105.360 ;
        RECT 244.570 104.795 245.320 104.985 ;
        RECT 244.060 104.140 244.575 104.550 ;
        RECT 244.810 103.790 244.980 104.550 ;
        RECT 245.150 104.130 245.320 104.795 ;
        RECT 245.490 104.810 245.680 106.170 ;
        RECT 245.850 105.320 246.125 106.170 ;
        RECT 246.315 105.805 246.845 106.170 ;
        RECT 247.270 105.940 247.600 106.340 ;
        RECT 246.670 105.770 246.845 105.805 ;
        RECT 245.850 105.150 246.130 105.320 ;
        RECT 245.850 105.010 246.125 105.150 ;
        RECT 246.330 104.810 246.500 105.610 ;
        RECT 245.490 104.640 246.500 104.810 ;
        RECT 246.670 105.600 247.600 105.770 ;
        RECT 247.770 105.600 248.025 106.170 ;
        RECT 248.260 105.860 248.540 106.340 ;
        RECT 248.710 105.690 248.970 106.080 ;
        RECT 249.145 105.860 249.400 106.340 ;
        RECT 249.570 105.690 249.865 106.080 ;
        RECT 250.045 105.860 250.320 106.340 ;
        RECT 250.490 105.840 250.790 106.170 ;
        RECT 246.670 104.470 246.840 105.600 ;
        RECT 247.430 105.430 247.600 105.600 ;
        RECT 245.715 104.300 246.840 104.470 ;
        RECT 247.010 105.100 247.205 105.430 ;
        RECT 247.430 105.100 247.685 105.430 ;
        RECT 247.010 104.130 247.180 105.100 ;
        RECT 247.855 104.930 248.025 105.600 ;
        RECT 245.150 103.960 247.180 104.130 ;
        RECT 247.350 103.790 247.520 104.930 ;
        RECT 247.690 103.960 248.025 104.930 ;
        RECT 248.215 105.520 249.865 105.690 ;
        RECT 248.215 105.010 248.620 105.520 ;
        RECT 248.790 105.180 249.930 105.350 ;
        RECT 248.215 104.840 248.970 105.010 ;
        RECT 248.255 103.790 248.540 104.660 ;
        RECT 248.710 104.590 248.970 104.840 ;
        RECT 249.760 104.930 249.930 105.180 ;
        RECT 250.100 105.100 250.450 105.670 ;
        RECT 250.620 104.930 250.790 105.840 ;
        RECT 250.960 105.590 252.170 106.340 ;
        RECT 252.340 105.615 252.630 106.340 ;
        RECT 252.860 105.860 253.140 106.340 ;
        RECT 253.310 105.690 253.570 106.080 ;
        RECT 253.745 105.860 254.000 106.340 ;
        RECT 254.170 105.690 254.465 106.080 ;
        RECT 254.645 105.860 254.920 106.340 ;
        RECT 255.090 105.840 255.390 106.170 ;
        RECT 255.620 105.860 255.900 106.340 ;
        RECT 250.960 105.050 251.480 105.590 ;
        RECT 252.815 105.520 254.465 105.690 ;
        RECT 249.760 104.760 250.790 104.930 ;
        RECT 251.650 104.880 252.170 105.420 ;
        RECT 252.815 105.010 253.220 105.520 ;
        RECT 253.390 105.180 254.530 105.350 ;
        RECT 248.710 104.420 249.830 104.590 ;
        RECT 248.710 103.960 248.970 104.420 ;
        RECT 249.145 103.790 249.400 104.250 ;
        RECT 249.570 103.960 249.830 104.420 ;
        RECT 250.000 103.790 250.310 104.590 ;
        RECT 250.480 103.960 250.790 104.760 ;
        RECT 250.960 103.790 252.170 104.880 ;
        RECT 252.340 103.790 252.630 104.955 ;
        RECT 252.815 104.840 253.570 105.010 ;
        RECT 252.855 103.790 253.140 104.660 ;
        RECT 253.310 104.590 253.570 104.840 ;
        RECT 254.360 104.930 254.530 105.180 ;
        RECT 254.700 105.100 255.050 105.670 ;
        RECT 255.220 104.930 255.390 105.840 ;
        RECT 256.070 105.690 256.330 106.080 ;
        RECT 256.505 105.860 256.760 106.340 ;
        RECT 256.930 105.690 257.225 106.080 ;
        RECT 257.405 105.860 257.680 106.340 ;
        RECT 257.850 105.840 258.150 106.170 ;
        RECT 254.360 104.760 255.390 104.930 ;
        RECT 255.575 105.520 257.225 105.690 ;
        RECT 255.575 105.010 255.980 105.520 ;
        RECT 256.150 105.180 257.290 105.350 ;
        RECT 255.575 104.840 256.330 105.010 ;
        RECT 253.310 104.420 254.430 104.590 ;
        RECT 253.310 103.960 253.570 104.420 ;
        RECT 253.745 103.790 254.000 104.250 ;
        RECT 254.170 103.960 254.430 104.420 ;
        RECT 254.600 103.790 254.910 104.590 ;
        RECT 255.080 103.960 255.390 104.760 ;
        RECT 255.615 103.790 255.900 104.660 ;
        RECT 256.070 104.590 256.330 104.840 ;
        RECT 257.120 104.930 257.290 105.180 ;
        RECT 257.460 105.100 257.810 105.670 ;
        RECT 257.980 104.930 258.150 105.840 ;
        RECT 258.325 105.500 258.585 106.340 ;
        RECT 258.760 105.595 259.015 106.170 ;
        RECT 259.185 105.960 259.515 106.340 ;
        RECT 259.730 105.790 259.900 106.170 ;
        RECT 261.140 105.860 261.420 106.340 ;
        RECT 259.185 105.620 259.900 105.790 ;
        RECT 261.590 105.690 261.850 106.080 ;
        RECT 262.025 105.860 262.280 106.340 ;
        RECT 262.450 105.690 262.745 106.080 ;
        RECT 262.925 105.860 263.200 106.340 ;
        RECT 263.370 105.840 263.670 106.170 ;
        RECT 257.120 104.760 258.150 104.930 ;
        RECT 256.070 104.420 257.190 104.590 ;
        RECT 256.070 103.960 256.330 104.420 ;
        RECT 256.505 103.790 256.760 104.250 ;
        RECT 256.930 103.960 257.190 104.420 ;
        RECT 257.360 103.790 257.670 104.590 ;
        RECT 257.840 103.960 258.150 104.760 ;
        RECT 258.325 103.790 258.585 104.940 ;
        RECT 258.760 104.865 258.930 105.595 ;
        RECT 259.185 105.430 259.355 105.620 ;
        RECT 261.095 105.520 262.745 105.690 ;
        RECT 259.100 105.100 259.355 105.430 ;
        RECT 259.185 104.890 259.355 105.100 ;
        RECT 259.635 105.070 259.990 105.440 ;
        RECT 261.095 105.010 261.500 105.520 ;
        RECT 261.670 105.180 262.810 105.350 ;
        RECT 258.760 103.960 259.015 104.865 ;
        RECT 259.185 104.720 259.900 104.890 ;
        RECT 261.095 104.840 261.850 105.010 ;
        RECT 259.185 103.790 259.515 104.550 ;
        RECT 259.730 103.960 259.900 104.720 ;
        RECT 261.135 103.790 261.420 104.660 ;
        RECT 261.590 104.590 261.850 104.840 ;
        RECT 262.640 104.930 262.810 105.180 ;
        RECT 262.980 105.100 263.330 105.670 ;
        RECT 263.500 104.930 263.670 105.840 ;
        RECT 263.840 105.590 265.050 106.340 ;
        RECT 265.220 105.615 265.510 106.340 ;
        RECT 263.840 105.050 264.360 105.590 ;
        RECT 265.685 105.500 265.945 106.340 ;
        RECT 266.120 105.595 266.375 106.170 ;
        RECT 266.545 105.960 266.875 106.340 ;
        RECT 267.090 105.790 267.260 106.170 ;
        RECT 268.500 105.860 268.780 106.340 ;
        RECT 266.545 105.620 267.260 105.790 ;
        RECT 268.950 105.690 269.210 106.080 ;
        RECT 269.385 105.860 269.640 106.340 ;
        RECT 269.810 105.690 270.105 106.080 ;
        RECT 270.285 105.860 270.560 106.340 ;
        RECT 270.730 105.840 271.030 106.170 ;
        RECT 271.260 105.860 271.540 106.340 ;
        RECT 262.640 104.760 263.670 104.930 ;
        RECT 264.530 104.880 265.050 105.420 ;
        RECT 261.590 104.420 262.710 104.590 ;
        RECT 261.590 103.960 261.850 104.420 ;
        RECT 262.025 103.790 262.280 104.250 ;
        RECT 262.450 103.960 262.710 104.420 ;
        RECT 262.880 103.790 263.190 104.590 ;
        RECT 263.360 103.960 263.670 104.760 ;
        RECT 263.840 103.790 265.050 104.880 ;
        RECT 265.220 103.790 265.510 104.955 ;
        RECT 265.685 103.790 265.945 104.940 ;
        RECT 266.120 104.865 266.290 105.595 ;
        RECT 266.545 105.430 266.715 105.620 ;
        RECT 268.455 105.520 270.105 105.690 ;
        RECT 266.460 105.100 266.715 105.430 ;
        RECT 266.545 104.890 266.715 105.100 ;
        RECT 266.995 105.070 267.350 105.440 ;
        RECT 268.455 105.010 268.860 105.520 ;
        RECT 269.030 105.180 270.170 105.350 ;
        RECT 266.120 103.960 266.375 104.865 ;
        RECT 266.545 104.720 267.260 104.890 ;
        RECT 268.455 104.840 269.210 105.010 ;
        RECT 266.545 103.790 266.875 104.550 ;
        RECT 267.090 103.960 267.260 104.720 ;
        RECT 268.495 103.790 268.780 104.660 ;
        RECT 268.950 104.590 269.210 104.840 ;
        RECT 270.000 104.930 270.170 105.180 ;
        RECT 270.340 105.100 270.690 105.670 ;
        RECT 270.860 104.930 271.030 105.840 ;
        RECT 271.710 105.690 271.970 106.080 ;
        RECT 272.145 105.860 272.400 106.340 ;
        RECT 272.570 105.690 272.865 106.080 ;
        RECT 273.045 105.860 273.320 106.340 ;
        RECT 273.490 105.840 273.790 106.170 ;
        RECT 270.000 104.760 271.030 104.930 ;
        RECT 271.215 105.520 272.865 105.690 ;
        RECT 271.215 105.010 271.620 105.520 ;
        RECT 271.790 105.180 272.930 105.350 ;
        RECT 271.215 104.840 271.970 105.010 ;
        RECT 268.950 104.420 270.070 104.590 ;
        RECT 268.950 103.960 269.210 104.420 ;
        RECT 269.385 103.790 269.640 104.250 ;
        RECT 269.810 103.960 270.070 104.420 ;
        RECT 270.240 103.790 270.550 104.590 ;
        RECT 270.720 103.960 271.030 104.760 ;
        RECT 271.255 103.790 271.540 104.660 ;
        RECT 271.710 104.590 271.970 104.840 ;
        RECT 272.760 104.930 272.930 105.180 ;
        RECT 273.100 105.100 273.450 105.670 ;
        RECT 273.620 104.930 273.790 105.840 ;
        RECT 273.965 105.500 274.225 106.340 ;
        RECT 274.400 105.595 274.655 106.170 ;
        RECT 274.825 105.960 275.155 106.340 ;
        RECT 275.370 105.790 275.540 106.170 ;
        RECT 274.825 105.620 275.540 105.790 ;
        RECT 272.760 104.760 273.790 104.930 ;
        RECT 271.710 104.420 272.830 104.590 ;
        RECT 271.710 103.960 271.970 104.420 ;
        RECT 272.145 103.790 272.400 104.250 ;
        RECT 272.570 103.960 272.830 104.420 ;
        RECT 273.000 103.790 273.310 104.590 ;
        RECT 273.480 103.960 273.790 104.760 ;
        RECT 273.965 103.790 274.225 104.940 ;
        RECT 274.400 104.865 274.570 105.595 ;
        RECT 274.825 105.430 274.995 105.620 ;
        RECT 275.805 105.500 276.065 106.340 ;
        RECT 276.240 105.595 276.495 106.170 ;
        RECT 276.665 105.960 276.995 106.340 ;
        RECT 277.210 105.790 277.380 106.170 ;
        RECT 276.665 105.620 277.380 105.790 ;
        RECT 274.740 105.100 274.995 105.430 ;
        RECT 274.825 104.890 274.995 105.100 ;
        RECT 275.275 105.070 275.630 105.440 ;
        RECT 274.400 103.960 274.655 104.865 ;
        RECT 274.825 104.720 275.540 104.890 ;
        RECT 274.825 103.790 275.155 104.550 ;
        RECT 275.370 103.960 275.540 104.720 ;
        RECT 275.805 103.790 276.065 104.940 ;
        RECT 276.240 104.865 276.410 105.595 ;
        RECT 276.665 105.430 276.835 105.620 ;
        RECT 278.100 105.615 278.390 106.340 ;
        RECT 278.620 105.860 278.900 106.340 ;
        RECT 279.070 105.690 279.330 106.080 ;
        RECT 279.505 105.860 279.760 106.340 ;
        RECT 279.930 105.690 280.225 106.080 ;
        RECT 280.405 105.860 280.680 106.340 ;
        RECT 280.850 105.840 281.150 106.170 ;
        RECT 278.575 105.520 280.225 105.690 ;
        RECT 276.580 105.100 276.835 105.430 ;
        RECT 276.665 104.890 276.835 105.100 ;
        RECT 277.115 105.070 277.470 105.440 ;
        RECT 278.575 105.010 278.980 105.520 ;
        RECT 279.150 105.180 280.290 105.350 ;
        RECT 276.240 103.960 276.495 104.865 ;
        RECT 276.665 104.720 277.380 104.890 ;
        RECT 276.665 103.790 276.995 104.550 ;
        RECT 277.210 103.960 277.380 104.720 ;
        RECT 278.100 103.790 278.390 104.955 ;
        RECT 278.575 104.840 279.330 105.010 ;
        RECT 278.615 103.790 278.900 104.660 ;
        RECT 279.070 104.590 279.330 104.840 ;
        RECT 280.120 104.930 280.290 105.180 ;
        RECT 280.460 105.100 280.810 105.670 ;
        RECT 280.980 104.930 281.150 105.840 ;
        RECT 281.325 105.500 281.585 106.340 ;
        RECT 281.760 105.595 282.015 106.170 ;
        RECT 282.185 105.960 282.515 106.340 ;
        RECT 282.730 105.790 282.900 106.170 ;
        RECT 283.220 105.860 283.500 106.340 ;
        RECT 282.185 105.620 282.900 105.790 ;
        RECT 283.670 105.690 283.930 106.080 ;
        RECT 284.105 105.860 284.360 106.340 ;
        RECT 284.530 105.690 284.825 106.080 ;
        RECT 285.005 105.860 285.280 106.340 ;
        RECT 285.450 105.840 285.750 106.170 ;
        RECT 280.120 104.760 281.150 104.930 ;
        RECT 279.070 104.420 280.190 104.590 ;
        RECT 279.070 103.960 279.330 104.420 ;
        RECT 279.505 103.790 279.760 104.250 ;
        RECT 279.930 103.960 280.190 104.420 ;
        RECT 280.360 103.790 280.670 104.590 ;
        RECT 280.840 103.960 281.150 104.760 ;
        RECT 281.325 103.790 281.585 104.940 ;
        RECT 281.760 104.865 281.930 105.595 ;
        RECT 282.185 105.430 282.355 105.620 ;
        RECT 283.175 105.520 284.825 105.690 ;
        RECT 282.100 105.100 282.355 105.430 ;
        RECT 282.185 104.890 282.355 105.100 ;
        RECT 282.635 105.070 282.990 105.440 ;
        RECT 283.175 105.010 283.580 105.520 ;
        RECT 283.750 105.180 284.890 105.350 ;
        RECT 281.760 103.960 282.015 104.865 ;
        RECT 282.185 104.720 282.900 104.890 ;
        RECT 283.175 104.840 283.930 105.010 ;
        RECT 282.185 103.790 282.515 104.550 ;
        RECT 282.730 103.960 282.900 104.720 ;
        RECT 283.215 103.790 283.500 104.660 ;
        RECT 283.670 104.590 283.930 104.840 ;
        RECT 284.720 104.930 284.890 105.180 ;
        RECT 285.060 105.100 285.410 105.670 ;
        RECT 285.580 104.930 285.750 105.840 ;
        RECT 285.925 105.500 286.185 106.340 ;
        RECT 286.360 105.595 286.615 106.170 ;
        RECT 286.785 105.960 287.115 106.340 ;
        RECT 287.330 105.790 287.500 106.170 ;
        RECT 286.785 105.620 287.500 105.790 ;
        RECT 284.720 104.760 285.750 104.930 ;
        RECT 283.670 104.420 284.790 104.590 ;
        RECT 283.670 103.960 283.930 104.420 ;
        RECT 284.105 103.790 284.360 104.250 ;
        RECT 284.530 103.960 284.790 104.420 ;
        RECT 284.960 103.790 285.270 104.590 ;
        RECT 285.440 103.960 285.750 104.760 ;
        RECT 285.925 103.790 286.185 104.940 ;
        RECT 286.360 104.865 286.530 105.595 ;
        RECT 286.785 105.430 286.955 105.620 ;
        RECT 287.765 105.500 288.025 106.340 ;
        RECT 288.200 105.595 288.455 106.170 ;
        RECT 288.625 105.960 288.955 106.340 ;
        RECT 289.170 105.790 289.340 106.170 ;
        RECT 288.625 105.620 289.340 105.790 ;
        RECT 289.600 105.665 289.860 106.170 ;
        RECT 290.040 105.960 290.370 106.340 ;
        RECT 290.550 105.790 290.720 106.170 ;
        RECT 286.700 105.100 286.955 105.430 ;
        RECT 286.785 104.890 286.955 105.100 ;
        RECT 287.235 105.070 287.590 105.440 ;
        RECT 286.360 103.960 286.615 104.865 ;
        RECT 286.785 104.720 287.500 104.890 ;
        RECT 286.785 103.790 287.115 104.550 ;
        RECT 287.330 103.960 287.500 104.720 ;
        RECT 287.765 103.790 288.025 104.940 ;
        RECT 288.200 104.865 288.370 105.595 ;
        RECT 288.625 105.430 288.795 105.620 ;
        RECT 288.540 105.100 288.795 105.430 ;
        RECT 288.625 104.890 288.795 105.100 ;
        RECT 289.075 105.070 289.430 105.440 ;
        RECT 288.200 103.960 288.455 104.865 ;
        RECT 288.625 104.720 289.340 104.890 ;
        RECT 288.625 103.790 288.955 104.550 ;
        RECT 289.170 103.960 289.340 104.720 ;
        RECT 289.600 104.865 289.770 105.665 ;
        RECT 290.055 105.620 290.720 105.790 ;
        RECT 290.055 105.365 290.225 105.620 ;
        RECT 290.980 105.615 291.270 106.340 ;
        RECT 291.500 105.860 291.780 106.340 ;
        RECT 291.950 105.690 292.210 106.080 ;
        RECT 292.385 105.860 292.640 106.340 ;
        RECT 292.810 105.690 293.105 106.080 ;
        RECT 293.285 105.860 293.560 106.340 ;
        RECT 293.730 105.840 294.030 106.170 ;
        RECT 291.455 105.520 293.105 105.690 ;
        RECT 289.940 105.035 290.225 105.365 ;
        RECT 290.460 105.070 290.790 105.440 ;
        RECT 290.055 104.890 290.225 105.035 ;
        RECT 291.455 105.010 291.860 105.520 ;
        RECT 292.030 105.180 293.170 105.350 ;
        RECT 289.600 103.960 289.870 104.865 ;
        RECT 290.055 104.720 290.720 104.890 ;
        RECT 290.040 103.790 290.370 104.550 ;
        RECT 290.550 103.960 290.720 104.720 ;
        RECT 290.980 103.790 291.270 104.955 ;
        RECT 291.455 104.840 292.210 105.010 ;
        RECT 291.495 103.790 291.780 104.660 ;
        RECT 291.950 104.590 292.210 104.840 ;
        RECT 293.000 104.930 293.170 105.180 ;
        RECT 293.340 105.100 293.690 105.670 ;
        RECT 293.860 104.930 294.030 105.840 ;
        RECT 294.290 105.790 294.460 106.170 ;
        RECT 294.675 105.960 295.005 106.340 ;
        RECT 294.290 105.620 295.005 105.790 ;
        RECT 294.200 105.070 294.555 105.440 ;
        RECT 294.835 105.430 295.005 105.620 ;
        RECT 295.175 105.595 295.430 106.170 ;
        RECT 294.835 105.100 295.090 105.430 ;
        RECT 293.000 104.760 294.030 104.930 ;
        RECT 294.835 104.890 295.005 105.100 ;
        RECT 291.950 104.420 293.070 104.590 ;
        RECT 291.950 103.960 292.210 104.420 ;
        RECT 292.385 103.790 292.640 104.250 ;
        RECT 292.810 103.960 293.070 104.420 ;
        RECT 293.240 103.790 293.550 104.590 ;
        RECT 293.720 103.960 294.030 104.760 ;
        RECT 294.290 104.720 295.005 104.890 ;
        RECT 295.260 104.865 295.430 105.595 ;
        RECT 295.605 105.500 295.865 106.340 ;
        RECT 297.020 105.860 297.300 106.340 ;
        RECT 297.470 105.690 297.730 106.080 ;
        RECT 297.905 105.860 298.160 106.340 ;
        RECT 298.330 105.690 298.625 106.080 ;
        RECT 298.805 105.860 299.080 106.340 ;
        RECT 299.250 105.840 299.550 106.170 ;
        RECT 296.975 105.520 298.625 105.690 ;
        RECT 296.975 105.010 297.380 105.520 ;
        RECT 297.550 105.180 298.690 105.350 ;
        RECT 294.290 103.960 294.460 104.720 ;
        RECT 294.675 103.790 295.005 104.550 ;
        RECT 295.175 103.960 295.430 104.865 ;
        RECT 295.605 103.790 295.865 104.940 ;
        RECT 296.975 104.840 297.730 105.010 ;
        RECT 297.015 103.790 297.300 104.660 ;
        RECT 297.470 104.590 297.730 104.840 ;
        RECT 298.520 104.930 298.690 105.180 ;
        RECT 298.860 105.100 299.210 105.670 ;
        RECT 299.380 104.930 299.550 105.840 ;
        RECT 299.725 105.500 299.985 106.340 ;
        RECT 300.160 105.595 300.415 106.170 ;
        RECT 300.585 105.960 300.915 106.340 ;
        RECT 301.130 105.790 301.300 106.170 ;
        RECT 300.585 105.620 301.300 105.790 ;
        RECT 301.650 105.790 301.820 106.170 ;
        RECT 302.035 105.960 302.365 106.340 ;
        RECT 301.650 105.620 302.365 105.790 ;
        RECT 298.520 104.760 299.550 104.930 ;
        RECT 297.470 104.420 298.590 104.590 ;
        RECT 297.470 103.960 297.730 104.420 ;
        RECT 297.905 103.790 298.160 104.250 ;
        RECT 298.330 103.960 298.590 104.420 ;
        RECT 298.760 103.790 299.070 104.590 ;
        RECT 299.240 103.960 299.550 104.760 ;
        RECT 299.725 103.790 299.985 104.940 ;
        RECT 300.160 104.865 300.330 105.595 ;
        RECT 300.585 105.430 300.755 105.620 ;
        RECT 300.500 105.100 300.755 105.430 ;
        RECT 300.585 104.890 300.755 105.100 ;
        RECT 301.035 105.070 301.390 105.440 ;
        RECT 301.560 105.070 301.915 105.440 ;
        RECT 302.195 105.430 302.365 105.620 ;
        RECT 302.535 105.595 302.790 106.170 ;
        RECT 302.195 105.100 302.450 105.430 ;
        RECT 302.195 104.890 302.365 105.100 ;
        RECT 300.160 103.960 300.415 104.865 ;
        RECT 300.585 104.720 301.300 104.890 ;
        RECT 300.585 103.790 300.915 104.550 ;
        RECT 301.130 103.960 301.300 104.720 ;
        RECT 301.650 104.720 302.365 104.890 ;
        RECT 302.620 104.865 302.790 105.595 ;
        RECT 302.965 105.500 303.225 106.340 ;
        RECT 303.860 105.615 304.150 106.340 ;
        RECT 304.320 105.840 304.620 106.170 ;
        RECT 304.790 105.860 305.065 106.340 ;
        RECT 301.650 103.960 301.820 104.720 ;
        RECT 302.035 103.790 302.365 104.550 ;
        RECT 302.535 103.960 302.790 104.865 ;
        RECT 302.965 103.790 303.225 104.940 ;
        RECT 303.860 103.790 304.150 104.955 ;
        RECT 304.320 104.930 304.490 105.840 ;
        RECT 305.245 105.690 305.540 106.080 ;
        RECT 305.710 105.860 305.965 106.340 ;
        RECT 306.140 105.690 306.400 106.080 ;
        RECT 306.570 105.860 306.850 106.340 ;
        RECT 304.660 105.100 305.010 105.670 ;
        RECT 305.245 105.520 306.895 105.690 ;
        RECT 305.180 105.180 306.320 105.350 ;
        RECT 305.180 104.930 305.350 105.180 ;
        RECT 306.490 105.010 306.895 105.520 ;
        RECT 307.085 105.500 307.345 106.340 ;
        RECT 307.520 105.595 307.775 106.170 ;
        RECT 307.945 105.960 308.275 106.340 ;
        RECT 308.490 105.790 308.660 106.170 ;
        RECT 307.945 105.620 308.660 105.790 ;
        RECT 304.320 104.760 305.350 104.930 ;
        RECT 306.140 104.840 306.895 105.010 ;
        RECT 304.320 103.960 304.630 104.760 ;
        RECT 306.140 104.590 306.400 104.840 ;
        RECT 304.800 103.790 305.110 104.590 ;
        RECT 305.280 104.420 306.400 104.590 ;
        RECT 305.280 103.960 305.540 104.420 ;
        RECT 305.710 103.790 305.965 104.250 ;
        RECT 306.140 103.960 306.400 104.420 ;
        RECT 306.570 103.790 306.855 104.660 ;
        RECT 307.085 103.790 307.345 104.940 ;
        RECT 307.520 104.865 307.690 105.595 ;
        RECT 307.945 105.430 308.115 105.620 ;
        RECT 309.840 105.590 311.050 106.340 ;
        RECT 307.860 105.100 308.115 105.430 ;
        RECT 307.945 104.890 308.115 105.100 ;
        RECT 308.395 105.070 308.750 105.440 ;
        RECT 307.520 103.960 307.775 104.865 ;
        RECT 307.945 104.720 308.660 104.890 ;
        RECT 307.945 103.790 308.275 104.550 ;
        RECT 308.490 103.960 308.660 104.720 ;
        RECT 309.840 104.880 310.360 105.420 ;
        RECT 310.530 105.050 311.050 105.590 ;
        RECT 309.840 103.790 311.050 104.880 ;
        RECT 162.095 103.620 311.135 103.790 ;
        RECT 162.180 102.530 163.390 103.620 ;
        RECT 163.560 102.530 165.230 103.620 ;
        RECT 165.405 102.950 165.660 103.450 ;
        RECT 165.830 103.120 166.160 103.620 ;
        RECT 165.405 102.780 166.155 102.950 ;
        RECT 162.180 101.820 162.700 102.360 ;
        RECT 162.870 101.990 163.390 102.530 ;
        RECT 163.560 101.840 164.310 102.360 ;
        RECT 164.480 102.010 165.230 102.530 ;
        RECT 165.405 101.960 165.755 102.610 ;
        RECT 162.180 101.070 163.390 101.820 ;
        RECT 163.560 101.070 165.230 101.840 ;
        RECT 165.925 101.790 166.155 102.780 ;
        RECT 165.405 101.620 166.155 101.790 ;
        RECT 165.405 101.330 165.660 101.620 ;
        RECT 165.830 101.070 166.160 101.450 ;
        RECT 166.330 101.330 166.500 103.450 ;
        RECT 166.670 102.650 166.995 103.435 ;
        RECT 167.165 103.160 167.415 103.620 ;
        RECT 167.585 103.120 167.835 103.450 ;
        RECT 168.050 103.120 168.730 103.450 ;
        RECT 167.585 102.990 167.755 103.120 ;
        RECT 167.360 102.820 167.755 102.990 ;
        RECT 166.730 101.600 167.190 102.650 ;
        RECT 167.360 101.460 167.530 102.820 ;
        RECT 167.925 102.560 168.390 102.950 ;
        RECT 167.700 101.750 168.050 102.370 ;
        RECT 168.220 101.970 168.390 102.560 ;
        RECT 168.560 102.340 168.730 103.120 ;
        RECT 168.900 103.020 169.070 103.360 ;
        RECT 169.305 103.190 169.635 103.620 ;
        RECT 169.805 103.020 169.975 103.360 ;
        RECT 170.270 103.160 170.640 103.620 ;
        RECT 168.900 102.850 169.975 103.020 ;
        RECT 170.810 102.990 170.980 103.450 ;
        RECT 171.215 103.110 172.085 103.450 ;
        RECT 172.255 103.160 172.505 103.620 ;
        RECT 170.420 102.820 170.980 102.990 ;
        RECT 170.420 102.680 170.590 102.820 ;
        RECT 169.090 102.510 170.590 102.680 ;
        RECT 171.285 102.650 171.745 102.940 ;
        RECT 168.560 102.170 170.250 102.340 ;
        RECT 168.220 101.750 168.575 101.970 ;
        RECT 168.745 101.460 168.915 102.170 ;
        RECT 169.120 101.750 169.910 102.000 ;
        RECT 170.080 101.990 170.250 102.170 ;
        RECT 170.420 101.820 170.590 102.510 ;
        RECT 166.860 101.070 167.190 101.430 ;
        RECT 167.360 101.290 167.855 101.460 ;
        RECT 168.060 101.290 168.915 101.460 ;
        RECT 169.790 101.070 170.120 101.530 ;
        RECT 170.330 101.430 170.590 101.820 ;
        RECT 170.780 102.640 171.745 102.650 ;
        RECT 171.915 102.730 172.085 103.110 ;
        RECT 172.675 103.070 172.845 103.360 ;
        RECT 173.025 103.240 173.355 103.620 ;
        RECT 172.675 102.900 173.475 103.070 ;
        RECT 170.780 102.480 171.455 102.640 ;
        RECT 171.915 102.560 173.135 102.730 ;
        RECT 170.780 101.690 170.990 102.480 ;
        RECT 171.915 102.470 172.085 102.560 ;
        RECT 171.160 101.690 171.510 102.310 ;
        RECT 171.680 102.300 172.085 102.470 ;
        RECT 171.680 101.520 171.850 102.300 ;
        RECT 172.020 101.850 172.240 102.130 ;
        RECT 172.420 102.020 172.960 102.390 ;
        RECT 173.305 102.310 173.475 102.900 ;
        RECT 173.695 102.480 174.000 103.620 ;
        RECT 174.170 102.430 174.420 103.310 ;
        RECT 174.590 102.480 174.840 103.620 ;
        RECT 175.060 102.455 175.350 103.620 ;
        RECT 175.525 102.480 175.860 103.450 ;
        RECT 176.030 102.480 176.200 103.620 ;
        RECT 176.370 103.280 178.400 103.450 ;
        RECT 173.305 102.280 174.045 102.310 ;
        RECT 172.020 101.680 172.550 101.850 ;
        RECT 170.330 101.260 170.680 101.430 ;
        RECT 170.900 101.240 171.850 101.520 ;
        RECT 172.020 101.070 172.210 101.510 ;
        RECT 172.380 101.450 172.550 101.680 ;
        RECT 172.720 101.620 172.960 102.020 ;
        RECT 173.130 101.980 174.045 102.280 ;
        RECT 173.130 101.805 173.455 101.980 ;
        RECT 173.130 101.450 173.450 101.805 ;
        RECT 174.215 101.780 174.420 102.430 ;
        RECT 172.380 101.280 173.450 101.450 ;
        RECT 173.695 101.070 174.000 101.530 ;
        RECT 174.170 101.250 174.420 101.780 ;
        RECT 174.590 101.070 174.840 101.825 ;
        RECT 175.525 101.810 175.695 102.480 ;
        RECT 176.370 102.310 176.540 103.280 ;
        RECT 175.865 101.980 176.120 102.310 ;
        RECT 176.345 101.980 176.540 102.310 ;
        RECT 176.710 102.940 177.835 103.110 ;
        RECT 175.950 101.810 176.120 101.980 ;
        RECT 176.710 101.810 176.880 102.940 ;
        RECT 175.060 101.070 175.350 101.795 ;
        RECT 175.525 101.240 175.780 101.810 ;
        RECT 175.950 101.640 176.880 101.810 ;
        RECT 177.050 102.600 178.060 102.770 ;
        RECT 177.050 101.800 177.220 102.600 ;
        RECT 177.425 102.260 177.700 102.400 ;
        RECT 177.420 102.090 177.700 102.260 ;
        RECT 176.705 101.605 176.880 101.640 ;
        RECT 175.950 101.070 176.280 101.470 ;
        RECT 176.705 101.240 177.235 101.605 ;
        RECT 177.425 101.240 177.700 102.090 ;
        RECT 177.870 101.240 178.060 102.600 ;
        RECT 178.230 102.615 178.400 103.280 ;
        RECT 178.570 102.860 178.740 103.620 ;
        RECT 178.975 102.860 179.490 103.270 ;
        RECT 178.230 102.425 178.980 102.615 ;
        RECT 179.150 102.050 179.490 102.860 ;
        RECT 179.665 102.470 179.925 103.620 ;
        RECT 180.100 102.545 180.355 103.450 ;
        RECT 180.525 102.860 180.855 103.620 ;
        RECT 181.070 102.690 181.240 103.450 ;
        RECT 181.505 102.950 181.760 103.450 ;
        RECT 181.930 103.120 182.260 103.620 ;
        RECT 181.505 102.780 182.255 102.950 ;
        RECT 178.260 101.880 179.490 102.050 ;
        RECT 178.240 101.070 178.750 101.605 ;
        RECT 178.970 101.275 179.215 101.880 ;
        RECT 179.665 101.070 179.925 101.910 ;
        RECT 180.100 101.815 180.270 102.545 ;
        RECT 180.525 102.520 181.240 102.690 ;
        RECT 180.525 102.310 180.695 102.520 ;
        RECT 180.440 101.980 180.695 102.310 ;
        RECT 180.100 101.240 180.355 101.815 ;
        RECT 180.525 101.790 180.695 101.980 ;
        RECT 180.975 101.970 181.330 102.340 ;
        RECT 181.505 101.960 181.855 102.610 ;
        RECT 182.025 101.790 182.255 102.780 ;
        RECT 180.525 101.620 181.240 101.790 ;
        RECT 180.525 101.070 180.855 101.450 ;
        RECT 181.070 101.240 181.240 101.620 ;
        RECT 181.505 101.620 182.255 101.790 ;
        RECT 181.505 101.330 181.760 101.620 ;
        RECT 181.930 101.070 182.260 101.450 ;
        RECT 182.430 101.330 182.600 103.450 ;
        RECT 182.770 102.650 183.095 103.435 ;
        RECT 183.265 103.160 183.515 103.620 ;
        RECT 183.685 103.120 183.935 103.450 ;
        RECT 184.150 103.120 184.830 103.450 ;
        RECT 183.685 102.990 183.855 103.120 ;
        RECT 183.460 102.820 183.855 102.990 ;
        RECT 182.830 101.600 183.290 102.650 ;
        RECT 183.460 101.460 183.630 102.820 ;
        RECT 184.025 102.560 184.490 102.950 ;
        RECT 183.800 101.750 184.150 102.370 ;
        RECT 184.320 101.970 184.490 102.560 ;
        RECT 184.660 102.340 184.830 103.120 ;
        RECT 185.000 103.020 185.170 103.360 ;
        RECT 185.405 103.190 185.735 103.620 ;
        RECT 185.905 103.020 186.075 103.360 ;
        RECT 186.370 103.160 186.740 103.620 ;
        RECT 185.000 102.850 186.075 103.020 ;
        RECT 186.910 102.990 187.080 103.450 ;
        RECT 187.315 103.110 188.185 103.450 ;
        RECT 188.355 103.160 188.605 103.620 ;
        RECT 186.520 102.820 187.080 102.990 ;
        RECT 186.520 102.680 186.690 102.820 ;
        RECT 185.190 102.510 186.690 102.680 ;
        RECT 187.385 102.650 187.845 102.940 ;
        RECT 184.660 102.170 186.350 102.340 ;
        RECT 184.320 101.750 184.675 101.970 ;
        RECT 184.845 101.460 185.015 102.170 ;
        RECT 185.220 101.750 186.010 102.000 ;
        RECT 186.180 101.990 186.350 102.170 ;
        RECT 186.520 101.820 186.690 102.510 ;
        RECT 182.960 101.070 183.290 101.430 ;
        RECT 183.460 101.290 183.955 101.460 ;
        RECT 184.160 101.290 185.015 101.460 ;
        RECT 185.890 101.070 186.220 101.530 ;
        RECT 186.430 101.430 186.690 101.820 ;
        RECT 186.880 102.640 187.845 102.650 ;
        RECT 188.015 102.730 188.185 103.110 ;
        RECT 188.775 103.070 188.945 103.360 ;
        RECT 189.125 103.240 189.455 103.620 ;
        RECT 188.775 102.900 189.575 103.070 ;
        RECT 186.880 102.480 187.555 102.640 ;
        RECT 188.015 102.560 189.235 102.730 ;
        RECT 186.880 101.690 187.090 102.480 ;
        RECT 188.015 102.470 188.185 102.560 ;
        RECT 187.260 101.690 187.610 102.310 ;
        RECT 187.780 102.300 188.185 102.470 ;
        RECT 187.780 101.520 187.950 102.300 ;
        RECT 188.120 101.850 188.340 102.130 ;
        RECT 188.520 102.020 189.060 102.390 ;
        RECT 189.405 102.310 189.575 102.900 ;
        RECT 189.795 102.480 190.100 103.620 ;
        RECT 190.270 102.430 190.520 103.310 ;
        RECT 190.690 102.480 190.940 103.620 ;
        RECT 191.165 102.950 191.420 103.450 ;
        RECT 191.590 103.120 191.920 103.620 ;
        RECT 191.165 102.780 191.915 102.950 ;
        RECT 189.405 102.280 190.145 102.310 ;
        RECT 188.120 101.680 188.650 101.850 ;
        RECT 186.430 101.260 186.780 101.430 ;
        RECT 187.000 101.240 187.950 101.520 ;
        RECT 188.120 101.070 188.310 101.510 ;
        RECT 188.480 101.450 188.650 101.680 ;
        RECT 188.820 101.620 189.060 102.020 ;
        RECT 189.230 101.980 190.145 102.280 ;
        RECT 189.230 101.805 189.555 101.980 ;
        RECT 189.230 101.450 189.550 101.805 ;
        RECT 190.315 101.780 190.520 102.430 ;
        RECT 191.165 101.960 191.515 102.610 ;
        RECT 188.480 101.280 189.550 101.450 ;
        RECT 189.795 101.070 190.100 101.530 ;
        RECT 190.270 101.250 190.520 101.780 ;
        RECT 190.690 101.070 190.940 101.825 ;
        RECT 191.685 101.790 191.915 102.780 ;
        RECT 191.165 101.620 191.915 101.790 ;
        RECT 191.165 101.330 191.420 101.620 ;
        RECT 191.590 101.070 191.920 101.450 ;
        RECT 192.090 101.330 192.260 103.450 ;
        RECT 192.430 102.650 192.755 103.435 ;
        RECT 192.925 103.160 193.175 103.620 ;
        RECT 193.345 103.120 193.595 103.450 ;
        RECT 193.810 103.120 194.490 103.450 ;
        RECT 193.345 102.990 193.515 103.120 ;
        RECT 193.120 102.820 193.515 102.990 ;
        RECT 192.490 101.600 192.950 102.650 ;
        RECT 193.120 101.460 193.290 102.820 ;
        RECT 193.685 102.560 194.150 102.950 ;
        RECT 193.460 101.750 193.810 102.370 ;
        RECT 193.980 101.970 194.150 102.560 ;
        RECT 194.320 102.340 194.490 103.120 ;
        RECT 194.660 103.020 194.830 103.360 ;
        RECT 195.065 103.190 195.395 103.620 ;
        RECT 195.565 103.020 195.735 103.360 ;
        RECT 196.030 103.160 196.400 103.620 ;
        RECT 194.660 102.850 195.735 103.020 ;
        RECT 196.570 102.990 196.740 103.450 ;
        RECT 196.975 103.110 197.845 103.450 ;
        RECT 198.015 103.160 198.265 103.620 ;
        RECT 196.180 102.820 196.740 102.990 ;
        RECT 196.180 102.680 196.350 102.820 ;
        RECT 194.850 102.510 196.350 102.680 ;
        RECT 197.045 102.650 197.505 102.940 ;
        RECT 194.320 102.170 196.010 102.340 ;
        RECT 193.980 101.750 194.335 101.970 ;
        RECT 194.505 101.460 194.675 102.170 ;
        RECT 194.880 101.750 195.670 102.000 ;
        RECT 195.840 101.990 196.010 102.170 ;
        RECT 196.180 101.820 196.350 102.510 ;
        RECT 192.620 101.070 192.950 101.430 ;
        RECT 193.120 101.290 193.615 101.460 ;
        RECT 193.820 101.290 194.675 101.460 ;
        RECT 195.550 101.070 195.880 101.530 ;
        RECT 196.090 101.430 196.350 101.820 ;
        RECT 196.540 102.640 197.505 102.650 ;
        RECT 197.675 102.730 197.845 103.110 ;
        RECT 198.435 103.070 198.605 103.360 ;
        RECT 198.785 103.240 199.115 103.620 ;
        RECT 198.435 102.900 199.235 103.070 ;
        RECT 196.540 102.480 197.215 102.640 ;
        RECT 197.675 102.560 198.895 102.730 ;
        RECT 196.540 101.690 196.750 102.480 ;
        RECT 197.675 102.470 197.845 102.560 ;
        RECT 196.920 101.690 197.270 102.310 ;
        RECT 197.440 102.300 197.845 102.470 ;
        RECT 197.440 101.520 197.610 102.300 ;
        RECT 197.780 101.850 198.000 102.130 ;
        RECT 198.180 102.020 198.720 102.390 ;
        RECT 199.065 102.310 199.235 102.900 ;
        RECT 199.455 102.480 199.760 103.620 ;
        RECT 199.930 102.430 200.180 103.310 ;
        RECT 200.350 102.480 200.600 103.620 ;
        RECT 200.820 102.455 201.110 103.620 ;
        RECT 201.830 102.690 202.000 103.450 ;
        RECT 202.180 102.860 202.510 103.620 ;
        RECT 201.830 102.520 202.495 102.690 ;
        RECT 202.680 102.545 202.950 103.450 ;
        RECT 199.065 102.280 199.805 102.310 ;
        RECT 197.780 101.680 198.310 101.850 ;
        RECT 196.090 101.260 196.440 101.430 ;
        RECT 196.660 101.240 197.610 101.520 ;
        RECT 197.780 101.070 197.970 101.510 ;
        RECT 198.140 101.450 198.310 101.680 ;
        RECT 198.480 101.620 198.720 102.020 ;
        RECT 198.890 101.980 199.805 102.280 ;
        RECT 198.890 101.805 199.215 101.980 ;
        RECT 198.890 101.450 199.210 101.805 ;
        RECT 199.975 101.780 200.180 102.430 ;
        RECT 202.325 102.375 202.495 102.520 ;
        RECT 201.760 101.970 202.090 102.340 ;
        RECT 202.325 102.045 202.610 102.375 ;
        RECT 198.140 101.280 199.210 101.450 ;
        RECT 199.455 101.070 199.760 101.530 ;
        RECT 199.930 101.250 200.180 101.780 ;
        RECT 200.350 101.070 200.600 101.825 ;
        RECT 200.820 101.070 201.110 101.795 ;
        RECT 202.325 101.790 202.495 102.045 ;
        RECT 201.830 101.620 202.495 101.790 ;
        RECT 202.780 101.745 202.950 102.545 ;
        RECT 203.210 102.690 203.380 103.450 ;
        RECT 203.595 102.860 203.925 103.620 ;
        RECT 203.210 102.520 203.925 102.690 ;
        RECT 204.095 102.545 204.350 103.450 ;
        RECT 203.120 101.970 203.475 102.340 ;
        RECT 203.755 102.310 203.925 102.520 ;
        RECT 203.755 101.980 204.010 102.310 ;
        RECT 203.755 101.790 203.925 101.980 ;
        RECT 204.180 101.815 204.350 102.545 ;
        RECT 204.525 102.470 204.785 103.620 ;
        RECT 205.425 102.950 205.680 103.450 ;
        RECT 205.850 103.120 206.180 103.620 ;
        RECT 205.425 102.780 206.175 102.950 ;
        RECT 205.425 101.960 205.775 102.610 ;
        RECT 201.830 101.240 202.000 101.620 ;
        RECT 202.180 101.070 202.510 101.450 ;
        RECT 202.690 101.240 202.950 101.745 ;
        RECT 203.210 101.620 203.925 101.790 ;
        RECT 203.210 101.240 203.380 101.620 ;
        RECT 203.595 101.070 203.925 101.450 ;
        RECT 204.095 101.240 204.350 101.815 ;
        RECT 204.525 101.070 204.785 101.910 ;
        RECT 205.945 101.790 206.175 102.780 ;
        RECT 205.425 101.620 206.175 101.790 ;
        RECT 205.425 101.330 205.680 101.620 ;
        RECT 205.850 101.070 206.180 101.450 ;
        RECT 206.350 101.330 206.520 103.450 ;
        RECT 206.690 102.650 207.015 103.435 ;
        RECT 207.185 103.160 207.435 103.620 ;
        RECT 207.605 103.120 207.855 103.450 ;
        RECT 208.070 103.120 208.750 103.450 ;
        RECT 207.605 102.990 207.775 103.120 ;
        RECT 207.380 102.820 207.775 102.990 ;
        RECT 206.750 101.600 207.210 102.650 ;
        RECT 207.380 101.460 207.550 102.820 ;
        RECT 207.945 102.560 208.410 102.950 ;
        RECT 207.720 101.750 208.070 102.370 ;
        RECT 208.240 101.970 208.410 102.560 ;
        RECT 208.580 102.340 208.750 103.120 ;
        RECT 208.920 103.020 209.090 103.360 ;
        RECT 209.325 103.190 209.655 103.620 ;
        RECT 209.825 103.020 209.995 103.360 ;
        RECT 210.290 103.160 210.660 103.620 ;
        RECT 208.920 102.850 209.995 103.020 ;
        RECT 210.830 102.990 211.000 103.450 ;
        RECT 211.235 103.110 212.105 103.450 ;
        RECT 212.275 103.160 212.525 103.620 ;
        RECT 210.440 102.820 211.000 102.990 ;
        RECT 210.440 102.680 210.610 102.820 ;
        RECT 209.110 102.510 210.610 102.680 ;
        RECT 211.305 102.650 211.765 102.940 ;
        RECT 208.580 102.170 210.270 102.340 ;
        RECT 208.240 101.750 208.595 101.970 ;
        RECT 208.765 101.460 208.935 102.170 ;
        RECT 209.140 101.750 209.930 102.000 ;
        RECT 210.100 101.990 210.270 102.170 ;
        RECT 210.440 101.820 210.610 102.510 ;
        RECT 206.880 101.070 207.210 101.430 ;
        RECT 207.380 101.290 207.875 101.460 ;
        RECT 208.080 101.290 208.935 101.460 ;
        RECT 209.810 101.070 210.140 101.530 ;
        RECT 210.350 101.430 210.610 101.820 ;
        RECT 210.800 102.640 211.765 102.650 ;
        RECT 211.935 102.730 212.105 103.110 ;
        RECT 212.695 103.070 212.865 103.360 ;
        RECT 213.045 103.240 213.375 103.620 ;
        RECT 212.695 102.900 213.495 103.070 ;
        RECT 210.800 102.480 211.475 102.640 ;
        RECT 211.935 102.560 213.155 102.730 ;
        RECT 210.800 101.690 211.010 102.480 ;
        RECT 211.935 102.470 212.105 102.560 ;
        RECT 211.180 101.690 211.530 102.310 ;
        RECT 211.700 102.300 212.105 102.470 ;
        RECT 211.700 101.520 211.870 102.300 ;
        RECT 212.040 101.850 212.260 102.130 ;
        RECT 212.440 102.020 212.980 102.390 ;
        RECT 213.325 102.310 213.495 102.900 ;
        RECT 213.715 102.480 214.020 103.620 ;
        RECT 214.190 102.430 214.445 103.310 ;
        RECT 214.675 102.750 214.960 103.620 ;
        RECT 215.130 102.990 215.390 103.450 ;
        RECT 215.565 103.160 215.820 103.620 ;
        RECT 215.990 102.990 216.250 103.450 ;
        RECT 215.130 102.820 216.250 102.990 ;
        RECT 216.420 102.820 216.730 103.620 ;
        RECT 215.130 102.570 215.390 102.820 ;
        RECT 216.900 102.650 217.210 103.450 ;
        RECT 217.385 102.950 217.640 103.450 ;
        RECT 217.810 103.120 218.140 103.620 ;
        RECT 217.385 102.780 218.135 102.950 ;
        RECT 213.325 102.280 214.065 102.310 ;
        RECT 212.040 101.680 212.570 101.850 ;
        RECT 210.350 101.260 210.700 101.430 ;
        RECT 210.920 101.240 211.870 101.520 ;
        RECT 212.040 101.070 212.230 101.510 ;
        RECT 212.400 101.450 212.570 101.680 ;
        RECT 212.740 101.620 212.980 102.020 ;
        RECT 213.150 101.980 214.065 102.280 ;
        RECT 213.150 101.805 213.475 101.980 ;
        RECT 213.150 101.450 213.470 101.805 ;
        RECT 214.235 101.780 214.445 102.430 ;
        RECT 212.400 101.280 213.470 101.450 ;
        RECT 213.715 101.070 214.020 101.530 ;
        RECT 214.190 101.250 214.445 101.780 ;
        RECT 214.635 102.400 215.390 102.570 ;
        RECT 216.180 102.480 217.210 102.650 ;
        RECT 214.635 101.890 215.040 102.400 ;
        RECT 216.180 102.230 216.350 102.480 ;
        RECT 215.210 102.060 216.350 102.230 ;
        RECT 214.635 101.720 216.285 101.890 ;
        RECT 216.520 101.740 216.870 102.310 ;
        RECT 214.680 101.070 214.960 101.550 ;
        RECT 215.130 101.330 215.390 101.720 ;
        RECT 215.565 101.070 215.820 101.550 ;
        RECT 215.990 101.330 216.285 101.720 ;
        RECT 217.040 101.570 217.210 102.480 ;
        RECT 217.385 101.960 217.735 102.610 ;
        RECT 217.905 101.790 218.135 102.780 ;
        RECT 216.465 101.070 216.740 101.550 ;
        RECT 216.910 101.240 217.210 101.570 ;
        RECT 217.385 101.620 218.135 101.790 ;
        RECT 217.385 101.330 217.640 101.620 ;
        RECT 217.810 101.070 218.140 101.450 ;
        RECT 218.310 101.330 218.480 103.450 ;
        RECT 218.650 102.650 218.975 103.435 ;
        RECT 219.145 103.160 219.395 103.620 ;
        RECT 219.565 103.120 219.815 103.450 ;
        RECT 220.030 103.120 220.710 103.450 ;
        RECT 219.565 102.990 219.735 103.120 ;
        RECT 219.340 102.820 219.735 102.990 ;
        RECT 218.710 101.600 219.170 102.650 ;
        RECT 219.340 101.460 219.510 102.820 ;
        RECT 219.905 102.560 220.370 102.950 ;
        RECT 219.680 101.750 220.030 102.370 ;
        RECT 220.200 101.970 220.370 102.560 ;
        RECT 220.540 102.340 220.710 103.120 ;
        RECT 220.880 103.020 221.050 103.360 ;
        RECT 221.285 103.190 221.615 103.620 ;
        RECT 221.785 103.020 221.955 103.360 ;
        RECT 222.250 103.160 222.620 103.620 ;
        RECT 220.880 102.850 221.955 103.020 ;
        RECT 222.790 102.990 222.960 103.450 ;
        RECT 223.195 103.110 224.065 103.450 ;
        RECT 224.235 103.160 224.485 103.620 ;
        RECT 222.400 102.820 222.960 102.990 ;
        RECT 222.400 102.680 222.570 102.820 ;
        RECT 221.070 102.510 222.570 102.680 ;
        RECT 223.265 102.650 223.725 102.940 ;
        RECT 220.540 102.170 222.230 102.340 ;
        RECT 220.200 101.750 220.555 101.970 ;
        RECT 220.725 101.460 220.895 102.170 ;
        RECT 221.100 101.750 221.890 102.000 ;
        RECT 222.060 101.990 222.230 102.170 ;
        RECT 222.400 101.820 222.570 102.510 ;
        RECT 218.840 101.070 219.170 101.430 ;
        RECT 219.340 101.290 219.835 101.460 ;
        RECT 220.040 101.290 220.895 101.460 ;
        RECT 221.770 101.070 222.100 101.530 ;
        RECT 222.310 101.430 222.570 101.820 ;
        RECT 222.760 102.640 223.725 102.650 ;
        RECT 223.895 102.730 224.065 103.110 ;
        RECT 224.655 103.070 224.825 103.360 ;
        RECT 225.005 103.240 225.335 103.620 ;
        RECT 224.655 102.900 225.455 103.070 ;
        RECT 222.760 102.480 223.435 102.640 ;
        RECT 223.895 102.560 225.115 102.730 ;
        RECT 222.760 101.690 222.970 102.480 ;
        RECT 223.895 102.470 224.065 102.560 ;
        RECT 223.140 101.690 223.490 102.310 ;
        RECT 223.660 102.300 224.065 102.470 ;
        RECT 223.660 101.520 223.830 102.300 ;
        RECT 224.000 101.850 224.220 102.130 ;
        RECT 224.400 102.020 224.940 102.390 ;
        RECT 225.285 102.310 225.455 102.900 ;
        RECT 225.675 102.480 225.980 103.620 ;
        RECT 226.150 102.430 226.405 103.310 ;
        RECT 226.580 102.455 226.870 103.620 ;
        RECT 227.045 102.950 227.300 103.450 ;
        RECT 227.470 103.120 227.800 103.620 ;
        RECT 227.045 102.780 227.795 102.950 ;
        RECT 225.285 102.280 226.025 102.310 ;
        RECT 224.000 101.680 224.530 101.850 ;
        RECT 222.310 101.260 222.660 101.430 ;
        RECT 222.880 101.240 223.830 101.520 ;
        RECT 224.000 101.070 224.190 101.510 ;
        RECT 224.360 101.450 224.530 101.680 ;
        RECT 224.700 101.620 224.940 102.020 ;
        RECT 225.110 101.980 226.025 102.280 ;
        RECT 225.110 101.805 225.435 101.980 ;
        RECT 225.110 101.450 225.430 101.805 ;
        RECT 226.195 101.780 226.405 102.430 ;
        RECT 227.045 101.960 227.395 102.610 ;
        RECT 224.360 101.280 225.430 101.450 ;
        RECT 225.675 101.070 225.980 101.530 ;
        RECT 226.150 101.250 226.405 101.780 ;
        RECT 226.580 101.070 226.870 101.795 ;
        RECT 227.565 101.790 227.795 102.780 ;
        RECT 227.045 101.620 227.795 101.790 ;
        RECT 227.045 101.330 227.300 101.620 ;
        RECT 227.470 101.070 227.800 101.450 ;
        RECT 227.970 101.330 228.140 103.450 ;
        RECT 228.310 102.650 228.635 103.435 ;
        RECT 228.805 103.160 229.055 103.620 ;
        RECT 229.225 103.120 229.475 103.450 ;
        RECT 229.690 103.120 230.370 103.450 ;
        RECT 229.225 102.990 229.395 103.120 ;
        RECT 229.000 102.820 229.395 102.990 ;
        RECT 228.370 101.600 228.830 102.650 ;
        RECT 229.000 101.460 229.170 102.820 ;
        RECT 229.565 102.560 230.030 102.950 ;
        RECT 229.340 101.750 229.690 102.370 ;
        RECT 229.860 101.970 230.030 102.560 ;
        RECT 230.200 102.340 230.370 103.120 ;
        RECT 230.540 103.020 230.710 103.360 ;
        RECT 230.945 103.190 231.275 103.620 ;
        RECT 231.445 103.020 231.615 103.360 ;
        RECT 231.910 103.160 232.280 103.620 ;
        RECT 230.540 102.850 231.615 103.020 ;
        RECT 232.450 102.990 232.620 103.450 ;
        RECT 232.855 103.110 233.725 103.450 ;
        RECT 233.895 103.160 234.145 103.620 ;
        RECT 232.060 102.820 232.620 102.990 ;
        RECT 232.060 102.680 232.230 102.820 ;
        RECT 230.730 102.510 232.230 102.680 ;
        RECT 232.925 102.650 233.385 102.940 ;
        RECT 230.200 102.170 231.890 102.340 ;
        RECT 229.860 101.750 230.215 101.970 ;
        RECT 230.385 101.460 230.555 102.170 ;
        RECT 230.760 101.750 231.550 102.000 ;
        RECT 231.720 101.990 231.890 102.170 ;
        RECT 232.060 101.820 232.230 102.510 ;
        RECT 228.500 101.070 228.830 101.430 ;
        RECT 229.000 101.290 229.495 101.460 ;
        RECT 229.700 101.290 230.555 101.460 ;
        RECT 231.430 101.070 231.760 101.530 ;
        RECT 231.970 101.430 232.230 101.820 ;
        RECT 232.420 102.640 233.385 102.650 ;
        RECT 233.555 102.730 233.725 103.110 ;
        RECT 234.315 103.070 234.485 103.360 ;
        RECT 234.665 103.240 234.995 103.620 ;
        RECT 234.315 102.900 235.115 103.070 ;
        RECT 232.420 102.480 233.095 102.640 ;
        RECT 233.555 102.560 234.775 102.730 ;
        RECT 232.420 101.690 232.630 102.480 ;
        RECT 233.555 102.470 233.725 102.560 ;
        RECT 232.800 101.690 233.150 102.310 ;
        RECT 233.320 102.300 233.725 102.470 ;
        RECT 233.320 101.520 233.490 102.300 ;
        RECT 233.660 101.850 233.880 102.130 ;
        RECT 234.060 102.020 234.600 102.390 ;
        RECT 234.945 102.310 235.115 102.900 ;
        RECT 235.335 102.480 235.640 103.620 ;
        RECT 235.810 102.430 236.065 103.310 ;
        RECT 236.245 102.470 236.505 103.620 ;
        RECT 236.680 102.545 236.935 103.450 ;
        RECT 237.105 102.860 237.435 103.620 ;
        RECT 237.650 102.690 237.820 103.450 ;
        RECT 238.545 102.950 238.800 103.450 ;
        RECT 238.970 103.120 239.300 103.620 ;
        RECT 238.545 102.780 239.295 102.950 ;
        RECT 234.945 102.280 235.685 102.310 ;
        RECT 233.660 101.680 234.190 101.850 ;
        RECT 231.970 101.260 232.320 101.430 ;
        RECT 232.540 101.240 233.490 101.520 ;
        RECT 233.660 101.070 233.850 101.510 ;
        RECT 234.020 101.450 234.190 101.680 ;
        RECT 234.360 101.620 234.600 102.020 ;
        RECT 234.770 101.980 235.685 102.280 ;
        RECT 234.770 101.805 235.095 101.980 ;
        RECT 234.770 101.450 235.090 101.805 ;
        RECT 235.855 101.780 236.065 102.430 ;
        RECT 234.020 101.280 235.090 101.450 ;
        RECT 235.335 101.070 235.640 101.530 ;
        RECT 235.810 101.250 236.065 101.780 ;
        RECT 236.245 101.070 236.505 101.910 ;
        RECT 236.680 101.815 236.850 102.545 ;
        RECT 237.105 102.520 237.820 102.690 ;
        RECT 237.105 102.310 237.275 102.520 ;
        RECT 237.020 101.980 237.275 102.310 ;
        RECT 236.680 101.240 236.935 101.815 ;
        RECT 237.105 101.790 237.275 101.980 ;
        RECT 237.555 101.970 237.910 102.340 ;
        RECT 238.545 101.960 238.895 102.610 ;
        RECT 239.065 101.790 239.295 102.780 ;
        RECT 237.105 101.620 237.820 101.790 ;
        RECT 237.105 101.070 237.435 101.450 ;
        RECT 237.650 101.240 237.820 101.620 ;
        RECT 238.545 101.620 239.295 101.790 ;
        RECT 238.545 101.330 238.800 101.620 ;
        RECT 238.970 101.070 239.300 101.450 ;
        RECT 239.470 101.330 239.640 103.450 ;
        RECT 239.810 102.650 240.135 103.435 ;
        RECT 240.305 103.160 240.555 103.620 ;
        RECT 240.725 103.120 240.975 103.450 ;
        RECT 241.190 103.120 241.870 103.450 ;
        RECT 240.725 102.990 240.895 103.120 ;
        RECT 240.500 102.820 240.895 102.990 ;
        RECT 239.870 101.600 240.330 102.650 ;
        RECT 240.500 101.460 240.670 102.820 ;
        RECT 241.065 102.560 241.530 102.950 ;
        RECT 240.840 101.750 241.190 102.370 ;
        RECT 241.360 101.970 241.530 102.560 ;
        RECT 241.700 102.340 241.870 103.120 ;
        RECT 242.040 103.020 242.210 103.360 ;
        RECT 242.445 103.190 242.775 103.620 ;
        RECT 242.945 103.020 243.115 103.360 ;
        RECT 243.410 103.160 243.780 103.620 ;
        RECT 242.040 102.850 243.115 103.020 ;
        RECT 243.950 102.990 244.120 103.450 ;
        RECT 244.355 103.110 245.225 103.450 ;
        RECT 245.395 103.160 245.645 103.620 ;
        RECT 243.560 102.820 244.120 102.990 ;
        RECT 243.560 102.680 243.730 102.820 ;
        RECT 242.230 102.510 243.730 102.680 ;
        RECT 244.425 102.650 244.885 102.940 ;
        RECT 241.700 102.170 243.390 102.340 ;
        RECT 241.360 101.750 241.715 101.970 ;
        RECT 241.885 101.460 242.055 102.170 ;
        RECT 242.260 101.750 243.050 102.000 ;
        RECT 243.220 101.990 243.390 102.170 ;
        RECT 243.560 101.820 243.730 102.510 ;
        RECT 240.000 101.070 240.330 101.430 ;
        RECT 240.500 101.290 240.995 101.460 ;
        RECT 241.200 101.290 242.055 101.460 ;
        RECT 242.930 101.070 243.260 101.530 ;
        RECT 243.470 101.430 243.730 101.820 ;
        RECT 243.920 102.640 244.885 102.650 ;
        RECT 245.055 102.730 245.225 103.110 ;
        RECT 245.815 103.070 245.985 103.360 ;
        RECT 246.165 103.240 246.495 103.620 ;
        RECT 245.815 102.900 246.615 103.070 ;
        RECT 243.920 102.480 244.595 102.640 ;
        RECT 245.055 102.560 246.275 102.730 ;
        RECT 243.920 101.690 244.130 102.480 ;
        RECT 245.055 102.470 245.225 102.560 ;
        RECT 244.300 101.690 244.650 102.310 ;
        RECT 244.820 102.300 245.225 102.470 ;
        RECT 244.820 101.520 244.990 102.300 ;
        RECT 245.160 101.850 245.380 102.130 ;
        RECT 245.560 102.020 246.100 102.390 ;
        RECT 246.445 102.310 246.615 102.900 ;
        RECT 246.835 102.480 247.140 103.620 ;
        RECT 247.310 102.430 247.565 103.310 ;
        RECT 247.795 102.750 248.080 103.620 ;
        RECT 248.250 102.990 248.510 103.450 ;
        RECT 248.685 103.160 248.940 103.620 ;
        RECT 249.110 102.990 249.370 103.450 ;
        RECT 248.250 102.820 249.370 102.990 ;
        RECT 249.540 102.820 249.850 103.620 ;
        RECT 248.250 102.570 248.510 102.820 ;
        RECT 250.020 102.650 250.330 103.450 ;
        RECT 246.445 102.280 247.185 102.310 ;
        RECT 245.160 101.680 245.690 101.850 ;
        RECT 243.470 101.260 243.820 101.430 ;
        RECT 244.040 101.240 244.990 101.520 ;
        RECT 245.160 101.070 245.350 101.510 ;
        RECT 245.520 101.450 245.690 101.680 ;
        RECT 245.860 101.620 246.100 102.020 ;
        RECT 246.270 101.980 247.185 102.280 ;
        RECT 246.270 101.805 246.595 101.980 ;
        RECT 246.270 101.450 246.590 101.805 ;
        RECT 247.355 101.780 247.565 102.430 ;
        RECT 245.520 101.280 246.590 101.450 ;
        RECT 246.835 101.070 247.140 101.530 ;
        RECT 247.310 101.250 247.565 101.780 ;
        RECT 247.755 102.400 248.510 102.570 ;
        RECT 249.300 102.480 250.330 102.650 ;
        RECT 247.755 101.890 248.160 102.400 ;
        RECT 249.300 102.230 249.470 102.480 ;
        RECT 248.330 102.060 249.470 102.230 ;
        RECT 247.755 101.720 249.405 101.890 ;
        RECT 249.640 101.740 249.990 102.310 ;
        RECT 247.800 101.070 248.080 101.550 ;
        RECT 248.250 101.330 248.510 101.720 ;
        RECT 248.685 101.070 248.940 101.550 ;
        RECT 249.110 101.330 249.405 101.720 ;
        RECT 250.160 101.570 250.330 102.480 ;
        RECT 249.585 101.070 249.860 101.550 ;
        RECT 250.030 101.240 250.330 101.570 ;
        RECT 250.500 102.545 250.770 103.450 ;
        RECT 250.940 102.860 251.270 103.620 ;
        RECT 251.450 102.690 251.620 103.450 ;
        RECT 250.500 101.745 250.670 102.545 ;
        RECT 250.955 102.520 251.620 102.690 ;
        RECT 250.955 102.375 251.125 102.520 ;
        RECT 252.340 102.455 252.630 103.620 ;
        RECT 252.805 102.470 253.065 103.620 ;
        RECT 253.240 102.545 253.495 103.450 ;
        RECT 253.665 102.860 253.995 103.620 ;
        RECT 254.210 102.690 254.380 103.450 ;
        RECT 250.840 102.045 251.125 102.375 ;
        RECT 250.955 101.790 251.125 102.045 ;
        RECT 251.360 101.970 251.690 102.340 ;
        RECT 250.500 101.240 250.760 101.745 ;
        RECT 250.955 101.620 251.620 101.790 ;
        RECT 250.940 101.070 251.270 101.450 ;
        RECT 251.450 101.240 251.620 101.620 ;
        RECT 252.340 101.070 252.630 101.795 ;
        RECT 252.805 101.070 253.065 101.910 ;
        RECT 253.240 101.815 253.410 102.545 ;
        RECT 253.665 102.520 254.380 102.690 ;
        RECT 255.565 103.230 255.900 103.450 ;
        RECT 256.905 103.240 257.260 103.620 ;
        RECT 255.565 102.610 255.820 103.230 ;
        RECT 256.070 103.070 256.300 103.110 ;
        RECT 257.430 103.070 257.680 103.450 ;
        RECT 256.070 102.870 257.680 103.070 ;
        RECT 256.070 102.780 256.255 102.870 ;
        RECT 256.845 102.860 257.680 102.870 ;
        RECT 257.930 102.840 258.180 103.620 ;
        RECT 258.350 102.770 258.610 103.450 ;
        RECT 256.410 102.670 256.740 102.700 ;
        RECT 256.410 102.610 258.210 102.670 ;
        RECT 253.665 102.310 253.835 102.520 ;
        RECT 255.565 102.500 258.270 102.610 ;
        RECT 255.565 102.440 256.740 102.500 ;
        RECT 258.070 102.465 258.270 102.500 ;
        RECT 253.580 101.980 253.835 102.310 ;
        RECT 253.240 101.240 253.495 101.815 ;
        RECT 253.665 101.790 253.835 101.980 ;
        RECT 254.115 101.970 254.470 102.340 ;
        RECT 255.560 102.060 256.050 102.260 ;
        RECT 256.240 102.060 256.715 102.270 ;
        RECT 253.665 101.620 254.380 101.790 ;
        RECT 253.665 101.070 253.995 101.450 ;
        RECT 254.210 101.240 254.380 101.620 ;
        RECT 255.565 101.070 256.020 101.835 ;
        RECT 256.495 101.660 256.715 102.060 ;
        RECT 256.960 102.060 257.290 102.270 ;
        RECT 256.960 101.660 257.170 102.060 ;
        RECT 257.460 102.025 257.870 102.330 ;
        RECT 258.100 101.890 258.270 102.465 ;
        RECT 258.000 101.770 258.270 101.890 ;
        RECT 257.425 101.725 258.270 101.770 ;
        RECT 257.425 101.600 258.180 101.725 ;
        RECT 257.425 101.450 257.595 101.600 ;
        RECT 258.440 101.570 258.610 102.770 ;
        RECT 258.870 102.610 259.040 103.450 ;
        RECT 259.210 103.280 260.380 103.450 ;
        RECT 259.210 102.780 259.540 103.280 ;
        RECT 260.050 103.240 260.380 103.280 ;
        RECT 260.570 103.200 260.925 103.620 ;
        RECT 259.710 103.020 259.940 103.110 ;
        RECT 261.095 103.020 261.345 103.450 ;
        RECT 259.710 102.780 261.345 103.020 ;
        RECT 261.515 102.860 261.845 103.620 ;
        RECT 262.015 102.780 262.270 103.450 ;
        RECT 262.060 102.770 262.270 102.780 ;
        RECT 258.870 102.440 261.930 102.610 ;
        RECT 258.785 102.060 259.135 102.270 ;
        RECT 259.305 102.060 259.750 102.260 ;
        RECT 259.920 102.060 260.395 102.260 ;
        RECT 256.295 101.240 257.595 101.450 ;
        RECT 257.850 101.070 258.180 101.430 ;
        RECT 258.350 101.240 258.610 101.570 ;
        RECT 258.870 101.720 259.935 101.890 ;
        RECT 258.870 101.240 259.040 101.720 ;
        RECT 259.210 101.070 259.540 101.550 ;
        RECT 259.765 101.490 259.935 101.720 ;
        RECT 260.115 101.660 260.395 102.060 ;
        RECT 260.665 102.060 260.995 102.260 ;
        RECT 261.165 102.060 261.530 102.260 ;
        RECT 260.665 101.660 260.950 102.060 ;
        RECT 261.760 101.890 261.930 102.440 ;
        RECT 261.130 101.720 261.930 101.890 ;
        RECT 261.130 101.490 261.300 101.720 ;
        RECT 262.100 101.650 262.270 102.770 ;
        RECT 262.465 103.230 262.800 103.450 ;
        RECT 263.805 103.240 264.160 103.620 ;
        RECT 262.465 102.610 262.720 103.230 ;
        RECT 262.970 103.070 263.200 103.110 ;
        RECT 264.330 103.070 264.580 103.450 ;
        RECT 262.970 102.870 264.580 103.070 ;
        RECT 262.970 102.780 263.155 102.870 ;
        RECT 263.745 102.860 264.580 102.870 ;
        RECT 264.830 102.840 265.080 103.620 ;
        RECT 265.250 102.770 265.510 103.450 ;
        RECT 263.310 102.670 263.640 102.700 ;
        RECT 263.310 102.610 265.110 102.670 ;
        RECT 262.465 102.500 265.170 102.610 ;
        RECT 262.465 102.440 263.640 102.500 ;
        RECT 264.970 102.465 265.170 102.500 ;
        RECT 262.460 102.060 262.950 102.260 ;
        RECT 263.140 102.060 263.615 102.270 ;
        RECT 262.085 101.570 262.270 101.650 ;
        RECT 259.765 101.240 261.300 101.490 ;
        RECT 261.470 101.070 261.800 101.550 ;
        RECT 262.015 101.240 262.270 101.570 ;
        RECT 262.465 101.070 262.920 101.835 ;
        RECT 263.395 101.660 263.615 102.060 ;
        RECT 263.860 102.060 264.190 102.270 ;
        RECT 263.860 101.660 264.070 102.060 ;
        RECT 264.360 102.025 264.770 102.330 ;
        RECT 265.000 101.890 265.170 102.465 ;
        RECT 264.900 101.770 265.170 101.890 ;
        RECT 264.325 101.725 265.170 101.770 ;
        RECT 264.325 101.600 265.080 101.725 ;
        RECT 264.325 101.450 264.495 101.600 ;
        RECT 265.340 101.570 265.510 102.770 ;
        RECT 265.685 102.470 265.945 103.620 ;
        RECT 266.120 102.545 266.375 103.450 ;
        RECT 266.545 102.860 266.875 103.620 ;
        RECT 267.090 102.690 267.260 103.450 ;
        RECT 263.195 101.240 264.495 101.450 ;
        RECT 264.750 101.070 265.080 101.430 ;
        RECT 265.250 101.240 265.510 101.570 ;
        RECT 265.685 101.070 265.945 101.910 ;
        RECT 266.120 101.815 266.290 102.545 ;
        RECT 266.545 102.520 267.260 102.690 ;
        RECT 267.520 102.530 268.730 103.620 ;
        RECT 266.545 102.310 266.715 102.520 ;
        RECT 266.460 101.980 266.715 102.310 ;
        RECT 266.120 101.240 266.375 101.815 ;
        RECT 266.545 101.790 266.715 101.980 ;
        RECT 266.995 101.970 267.350 102.340 ;
        RECT 267.520 101.820 268.040 102.360 ;
        RECT 268.210 101.990 268.730 102.530 ;
        RECT 268.905 102.430 269.160 103.310 ;
        RECT 269.330 102.480 269.635 103.620 ;
        RECT 269.975 103.240 270.305 103.620 ;
        RECT 270.485 103.070 270.655 103.360 ;
        RECT 270.825 103.160 271.075 103.620 ;
        RECT 269.855 102.900 270.655 103.070 ;
        RECT 271.245 103.110 272.115 103.450 ;
        RECT 266.545 101.620 267.260 101.790 ;
        RECT 266.545 101.070 266.875 101.450 ;
        RECT 267.090 101.240 267.260 101.620 ;
        RECT 267.520 101.070 268.730 101.820 ;
        RECT 268.905 101.780 269.115 102.430 ;
        RECT 269.855 102.310 270.025 102.900 ;
        RECT 271.245 102.730 271.415 103.110 ;
        RECT 272.350 102.990 272.520 103.450 ;
        RECT 272.690 103.160 273.060 103.620 ;
        RECT 273.355 103.020 273.525 103.360 ;
        RECT 273.695 103.190 274.025 103.620 ;
        RECT 274.260 103.020 274.430 103.360 ;
        RECT 270.195 102.560 271.415 102.730 ;
        RECT 271.585 102.650 272.045 102.940 ;
        RECT 272.350 102.820 272.910 102.990 ;
        RECT 273.355 102.850 274.430 103.020 ;
        RECT 274.600 103.120 275.280 103.450 ;
        RECT 275.495 103.120 275.745 103.450 ;
        RECT 275.915 103.160 276.165 103.620 ;
        RECT 272.740 102.680 272.910 102.820 ;
        RECT 271.585 102.640 272.550 102.650 ;
        RECT 271.245 102.470 271.415 102.560 ;
        RECT 271.875 102.480 272.550 102.640 ;
        RECT 269.285 102.280 270.025 102.310 ;
        RECT 269.285 101.980 270.200 102.280 ;
        RECT 269.875 101.805 270.200 101.980 ;
        RECT 268.905 101.250 269.160 101.780 ;
        RECT 269.330 101.070 269.635 101.530 ;
        RECT 269.880 101.450 270.200 101.805 ;
        RECT 270.370 102.020 270.910 102.390 ;
        RECT 271.245 102.300 271.650 102.470 ;
        RECT 270.370 101.620 270.610 102.020 ;
        RECT 271.090 101.850 271.310 102.130 ;
        RECT 270.780 101.680 271.310 101.850 ;
        RECT 270.780 101.450 270.950 101.680 ;
        RECT 271.480 101.520 271.650 102.300 ;
        RECT 271.820 101.690 272.170 102.310 ;
        RECT 272.340 101.690 272.550 102.480 ;
        RECT 272.740 102.510 274.240 102.680 ;
        RECT 272.740 101.820 272.910 102.510 ;
        RECT 274.600 102.340 274.770 103.120 ;
        RECT 275.575 102.990 275.745 103.120 ;
        RECT 273.080 102.170 274.770 102.340 ;
        RECT 274.940 102.560 275.405 102.950 ;
        RECT 275.575 102.820 275.970 102.990 ;
        RECT 273.080 101.990 273.250 102.170 ;
        RECT 269.880 101.280 270.950 101.450 ;
        RECT 271.120 101.070 271.310 101.510 ;
        RECT 271.480 101.240 272.430 101.520 ;
        RECT 272.740 101.430 273.000 101.820 ;
        RECT 273.420 101.750 274.210 102.000 ;
        RECT 272.650 101.260 273.000 101.430 ;
        RECT 273.210 101.070 273.540 101.530 ;
        RECT 274.415 101.460 274.585 102.170 ;
        RECT 274.940 101.970 275.110 102.560 ;
        RECT 274.755 101.750 275.110 101.970 ;
        RECT 275.280 101.750 275.630 102.370 ;
        RECT 275.800 101.460 275.970 102.820 ;
        RECT 276.335 102.650 276.660 103.435 ;
        RECT 276.140 101.600 276.600 102.650 ;
        RECT 274.415 101.290 275.270 101.460 ;
        RECT 275.475 101.290 275.970 101.460 ;
        RECT 276.140 101.070 276.470 101.430 ;
        RECT 276.830 101.330 277.000 103.450 ;
        RECT 277.170 103.120 277.500 103.620 ;
        RECT 277.670 102.950 277.925 103.450 ;
        RECT 277.175 102.780 277.925 102.950 ;
        RECT 277.175 101.790 277.405 102.780 ;
        RECT 277.575 101.960 277.925 102.610 ;
        RECT 278.100 102.455 278.390 103.620 ;
        RECT 278.560 102.860 279.075 103.270 ;
        RECT 279.310 102.860 279.480 103.620 ;
        RECT 279.650 103.280 281.680 103.450 ;
        RECT 278.560 102.050 278.900 102.860 ;
        RECT 279.650 102.615 279.820 103.280 ;
        RECT 280.215 102.940 281.340 103.110 ;
        RECT 279.070 102.425 279.820 102.615 ;
        RECT 279.990 102.600 281.000 102.770 ;
        RECT 278.560 101.880 279.790 102.050 ;
        RECT 277.175 101.620 277.925 101.790 ;
        RECT 277.170 101.070 277.500 101.450 ;
        RECT 277.670 101.330 277.925 101.620 ;
        RECT 278.100 101.070 278.390 101.795 ;
        RECT 278.835 101.275 279.080 101.880 ;
        RECT 279.300 101.070 279.810 101.605 ;
        RECT 279.990 101.240 280.180 102.600 ;
        RECT 280.350 101.920 280.625 102.400 ;
        RECT 280.350 101.750 280.630 101.920 ;
        RECT 280.830 101.800 281.000 102.600 ;
        RECT 281.170 101.810 281.340 102.940 ;
        RECT 281.510 102.310 281.680 103.280 ;
        RECT 281.850 102.480 282.020 103.620 ;
        RECT 282.190 102.480 282.525 103.450 ;
        RECT 281.510 101.980 281.705 102.310 ;
        RECT 281.930 101.980 282.185 102.310 ;
        RECT 281.930 101.810 282.100 101.980 ;
        RECT 282.355 101.810 282.525 102.480 ;
        RECT 282.705 102.470 282.965 103.620 ;
        RECT 283.140 102.545 283.395 103.450 ;
        RECT 283.565 102.860 283.895 103.620 ;
        RECT 284.110 102.690 284.280 103.450 ;
        RECT 285.005 102.950 285.260 103.450 ;
        RECT 285.430 103.120 285.760 103.620 ;
        RECT 285.005 102.780 285.755 102.950 ;
        RECT 280.350 101.240 280.625 101.750 ;
        RECT 281.170 101.640 282.100 101.810 ;
        RECT 281.170 101.605 281.345 101.640 ;
        RECT 280.815 101.240 281.345 101.605 ;
        RECT 281.770 101.070 282.100 101.470 ;
        RECT 282.270 101.240 282.525 101.810 ;
        RECT 282.705 101.070 282.965 101.910 ;
        RECT 283.140 101.815 283.310 102.545 ;
        RECT 283.565 102.520 284.280 102.690 ;
        RECT 283.565 102.310 283.735 102.520 ;
        RECT 283.480 101.980 283.735 102.310 ;
        RECT 283.140 101.240 283.395 101.815 ;
        RECT 283.565 101.790 283.735 101.980 ;
        RECT 284.015 101.970 284.370 102.340 ;
        RECT 285.005 101.960 285.355 102.610 ;
        RECT 285.525 101.790 285.755 102.780 ;
        RECT 283.565 101.620 284.280 101.790 ;
        RECT 283.565 101.070 283.895 101.450 ;
        RECT 284.110 101.240 284.280 101.620 ;
        RECT 285.005 101.620 285.755 101.790 ;
        RECT 285.005 101.330 285.260 101.620 ;
        RECT 285.430 101.070 285.760 101.450 ;
        RECT 285.930 101.330 286.100 103.450 ;
        RECT 286.270 102.650 286.595 103.435 ;
        RECT 286.765 103.160 287.015 103.620 ;
        RECT 287.185 103.120 287.435 103.450 ;
        RECT 287.650 103.120 288.330 103.450 ;
        RECT 287.185 102.990 287.355 103.120 ;
        RECT 286.960 102.820 287.355 102.990 ;
        RECT 286.330 101.600 286.790 102.650 ;
        RECT 286.960 101.460 287.130 102.820 ;
        RECT 287.525 102.560 287.990 102.950 ;
        RECT 287.300 101.750 287.650 102.370 ;
        RECT 287.820 101.970 287.990 102.560 ;
        RECT 288.160 102.340 288.330 103.120 ;
        RECT 288.500 103.020 288.670 103.360 ;
        RECT 288.905 103.190 289.235 103.620 ;
        RECT 289.405 103.020 289.575 103.360 ;
        RECT 289.870 103.160 290.240 103.620 ;
        RECT 288.500 102.850 289.575 103.020 ;
        RECT 290.410 102.990 290.580 103.450 ;
        RECT 290.815 103.110 291.685 103.450 ;
        RECT 291.855 103.160 292.105 103.620 ;
        RECT 290.020 102.820 290.580 102.990 ;
        RECT 290.020 102.680 290.190 102.820 ;
        RECT 288.690 102.510 290.190 102.680 ;
        RECT 290.885 102.650 291.345 102.940 ;
        RECT 288.160 102.170 289.850 102.340 ;
        RECT 287.820 101.750 288.175 101.970 ;
        RECT 288.345 101.460 288.515 102.170 ;
        RECT 288.720 101.750 289.510 102.000 ;
        RECT 289.680 101.990 289.850 102.170 ;
        RECT 290.020 101.820 290.190 102.510 ;
        RECT 286.460 101.070 286.790 101.430 ;
        RECT 286.960 101.290 287.455 101.460 ;
        RECT 287.660 101.290 288.515 101.460 ;
        RECT 289.390 101.070 289.720 101.530 ;
        RECT 289.930 101.430 290.190 101.820 ;
        RECT 290.380 102.640 291.345 102.650 ;
        RECT 291.515 102.730 291.685 103.110 ;
        RECT 292.275 103.070 292.445 103.360 ;
        RECT 292.625 103.240 292.955 103.620 ;
        RECT 292.275 102.900 293.075 103.070 ;
        RECT 290.380 102.480 291.055 102.640 ;
        RECT 291.515 102.560 292.735 102.730 ;
        RECT 290.380 101.690 290.590 102.480 ;
        RECT 291.515 102.470 291.685 102.560 ;
        RECT 290.760 101.690 291.110 102.310 ;
        RECT 291.280 102.300 291.685 102.470 ;
        RECT 291.280 101.520 291.450 102.300 ;
        RECT 291.620 101.850 291.840 102.130 ;
        RECT 292.020 102.020 292.560 102.390 ;
        RECT 292.905 102.310 293.075 102.900 ;
        RECT 293.295 102.480 293.600 103.620 ;
        RECT 293.770 102.430 294.020 103.310 ;
        RECT 294.190 102.480 294.440 103.620 ;
        RECT 292.905 102.280 293.645 102.310 ;
        RECT 291.620 101.680 292.150 101.850 ;
        RECT 289.930 101.260 290.280 101.430 ;
        RECT 290.500 101.240 291.450 101.520 ;
        RECT 291.620 101.070 291.810 101.510 ;
        RECT 291.980 101.450 292.150 101.680 ;
        RECT 292.320 101.620 292.560 102.020 ;
        RECT 292.730 101.980 293.645 102.280 ;
        RECT 292.730 101.805 293.055 101.980 ;
        RECT 292.730 101.450 293.050 101.805 ;
        RECT 293.815 101.780 294.020 102.430 ;
        RECT 294.665 102.430 294.920 103.310 ;
        RECT 295.090 102.480 295.395 103.620 ;
        RECT 295.735 103.240 296.065 103.620 ;
        RECT 296.245 103.070 296.415 103.360 ;
        RECT 296.585 103.160 296.835 103.620 ;
        RECT 295.615 102.900 296.415 103.070 ;
        RECT 297.005 103.110 297.875 103.450 ;
        RECT 291.980 101.280 293.050 101.450 ;
        RECT 293.295 101.070 293.600 101.530 ;
        RECT 293.770 101.250 294.020 101.780 ;
        RECT 294.190 101.070 294.440 101.825 ;
        RECT 294.665 101.780 294.875 102.430 ;
        RECT 295.615 102.310 295.785 102.900 ;
        RECT 297.005 102.730 297.175 103.110 ;
        RECT 298.110 102.990 298.280 103.450 ;
        RECT 298.450 103.160 298.820 103.620 ;
        RECT 299.115 103.020 299.285 103.360 ;
        RECT 299.455 103.190 299.785 103.620 ;
        RECT 300.020 103.020 300.190 103.360 ;
        RECT 295.955 102.560 297.175 102.730 ;
        RECT 297.345 102.650 297.805 102.940 ;
        RECT 298.110 102.820 298.670 102.990 ;
        RECT 299.115 102.850 300.190 103.020 ;
        RECT 300.360 103.120 301.040 103.450 ;
        RECT 301.255 103.120 301.505 103.450 ;
        RECT 301.675 103.160 301.925 103.620 ;
        RECT 298.500 102.680 298.670 102.820 ;
        RECT 297.345 102.640 298.310 102.650 ;
        RECT 297.005 102.470 297.175 102.560 ;
        RECT 297.635 102.480 298.310 102.640 ;
        RECT 295.045 102.280 295.785 102.310 ;
        RECT 295.045 101.980 295.960 102.280 ;
        RECT 295.635 101.805 295.960 101.980 ;
        RECT 294.665 101.250 294.920 101.780 ;
        RECT 295.090 101.070 295.395 101.530 ;
        RECT 295.640 101.450 295.960 101.805 ;
        RECT 296.130 102.020 296.670 102.390 ;
        RECT 297.005 102.300 297.410 102.470 ;
        RECT 296.130 101.620 296.370 102.020 ;
        RECT 296.850 101.850 297.070 102.130 ;
        RECT 296.540 101.680 297.070 101.850 ;
        RECT 296.540 101.450 296.710 101.680 ;
        RECT 297.240 101.520 297.410 102.300 ;
        RECT 297.580 101.690 297.930 102.310 ;
        RECT 298.100 101.690 298.310 102.480 ;
        RECT 298.500 102.510 300.000 102.680 ;
        RECT 298.500 101.820 298.670 102.510 ;
        RECT 300.360 102.340 300.530 103.120 ;
        RECT 301.335 102.990 301.505 103.120 ;
        RECT 298.840 102.170 300.530 102.340 ;
        RECT 300.700 102.560 301.165 102.950 ;
        RECT 301.335 102.820 301.730 102.990 ;
        RECT 298.840 101.990 299.010 102.170 ;
        RECT 295.640 101.280 296.710 101.450 ;
        RECT 296.880 101.070 297.070 101.510 ;
        RECT 297.240 101.240 298.190 101.520 ;
        RECT 298.500 101.430 298.760 101.820 ;
        RECT 299.180 101.750 299.970 102.000 ;
        RECT 298.410 101.260 298.760 101.430 ;
        RECT 298.970 101.070 299.300 101.530 ;
        RECT 300.175 101.460 300.345 102.170 ;
        RECT 300.700 101.970 300.870 102.560 ;
        RECT 300.515 101.750 300.870 101.970 ;
        RECT 301.040 101.750 301.390 102.370 ;
        RECT 301.560 101.460 301.730 102.820 ;
        RECT 302.095 102.650 302.420 103.435 ;
        RECT 301.900 101.600 302.360 102.650 ;
        RECT 300.175 101.290 301.030 101.460 ;
        RECT 301.235 101.290 301.730 101.460 ;
        RECT 301.900 101.070 302.230 101.430 ;
        RECT 302.590 101.330 302.760 103.450 ;
        RECT 302.930 103.120 303.260 103.620 ;
        RECT 303.430 102.950 303.685 103.450 ;
        RECT 302.935 102.780 303.685 102.950 ;
        RECT 302.935 101.790 303.165 102.780 ;
        RECT 303.335 101.960 303.685 102.610 ;
        RECT 303.860 102.455 304.150 103.620 ;
        RECT 304.410 102.690 304.580 103.450 ;
        RECT 304.795 102.860 305.125 103.620 ;
        RECT 304.410 102.520 305.125 102.690 ;
        RECT 305.295 102.545 305.550 103.450 ;
        RECT 304.320 101.970 304.675 102.340 ;
        RECT 304.955 102.310 305.125 102.520 ;
        RECT 304.955 101.980 305.210 102.310 ;
        RECT 302.935 101.620 303.685 101.790 ;
        RECT 302.930 101.070 303.260 101.450 ;
        RECT 303.430 101.330 303.685 101.620 ;
        RECT 303.860 101.070 304.150 101.795 ;
        RECT 304.955 101.790 305.125 101.980 ;
        RECT 305.380 101.815 305.550 102.545 ;
        RECT 305.725 102.470 305.985 103.620 ;
        RECT 307.080 102.650 307.390 103.450 ;
        RECT 307.560 102.820 307.870 103.620 ;
        RECT 308.040 102.990 308.300 103.450 ;
        RECT 308.470 103.160 308.725 103.620 ;
        RECT 308.900 102.990 309.160 103.450 ;
        RECT 308.040 102.820 309.160 102.990 ;
        RECT 307.080 102.480 308.110 102.650 ;
        RECT 304.410 101.620 305.125 101.790 ;
        RECT 304.410 101.240 304.580 101.620 ;
        RECT 304.795 101.070 305.125 101.450 ;
        RECT 305.295 101.240 305.550 101.815 ;
        RECT 305.725 101.070 305.985 101.910 ;
        RECT 307.080 101.570 307.250 102.480 ;
        RECT 307.420 101.740 307.770 102.310 ;
        RECT 307.940 102.230 308.110 102.480 ;
        RECT 308.900 102.570 309.160 102.820 ;
        RECT 309.330 102.750 309.615 103.620 ;
        RECT 308.900 102.400 309.655 102.570 ;
        RECT 307.940 102.060 309.080 102.230 ;
        RECT 309.250 101.890 309.655 102.400 ;
        RECT 309.840 102.530 311.050 103.620 ;
        RECT 309.840 101.990 310.360 102.530 ;
        RECT 308.005 101.720 309.655 101.890 ;
        RECT 310.530 101.820 311.050 102.360 ;
        RECT 307.080 101.240 307.380 101.570 ;
        RECT 307.550 101.070 307.825 101.550 ;
        RECT 308.005 101.330 308.300 101.720 ;
        RECT 308.470 101.070 308.725 101.550 ;
        RECT 308.900 101.330 309.160 101.720 ;
        RECT 309.330 101.070 309.610 101.550 ;
        RECT 309.840 101.070 311.050 101.820 ;
        RECT 162.095 100.900 311.135 101.070 ;
        RECT 162.180 100.150 163.390 100.900 ;
        RECT 162.180 99.610 162.700 100.150 ;
        RECT 163.560 100.130 165.230 100.900 ;
        RECT 165.490 100.350 165.660 100.730 ;
        RECT 165.840 100.520 166.170 100.900 ;
        RECT 165.490 100.180 166.155 100.350 ;
        RECT 166.350 100.225 166.610 100.730 ;
        RECT 162.870 99.440 163.390 99.980 ;
        RECT 163.560 99.610 164.310 100.130 ;
        RECT 164.480 99.440 165.230 99.960 ;
        RECT 165.420 99.630 165.750 100.000 ;
        RECT 165.985 99.925 166.155 100.180 ;
        RECT 165.985 99.595 166.270 99.925 ;
        RECT 165.985 99.450 166.155 99.595 ;
        RECT 162.180 98.350 163.390 99.440 ;
        RECT 163.560 98.350 165.230 99.440 ;
        RECT 165.490 99.280 166.155 99.450 ;
        RECT 166.440 99.425 166.610 100.225 ;
        RECT 166.785 100.060 167.045 100.900 ;
        RECT 167.220 100.155 167.475 100.730 ;
        RECT 167.645 100.520 167.975 100.900 ;
        RECT 168.190 100.350 168.360 100.730 ;
        RECT 167.645 100.180 168.360 100.350 ;
        RECT 168.625 100.350 168.880 100.640 ;
        RECT 169.050 100.520 169.380 100.900 ;
        RECT 168.625 100.180 169.375 100.350 ;
        RECT 165.490 98.520 165.660 99.280 ;
        RECT 165.840 98.350 166.170 99.110 ;
        RECT 166.340 98.520 166.610 99.425 ;
        RECT 166.785 98.350 167.045 99.500 ;
        RECT 167.220 99.425 167.390 100.155 ;
        RECT 167.645 99.990 167.815 100.180 ;
        RECT 167.560 99.660 167.815 99.990 ;
        RECT 167.645 99.450 167.815 99.660 ;
        RECT 168.095 99.630 168.450 100.000 ;
        RECT 167.220 98.520 167.475 99.425 ;
        RECT 167.645 99.280 168.360 99.450 ;
        RECT 168.625 99.360 168.975 100.010 ;
        RECT 167.645 98.350 167.975 99.110 ;
        RECT 168.190 98.520 168.360 99.280 ;
        RECT 169.145 99.190 169.375 100.180 ;
        RECT 168.625 99.020 169.375 99.190 ;
        RECT 168.625 98.520 168.880 99.020 ;
        RECT 169.050 98.350 169.380 98.850 ;
        RECT 169.550 98.520 169.720 100.640 ;
        RECT 170.080 100.540 170.410 100.900 ;
        RECT 170.580 100.510 171.075 100.680 ;
        RECT 171.280 100.510 172.135 100.680 ;
        RECT 169.950 99.320 170.410 100.370 ;
        RECT 169.890 98.535 170.215 99.320 ;
        RECT 170.580 99.150 170.750 100.510 ;
        RECT 170.920 99.600 171.270 100.220 ;
        RECT 171.440 100.000 171.795 100.220 ;
        RECT 171.440 99.410 171.610 100.000 ;
        RECT 171.965 99.800 172.135 100.510 ;
        RECT 173.010 100.440 173.340 100.900 ;
        RECT 173.550 100.540 173.900 100.710 ;
        RECT 172.340 99.970 173.130 100.220 ;
        RECT 173.550 100.150 173.810 100.540 ;
        RECT 174.120 100.450 175.070 100.730 ;
        RECT 175.240 100.460 175.430 100.900 ;
        RECT 175.600 100.520 176.670 100.690 ;
        RECT 173.300 99.800 173.470 99.980 ;
        RECT 170.580 98.980 170.975 99.150 ;
        RECT 171.145 99.020 171.610 99.410 ;
        RECT 171.780 99.630 173.470 99.800 ;
        RECT 170.805 98.850 170.975 98.980 ;
        RECT 171.780 98.850 171.950 99.630 ;
        RECT 173.640 99.460 173.810 100.150 ;
        RECT 172.310 99.290 173.810 99.460 ;
        RECT 174.000 99.490 174.210 100.280 ;
        RECT 174.380 99.660 174.730 100.280 ;
        RECT 174.900 99.670 175.070 100.450 ;
        RECT 175.600 100.290 175.770 100.520 ;
        RECT 175.240 100.120 175.770 100.290 ;
        RECT 175.240 99.840 175.460 100.120 ;
        RECT 175.940 99.950 176.180 100.350 ;
        RECT 174.900 99.500 175.305 99.670 ;
        RECT 175.640 99.580 176.180 99.950 ;
        RECT 176.350 100.165 176.670 100.520 ;
        RECT 176.915 100.440 177.220 100.900 ;
        RECT 177.390 100.190 177.645 100.720 ;
        RECT 176.350 99.990 176.675 100.165 ;
        RECT 176.350 99.690 177.265 99.990 ;
        RECT 176.525 99.660 177.265 99.690 ;
        RECT 174.000 99.330 174.675 99.490 ;
        RECT 175.135 99.410 175.305 99.500 ;
        RECT 174.000 99.320 174.965 99.330 ;
        RECT 173.640 99.150 173.810 99.290 ;
        RECT 170.385 98.350 170.635 98.810 ;
        RECT 170.805 98.520 171.055 98.850 ;
        RECT 171.270 98.520 171.950 98.850 ;
        RECT 172.120 98.950 173.195 99.120 ;
        RECT 173.640 98.980 174.200 99.150 ;
        RECT 174.505 99.030 174.965 99.320 ;
        RECT 175.135 99.240 176.355 99.410 ;
        RECT 172.120 98.610 172.290 98.950 ;
        RECT 172.525 98.350 172.855 98.780 ;
        RECT 173.025 98.610 173.195 98.950 ;
        RECT 173.490 98.350 173.860 98.810 ;
        RECT 174.030 98.520 174.200 98.980 ;
        RECT 175.135 98.860 175.305 99.240 ;
        RECT 176.525 99.070 176.695 99.660 ;
        RECT 177.435 99.540 177.645 100.190 ;
        RECT 174.435 98.520 175.305 98.860 ;
        RECT 175.895 98.900 176.695 99.070 ;
        RECT 175.475 98.350 175.725 98.810 ;
        RECT 175.895 98.610 176.065 98.900 ;
        RECT 176.245 98.350 176.575 98.730 ;
        RECT 176.915 98.350 177.220 99.490 ;
        RECT 177.390 98.660 177.645 99.540 ;
        RECT 177.825 100.160 178.080 100.730 ;
        RECT 178.250 100.500 178.580 100.900 ;
        RECT 179.005 100.365 179.535 100.730 ;
        RECT 179.005 100.330 179.180 100.365 ;
        RECT 178.250 100.160 179.180 100.330 ;
        RECT 179.725 100.220 180.000 100.730 ;
        RECT 177.825 99.490 177.995 100.160 ;
        RECT 178.250 99.990 178.420 100.160 ;
        RECT 178.165 99.660 178.420 99.990 ;
        RECT 178.645 99.660 178.840 99.990 ;
        RECT 177.825 98.520 178.160 99.490 ;
        RECT 178.330 98.350 178.500 99.490 ;
        RECT 178.670 98.690 178.840 99.660 ;
        RECT 179.010 99.030 179.180 100.160 ;
        RECT 179.350 99.370 179.520 100.170 ;
        RECT 179.720 100.050 180.000 100.220 ;
        RECT 179.725 99.570 180.000 100.050 ;
        RECT 180.170 99.370 180.360 100.730 ;
        RECT 180.540 100.365 181.050 100.900 ;
        RECT 181.270 100.090 181.515 100.695 ;
        RECT 182.050 100.350 182.220 100.730 ;
        RECT 182.400 100.520 182.730 100.900 ;
        RECT 182.050 100.180 182.715 100.350 ;
        RECT 182.910 100.225 183.170 100.730 ;
        RECT 180.560 99.920 181.790 100.090 ;
        RECT 179.350 99.200 180.360 99.370 ;
        RECT 180.530 99.355 181.280 99.545 ;
        RECT 179.010 98.860 180.135 99.030 ;
        RECT 180.530 98.690 180.700 99.355 ;
        RECT 181.450 99.110 181.790 99.920 ;
        RECT 181.980 99.630 182.310 100.000 ;
        RECT 182.545 99.925 182.715 100.180 ;
        RECT 182.545 99.595 182.830 99.925 ;
        RECT 182.545 99.450 182.715 99.595 ;
        RECT 178.670 98.520 180.700 98.690 ;
        RECT 180.870 98.350 181.040 99.110 ;
        RECT 181.275 98.700 181.790 99.110 ;
        RECT 182.050 99.280 182.715 99.450 ;
        RECT 183.000 99.425 183.170 100.225 ;
        RECT 182.050 98.520 182.220 99.280 ;
        RECT 182.400 98.350 182.730 99.110 ;
        RECT 182.900 98.520 183.170 99.425 ;
        RECT 183.805 100.160 184.060 100.730 ;
        RECT 184.230 100.500 184.560 100.900 ;
        RECT 184.985 100.365 185.515 100.730 ;
        RECT 184.985 100.330 185.160 100.365 ;
        RECT 184.230 100.160 185.160 100.330 ;
        RECT 185.705 100.220 185.980 100.730 ;
        RECT 183.805 99.490 183.975 100.160 ;
        RECT 184.230 99.990 184.400 100.160 ;
        RECT 184.145 99.660 184.400 99.990 ;
        RECT 184.625 99.660 184.820 99.990 ;
        RECT 183.805 98.520 184.140 99.490 ;
        RECT 184.310 98.350 184.480 99.490 ;
        RECT 184.650 98.690 184.820 99.660 ;
        RECT 184.990 99.030 185.160 100.160 ;
        RECT 185.330 99.370 185.500 100.170 ;
        RECT 185.700 100.050 185.980 100.220 ;
        RECT 185.705 99.570 185.980 100.050 ;
        RECT 186.150 99.370 186.340 100.730 ;
        RECT 186.520 100.365 187.030 100.900 ;
        RECT 187.250 100.090 187.495 100.695 ;
        RECT 187.940 100.175 188.230 100.900 ;
        RECT 188.405 100.350 188.660 100.640 ;
        RECT 188.830 100.520 189.160 100.900 ;
        RECT 188.405 100.180 189.155 100.350 ;
        RECT 186.540 99.920 187.770 100.090 ;
        RECT 185.330 99.200 186.340 99.370 ;
        RECT 186.510 99.355 187.260 99.545 ;
        RECT 184.990 98.860 186.115 99.030 ;
        RECT 186.510 98.690 186.680 99.355 ;
        RECT 187.430 99.110 187.770 99.920 ;
        RECT 184.650 98.520 186.680 98.690 ;
        RECT 186.850 98.350 187.020 99.110 ;
        RECT 187.255 98.700 187.770 99.110 ;
        RECT 187.940 98.350 188.230 99.515 ;
        RECT 188.405 99.360 188.755 100.010 ;
        RECT 188.925 99.190 189.155 100.180 ;
        RECT 188.405 99.020 189.155 99.190 ;
        RECT 188.405 98.520 188.660 99.020 ;
        RECT 188.830 98.350 189.160 98.850 ;
        RECT 189.330 98.520 189.500 100.640 ;
        RECT 189.860 100.540 190.190 100.900 ;
        RECT 190.360 100.510 190.855 100.680 ;
        RECT 191.060 100.510 191.915 100.680 ;
        RECT 189.730 99.320 190.190 100.370 ;
        RECT 189.670 98.535 189.995 99.320 ;
        RECT 190.360 99.150 190.530 100.510 ;
        RECT 190.700 99.600 191.050 100.220 ;
        RECT 191.220 100.000 191.575 100.220 ;
        RECT 191.220 99.410 191.390 100.000 ;
        RECT 191.745 99.800 191.915 100.510 ;
        RECT 192.790 100.440 193.120 100.900 ;
        RECT 193.330 100.540 193.680 100.710 ;
        RECT 192.120 99.970 192.910 100.220 ;
        RECT 193.330 100.150 193.590 100.540 ;
        RECT 193.900 100.450 194.850 100.730 ;
        RECT 195.020 100.460 195.210 100.900 ;
        RECT 195.380 100.520 196.450 100.690 ;
        RECT 193.080 99.800 193.250 99.980 ;
        RECT 190.360 98.980 190.755 99.150 ;
        RECT 190.925 99.020 191.390 99.410 ;
        RECT 191.560 99.630 193.250 99.800 ;
        RECT 190.585 98.850 190.755 98.980 ;
        RECT 191.560 98.850 191.730 99.630 ;
        RECT 193.420 99.460 193.590 100.150 ;
        RECT 192.090 99.290 193.590 99.460 ;
        RECT 193.780 99.490 193.990 100.280 ;
        RECT 194.160 99.660 194.510 100.280 ;
        RECT 194.680 99.670 194.850 100.450 ;
        RECT 195.380 100.290 195.550 100.520 ;
        RECT 195.020 100.120 195.550 100.290 ;
        RECT 195.020 99.840 195.240 100.120 ;
        RECT 195.720 99.950 195.960 100.350 ;
        RECT 194.680 99.500 195.085 99.670 ;
        RECT 195.420 99.580 195.960 99.950 ;
        RECT 196.130 100.165 196.450 100.520 ;
        RECT 196.695 100.440 197.000 100.900 ;
        RECT 197.170 100.190 197.425 100.720 ;
        RECT 196.130 99.990 196.455 100.165 ;
        RECT 196.130 99.690 197.045 99.990 ;
        RECT 196.305 99.660 197.045 99.690 ;
        RECT 193.780 99.330 194.455 99.490 ;
        RECT 194.915 99.410 195.085 99.500 ;
        RECT 193.780 99.320 194.745 99.330 ;
        RECT 193.420 99.150 193.590 99.290 ;
        RECT 190.165 98.350 190.415 98.810 ;
        RECT 190.585 98.520 190.835 98.850 ;
        RECT 191.050 98.520 191.730 98.850 ;
        RECT 191.900 98.950 192.975 99.120 ;
        RECT 193.420 98.980 193.980 99.150 ;
        RECT 194.285 99.030 194.745 99.320 ;
        RECT 194.915 99.240 196.135 99.410 ;
        RECT 191.900 98.610 192.070 98.950 ;
        RECT 192.305 98.350 192.635 98.780 ;
        RECT 192.805 98.610 192.975 98.950 ;
        RECT 193.270 98.350 193.640 98.810 ;
        RECT 193.810 98.520 193.980 98.980 ;
        RECT 194.915 98.860 195.085 99.240 ;
        RECT 196.305 99.070 196.475 99.660 ;
        RECT 197.215 99.540 197.425 100.190 ;
        RECT 197.875 100.090 198.120 100.695 ;
        RECT 198.340 100.365 198.850 100.900 ;
        RECT 194.215 98.520 195.085 98.860 ;
        RECT 195.675 98.900 196.475 99.070 ;
        RECT 195.255 98.350 195.505 98.810 ;
        RECT 195.675 98.610 195.845 98.900 ;
        RECT 196.025 98.350 196.355 98.730 ;
        RECT 196.695 98.350 197.000 99.490 ;
        RECT 197.170 98.660 197.425 99.540 ;
        RECT 197.600 99.920 198.830 100.090 ;
        RECT 197.600 99.110 197.940 99.920 ;
        RECT 198.110 99.355 198.860 99.545 ;
        RECT 197.600 98.700 198.115 99.110 ;
        RECT 198.350 98.350 198.520 99.110 ;
        RECT 198.690 98.690 198.860 99.355 ;
        RECT 199.030 99.370 199.220 100.730 ;
        RECT 199.390 100.560 199.665 100.730 ;
        RECT 199.390 100.390 199.670 100.560 ;
        RECT 199.390 99.570 199.665 100.390 ;
        RECT 199.855 100.365 200.385 100.730 ;
        RECT 200.810 100.500 201.140 100.900 ;
        RECT 200.210 100.330 200.385 100.365 ;
        RECT 199.870 99.370 200.040 100.170 ;
        RECT 199.030 99.200 200.040 99.370 ;
        RECT 200.210 100.160 201.140 100.330 ;
        RECT 201.310 100.160 201.565 100.730 ;
        RECT 200.210 99.030 200.380 100.160 ;
        RECT 200.970 99.990 201.140 100.160 ;
        RECT 199.255 98.860 200.380 99.030 ;
        RECT 200.550 99.660 200.745 99.990 ;
        RECT 200.970 99.660 201.225 99.990 ;
        RECT 200.550 98.690 200.720 99.660 ;
        RECT 201.395 99.490 201.565 100.160 ;
        RECT 198.690 98.520 200.720 98.690 ;
        RECT 200.890 98.350 201.060 99.490 ;
        RECT 201.230 98.520 201.565 99.490 ;
        RECT 201.745 100.190 202.000 100.720 ;
        RECT 202.170 100.440 202.475 100.900 ;
        RECT 202.720 100.520 203.790 100.690 ;
        RECT 201.745 99.540 201.955 100.190 ;
        RECT 202.720 100.165 203.040 100.520 ;
        RECT 202.715 99.990 203.040 100.165 ;
        RECT 202.125 99.690 203.040 99.990 ;
        RECT 203.210 99.950 203.450 100.350 ;
        RECT 203.620 100.290 203.790 100.520 ;
        RECT 203.960 100.460 204.150 100.900 ;
        RECT 204.320 100.450 205.270 100.730 ;
        RECT 205.490 100.540 205.840 100.710 ;
        RECT 203.620 100.120 204.150 100.290 ;
        RECT 202.125 99.660 202.865 99.690 ;
        RECT 201.745 98.660 202.000 99.540 ;
        RECT 202.170 98.350 202.475 99.490 ;
        RECT 202.695 99.070 202.865 99.660 ;
        RECT 203.210 99.580 203.750 99.950 ;
        RECT 203.930 99.840 204.150 100.120 ;
        RECT 204.320 99.670 204.490 100.450 ;
        RECT 204.085 99.500 204.490 99.670 ;
        RECT 204.660 99.660 205.010 100.280 ;
        RECT 204.085 99.410 204.255 99.500 ;
        RECT 205.180 99.490 205.390 100.280 ;
        RECT 203.035 99.240 204.255 99.410 ;
        RECT 204.715 99.330 205.390 99.490 ;
        RECT 202.695 98.900 203.495 99.070 ;
        RECT 202.815 98.350 203.145 98.730 ;
        RECT 203.325 98.610 203.495 98.900 ;
        RECT 204.085 98.860 204.255 99.240 ;
        RECT 204.425 99.320 205.390 99.330 ;
        RECT 205.580 100.150 205.840 100.540 ;
        RECT 206.050 100.440 206.380 100.900 ;
        RECT 207.255 100.510 208.110 100.680 ;
        RECT 208.315 100.510 208.810 100.680 ;
        RECT 208.980 100.540 209.310 100.900 ;
        RECT 205.580 99.460 205.750 100.150 ;
        RECT 205.920 99.800 206.090 99.980 ;
        RECT 206.260 99.970 207.050 100.220 ;
        RECT 207.255 99.800 207.425 100.510 ;
        RECT 207.595 100.000 207.950 100.220 ;
        RECT 205.920 99.630 207.610 99.800 ;
        RECT 204.425 99.030 204.885 99.320 ;
        RECT 205.580 99.290 207.080 99.460 ;
        RECT 205.580 99.150 205.750 99.290 ;
        RECT 205.190 98.980 205.750 99.150 ;
        RECT 203.665 98.350 203.915 98.810 ;
        RECT 204.085 98.520 204.955 98.860 ;
        RECT 205.190 98.520 205.360 98.980 ;
        RECT 206.195 98.950 207.270 99.120 ;
        RECT 205.530 98.350 205.900 98.810 ;
        RECT 206.195 98.610 206.365 98.950 ;
        RECT 206.535 98.350 206.865 98.780 ;
        RECT 207.100 98.610 207.270 98.950 ;
        RECT 207.440 98.850 207.610 99.630 ;
        RECT 207.780 99.410 207.950 100.000 ;
        RECT 208.120 99.600 208.470 100.220 ;
        RECT 207.780 99.020 208.245 99.410 ;
        RECT 208.640 99.150 208.810 100.510 ;
        RECT 208.980 99.320 209.440 100.370 ;
        RECT 208.415 98.980 208.810 99.150 ;
        RECT 208.415 98.850 208.585 98.980 ;
        RECT 207.440 98.520 208.120 98.850 ;
        RECT 208.335 98.520 208.585 98.850 ;
        RECT 208.755 98.350 209.005 98.810 ;
        RECT 209.175 98.535 209.500 99.320 ;
        RECT 209.670 98.520 209.840 100.640 ;
        RECT 210.010 100.520 210.340 100.900 ;
        RECT 210.510 100.350 210.765 100.640 ;
        RECT 210.015 100.180 210.765 100.350 ;
        RECT 210.940 100.225 211.200 100.730 ;
        RECT 211.380 100.520 211.710 100.900 ;
        RECT 211.890 100.350 212.060 100.730 ;
        RECT 210.015 99.190 210.245 100.180 ;
        RECT 210.415 99.360 210.765 100.010 ;
        RECT 210.940 99.425 211.110 100.225 ;
        RECT 211.395 100.180 212.060 100.350 ;
        RECT 211.395 99.925 211.565 100.180 ;
        RECT 212.320 100.150 213.530 100.900 ;
        RECT 213.700 100.175 213.990 100.900 ;
        RECT 215.170 100.350 215.340 100.730 ;
        RECT 215.555 100.520 215.885 100.900 ;
        RECT 215.170 100.180 215.885 100.350 ;
        RECT 211.280 99.595 211.565 99.925 ;
        RECT 211.800 99.630 212.130 100.000 ;
        RECT 212.320 99.610 212.840 100.150 ;
        RECT 211.395 99.450 211.565 99.595 ;
        RECT 210.015 99.020 210.765 99.190 ;
        RECT 210.010 98.350 210.340 98.850 ;
        RECT 210.510 98.520 210.765 99.020 ;
        RECT 210.940 98.520 211.210 99.425 ;
        RECT 211.395 99.280 212.060 99.450 ;
        RECT 213.010 99.440 213.530 99.980 ;
        RECT 215.080 99.630 215.435 100.000 ;
        RECT 215.715 99.990 215.885 100.180 ;
        RECT 216.055 100.155 216.310 100.730 ;
        RECT 215.715 99.660 215.970 99.990 ;
        RECT 211.380 98.350 211.710 99.110 ;
        RECT 211.890 98.520 212.060 99.280 ;
        RECT 212.320 98.350 213.530 99.440 ;
        RECT 213.700 98.350 213.990 99.515 ;
        RECT 215.715 99.450 215.885 99.660 ;
        RECT 215.170 99.280 215.885 99.450 ;
        RECT 216.140 99.425 216.310 100.155 ;
        RECT 216.485 100.060 216.745 100.900 ;
        RECT 217.010 100.350 217.180 100.730 ;
        RECT 217.395 100.520 217.725 100.900 ;
        RECT 217.010 100.180 217.725 100.350 ;
        RECT 216.920 99.630 217.275 100.000 ;
        RECT 217.555 99.990 217.725 100.180 ;
        RECT 217.895 100.155 218.150 100.730 ;
        RECT 217.555 99.660 217.810 99.990 ;
        RECT 215.170 98.520 215.340 99.280 ;
        RECT 215.555 98.350 215.885 99.110 ;
        RECT 216.055 98.520 216.310 99.425 ;
        RECT 216.485 98.350 216.745 99.500 ;
        RECT 217.555 99.450 217.725 99.660 ;
        RECT 217.010 99.280 217.725 99.450 ;
        RECT 217.980 99.425 218.150 100.155 ;
        RECT 218.325 100.060 218.585 100.900 ;
        RECT 217.010 98.520 217.180 99.280 ;
        RECT 217.395 98.350 217.725 99.110 ;
        RECT 217.895 98.520 218.150 99.425 ;
        RECT 218.325 98.350 218.585 99.500 ;
        RECT 219.680 98.520 220.430 100.730 ;
        RECT 221.525 100.160 221.780 100.730 ;
        RECT 221.950 100.500 222.280 100.900 ;
        RECT 222.705 100.365 223.235 100.730 ;
        RECT 222.705 100.330 222.880 100.365 ;
        RECT 221.950 100.160 222.880 100.330 ;
        RECT 221.525 99.490 221.695 100.160 ;
        RECT 221.950 99.990 222.120 100.160 ;
        RECT 221.865 99.660 222.120 99.990 ;
        RECT 222.345 99.660 222.540 99.990 ;
        RECT 221.525 98.520 221.860 99.490 ;
        RECT 222.030 98.350 222.200 99.490 ;
        RECT 222.370 98.690 222.540 99.660 ;
        RECT 222.710 99.030 222.880 100.160 ;
        RECT 223.050 99.370 223.220 100.170 ;
        RECT 223.425 99.880 223.700 100.730 ;
        RECT 223.420 99.710 223.700 99.880 ;
        RECT 223.425 99.570 223.700 99.710 ;
        RECT 223.870 99.370 224.060 100.730 ;
        RECT 224.240 100.365 224.750 100.900 ;
        RECT 224.970 100.090 225.215 100.695 ;
        RECT 225.660 100.130 228.250 100.900 ;
        RECT 228.420 100.225 228.680 100.730 ;
        RECT 228.860 100.520 229.190 100.900 ;
        RECT 229.370 100.350 229.540 100.730 ;
        RECT 224.260 99.920 225.490 100.090 ;
        RECT 223.050 99.200 224.060 99.370 ;
        RECT 224.230 99.355 224.980 99.545 ;
        RECT 222.710 98.860 223.835 99.030 ;
        RECT 224.230 98.690 224.400 99.355 ;
        RECT 225.150 99.110 225.490 99.920 ;
        RECT 225.660 99.610 226.870 100.130 ;
        RECT 227.040 99.440 228.250 99.960 ;
        RECT 222.370 98.520 224.400 98.690 ;
        RECT 224.570 98.350 224.740 99.110 ;
        RECT 224.975 98.700 225.490 99.110 ;
        RECT 225.660 98.350 228.250 99.440 ;
        RECT 228.420 99.425 228.590 100.225 ;
        RECT 228.875 100.180 229.540 100.350 ;
        RECT 228.875 99.925 229.045 100.180 ;
        RECT 229.805 100.160 230.060 100.730 ;
        RECT 230.230 100.500 230.560 100.900 ;
        RECT 230.985 100.365 231.515 100.730 ;
        RECT 230.985 100.330 231.160 100.365 ;
        RECT 230.230 100.160 231.160 100.330 ;
        RECT 228.760 99.595 229.045 99.925 ;
        RECT 229.280 99.630 229.610 100.000 ;
        RECT 228.875 99.450 229.045 99.595 ;
        RECT 229.805 99.490 229.975 100.160 ;
        RECT 230.230 99.990 230.400 100.160 ;
        RECT 230.145 99.660 230.400 99.990 ;
        RECT 230.625 99.660 230.820 99.990 ;
        RECT 228.420 98.520 228.690 99.425 ;
        RECT 228.875 99.280 229.540 99.450 ;
        RECT 228.860 98.350 229.190 99.110 ;
        RECT 229.370 98.520 229.540 99.280 ;
        RECT 229.805 98.520 230.140 99.490 ;
        RECT 230.310 98.350 230.480 99.490 ;
        RECT 230.650 98.690 230.820 99.660 ;
        RECT 230.990 99.030 231.160 100.160 ;
        RECT 231.330 99.370 231.500 100.170 ;
        RECT 231.705 99.880 231.980 100.730 ;
        RECT 231.700 99.710 231.980 99.880 ;
        RECT 231.705 99.570 231.980 99.710 ;
        RECT 232.150 99.370 232.340 100.730 ;
        RECT 232.520 100.365 233.030 100.900 ;
        RECT 233.250 100.090 233.495 100.695 ;
        RECT 233.940 100.355 239.285 100.900 ;
        RECT 232.540 99.920 233.770 100.090 ;
        RECT 231.330 99.200 232.340 99.370 ;
        RECT 232.510 99.355 233.260 99.545 ;
        RECT 230.990 98.860 232.115 99.030 ;
        RECT 232.510 98.690 232.680 99.355 ;
        RECT 233.430 99.110 233.770 99.920 ;
        RECT 235.525 99.525 235.865 100.355 ;
        RECT 239.460 100.175 239.750 100.900 ;
        RECT 239.920 100.225 240.180 100.730 ;
        RECT 240.360 100.520 240.690 100.900 ;
        RECT 240.870 100.350 241.040 100.730 ;
        RECT 230.650 98.520 232.680 98.690 ;
        RECT 232.850 98.350 233.020 99.110 ;
        RECT 233.255 98.700 233.770 99.110 ;
        RECT 237.345 98.785 237.695 100.035 ;
        RECT 233.940 98.350 239.285 98.785 ;
        RECT 239.460 98.350 239.750 99.515 ;
        RECT 239.920 99.425 240.090 100.225 ;
        RECT 240.375 100.180 241.040 100.350 ;
        RECT 240.375 99.925 240.545 100.180 ;
        RECT 241.300 100.130 242.970 100.900 ;
        RECT 243.605 100.190 243.860 100.720 ;
        RECT 244.030 100.440 244.335 100.900 ;
        RECT 244.580 100.520 245.650 100.690 ;
        RECT 240.260 99.595 240.545 99.925 ;
        RECT 240.780 99.630 241.110 100.000 ;
        RECT 241.300 99.610 242.050 100.130 ;
        RECT 240.375 99.450 240.545 99.595 ;
        RECT 239.920 98.520 240.190 99.425 ;
        RECT 240.375 99.280 241.040 99.450 ;
        RECT 242.220 99.440 242.970 99.960 ;
        RECT 240.360 98.350 240.690 99.110 ;
        RECT 240.870 98.520 241.040 99.280 ;
        RECT 241.300 98.350 242.970 99.440 ;
        RECT 243.605 99.540 243.815 100.190 ;
        RECT 244.580 100.165 244.900 100.520 ;
        RECT 244.575 99.990 244.900 100.165 ;
        RECT 243.985 99.690 244.900 99.990 ;
        RECT 245.070 99.950 245.310 100.350 ;
        RECT 245.480 100.290 245.650 100.520 ;
        RECT 245.820 100.460 246.010 100.900 ;
        RECT 246.180 100.450 247.130 100.730 ;
        RECT 247.350 100.540 247.700 100.710 ;
        RECT 245.480 100.120 246.010 100.290 ;
        RECT 243.985 99.660 244.725 99.690 ;
        RECT 243.605 98.660 243.860 99.540 ;
        RECT 244.030 98.350 244.335 99.490 ;
        RECT 244.555 99.070 244.725 99.660 ;
        RECT 245.070 99.580 245.610 99.950 ;
        RECT 245.790 99.840 246.010 100.120 ;
        RECT 246.180 99.670 246.350 100.450 ;
        RECT 245.945 99.500 246.350 99.670 ;
        RECT 246.520 99.660 246.870 100.280 ;
        RECT 245.945 99.410 246.115 99.500 ;
        RECT 247.040 99.490 247.250 100.280 ;
        RECT 244.895 99.240 246.115 99.410 ;
        RECT 246.575 99.330 247.250 99.490 ;
        RECT 244.555 98.900 245.355 99.070 ;
        RECT 244.675 98.350 245.005 98.730 ;
        RECT 245.185 98.610 245.355 98.900 ;
        RECT 245.945 98.860 246.115 99.240 ;
        RECT 246.285 99.320 247.250 99.330 ;
        RECT 247.440 100.150 247.700 100.540 ;
        RECT 247.910 100.440 248.240 100.900 ;
        RECT 249.115 100.510 249.970 100.680 ;
        RECT 250.175 100.510 250.670 100.680 ;
        RECT 250.840 100.540 251.170 100.900 ;
        RECT 247.440 99.460 247.610 100.150 ;
        RECT 247.780 99.800 247.950 99.980 ;
        RECT 248.120 99.970 248.910 100.220 ;
        RECT 249.115 99.800 249.285 100.510 ;
        RECT 249.455 100.000 249.810 100.220 ;
        RECT 247.780 99.630 249.470 99.800 ;
        RECT 246.285 99.030 246.745 99.320 ;
        RECT 247.440 99.290 248.940 99.460 ;
        RECT 247.440 99.150 247.610 99.290 ;
        RECT 247.050 98.980 247.610 99.150 ;
        RECT 245.525 98.350 245.775 98.810 ;
        RECT 245.945 98.520 246.815 98.860 ;
        RECT 247.050 98.520 247.220 98.980 ;
        RECT 248.055 98.950 249.130 99.120 ;
        RECT 247.390 98.350 247.760 98.810 ;
        RECT 248.055 98.610 248.225 98.950 ;
        RECT 248.395 98.350 248.725 98.780 ;
        RECT 248.960 98.610 249.130 98.950 ;
        RECT 249.300 98.850 249.470 99.630 ;
        RECT 249.640 99.410 249.810 100.000 ;
        RECT 249.980 99.600 250.330 100.220 ;
        RECT 249.640 99.020 250.105 99.410 ;
        RECT 250.500 99.150 250.670 100.510 ;
        RECT 250.840 99.320 251.300 100.370 ;
        RECT 250.275 98.980 250.670 99.150 ;
        RECT 250.275 98.850 250.445 98.980 ;
        RECT 249.300 98.520 249.980 98.850 ;
        RECT 250.195 98.520 250.445 98.850 ;
        RECT 250.615 98.350 250.865 98.810 ;
        RECT 251.035 98.535 251.360 99.320 ;
        RECT 251.530 98.520 251.700 100.640 ;
        RECT 251.870 100.520 252.200 100.900 ;
        RECT 252.370 100.350 252.625 100.640 ;
        RECT 251.875 100.180 252.625 100.350 ;
        RECT 251.875 99.190 252.105 100.180 ;
        RECT 253.725 100.135 254.180 100.900 ;
        RECT 254.455 100.520 255.755 100.730 ;
        RECT 256.010 100.540 256.340 100.900 ;
        RECT 255.585 100.370 255.755 100.520 ;
        RECT 256.510 100.400 256.770 100.730 ;
        RECT 256.540 100.390 256.770 100.400 ;
        RECT 252.275 99.360 252.625 100.010 ;
        RECT 254.655 99.910 254.875 100.310 ;
        RECT 253.720 99.710 254.210 99.910 ;
        RECT 254.400 99.700 254.875 99.910 ;
        RECT 255.120 99.910 255.330 100.310 ;
        RECT 255.585 100.245 256.340 100.370 ;
        RECT 255.585 100.200 256.430 100.245 ;
        RECT 256.160 100.080 256.430 100.200 ;
        RECT 255.120 99.700 255.450 99.910 ;
        RECT 255.620 99.640 256.030 99.945 ;
        RECT 253.725 99.470 254.900 99.530 ;
        RECT 256.260 99.505 256.430 100.080 ;
        RECT 256.230 99.470 256.430 99.505 ;
        RECT 253.725 99.360 256.430 99.470 ;
        RECT 251.875 99.020 252.625 99.190 ;
        RECT 251.870 98.350 252.200 98.850 ;
        RECT 252.370 98.520 252.625 99.020 ;
        RECT 253.725 98.740 253.980 99.360 ;
        RECT 254.570 99.300 256.370 99.360 ;
        RECT 254.570 99.270 254.900 99.300 ;
        RECT 256.600 99.200 256.770 100.390 ;
        RECT 256.940 100.130 258.610 100.900 ;
        RECT 258.870 100.250 259.040 100.730 ;
        RECT 259.210 100.420 259.540 100.900 ;
        RECT 259.765 100.480 261.300 100.730 ;
        RECT 259.765 100.250 259.935 100.480 ;
        RECT 256.940 99.610 257.690 100.130 ;
        RECT 258.870 100.080 259.935 100.250 ;
        RECT 257.860 99.440 258.610 99.960 ;
        RECT 260.115 99.910 260.395 100.310 ;
        RECT 258.785 99.700 259.135 99.910 ;
        RECT 259.305 99.710 259.750 99.910 ;
        RECT 259.920 99.710 260.395 99.910 ;
        RECT 260.665 99.910 260.950 100.310 ;
        RECT 261.130 100.250 261.300 100.480 ;
        RECT 261.470 100.420 261.800 100.900 ;
        RECT 262.015 100.400 262.270 100.730 ;
        RECT 262.085 100.320 262.270 100.400 ;
        RECT 261.130 100.080 261.930 100.250 ;
        RECT 260.665 99.710 260.995 99.910 ;
        RECT 261.165 99.880 261.530 99.910 ;
        RECT 261.165 99.710 261.540 99.880 ;
        RECT 261.760 99.530 261.930 100.080 ;
        RECT 254.230 99.100 254.415 99.190 ;
        RECT 255.005 99.100 255.840 99.110 ;
        RECT 254.230 98.900 255.840 99.100 ;
        RECT 254.230 98.860 254.460 98.900 ;
        RECT 253.725 98.520 254.060 98.740 ;
        RECT 255.065 98.350 255.420 98.730 ;
        RECT 255.590 98.520 255.840 98.900 ;
        RECT 256.090 98.350 256.340 99.130 ;
        RECT 256.510 98.520 256.770 99.200 ;
        RECT 256.940 98.350 258.610 99.440 ;
        RECT 258.870 99.360 261.930 99.530 ;
        RECT 258.870 98.520 259.040 99.360 ;
        RECT 262.100 99.190 262.270 100.320 ;
        RECT 263.120 100.270 263.450 100.630 ;
        RECT 264.070 100.440 264.320 100.900 ;
        RECT 264.490 100.440 265.050 100.730 ;
        RECT 263.120 100.080 264.510 100.270 ;
        RECT 264.340 99.990 264.510 100.080 ;
        RECT 262.935 99.660 263.610 99.910 ;
        RECT 263.830 99.660 264.170 99.910 ;
        RECT 264.340 99.660 264.630 99.990 ;
        RECT 262.935 99.300 263.200 99.660 ;
        RECT 264.340 99.410 264.510 99.660 ;
        RECT 259.210 98.690 259.540 99.190 ;
        RECT 259.710 98.950 261.345 99.190 ;
        RECT 259.710 98.860 259.940 98.950 ;
        RECT 260.050 98.690 260.380 98.730 ;
        RECT 259.210 98.520 260.380 98.690 ;
        RECT 260.570 98.350 260.925 98.770 ;
        RECT 261.095 98.520 261.345 98.950 ;
        RECT 261.515 98.350 261.845 99.110 ;
        RECT 262.015 98.520 262.270 99.190 ;
        RECT 263.570 99.240 264.510 99.410 ;
        RECT 263.120 98.350 263.400 99.020 ;
        RECT 263.570 98.690 263.870 99.240 ;
        RECT 264.800 99.070 265.050 100.440 ;
        RECT 265.220 100.175 265.510 100.900 ;
        RECT 265.680 100.355 271.025 100.900 ;
        RECT 267.265 99.525 267.605 100.355 ;
        RECT 271.205 100.350 271.460 100.640 ;
        RECT 271.630 100.520 271.960 100.900 ;
        RECT 271.205 100.180 271.955 100.350 ;
        RECT 264.070 98.350 264.400 99.070 ;
        RECT 264.590 98.520 265.050 99.070 ;
        RECT 265.220 98.350 265.510 99.515 ;
        RECT 269.085 98.785 269.435 100.035 ;
        RECT 271.205 99.360 271.555 100.010 ;
        RECT 271.725 99.190 271.955 100.180 ;
        RECT 271.205 99.020 271.955 99.190 ;
        RECT 265.680 98.350 271.025 98.785 ;
        RECT 271.205 98.520 271.460 99.020 ;
        RECT 271.630 98.350 271.960 98.850 ;
        RECT 272.130 98.520 272.300 100.640 ;
        RECT 272.660 100.540 272.990 100.900 ;
        RECT 273.160 100.510 273.655 100.680 ;
        RECT 273.860 100.510 274.715 100.680 ;
        RECT 272.530 99.320 272.990 100.370 ;
        RECT 272.470 98.535 272.795 99.320 ;
        RECT 273.160 99.150 273.330 100.510 ;
        RECT 273.500 99.600 273.850 100.220 ;
        RECT 274.020 100.000 274.375 100.220 ;
        RECT 274.020 99.410 274.190 100.000 ;
        RECT 274.545 99.800 274.715 100.510 ;
        RECT 275.590 100.440 275.920 100.900 ;
        RECT 276.130 100.540 276.480 100.710 ;
        RECT 274.920 99.970 275.710 100.220 ;
        RECT 276.130 100.150 276.390 100.540 ;
        RECT 276.700 100.450 277.650 100.730 ;
        RECT 277.820 100.460 278.010 100.900 ;
        RECT 278.180 100.520 279.250 100.690 ;
        RECT 275.880 99.800 276.050 99.980 ;
        RECT 273.160 98.980 273.555 99.150 ;
        RECT 273.725 99.020 274.190 99.410 ;
        RECT 274.360 99.630 276.050 99.800 ;
        RECT 273.385 98.850 273.555 98.980 ;
        RECT 274.360 98.850 274.530 99.630 ;
        RECT 276.220 99.460 276.390 100.150 ;
        RECT 274.890 99.290 276.390 99.460 ;
        RECT 276.580 99.490 276.790 100.280 ;
        RECT 276.960 99.660 277.310 100.280 ;
        RECT 277.480 99.670 277.650 100.450 ;
        RECT 278.180 100.290 278.350 100.520 ;
        RECT 277.820 100.120 278.350 100.290 ;
        RECT 277.820 99.840 278.040 100.120 ;
        RECT 278.520 99.950 278.760 100.350 ;
        RECT 277.480 99.500 277.885 99.670 ;
        RECT 278.220 99.580 278.760 99.950 ;
        RECT 278.930 100.165 279.250 100.520 ;
        RECT 279.495 100.440 279.800 100.900 ;
        RECT 279.970 100.190 280.225 100.720 ;
        RECT 278.930 99.990 279.255 100.165 ;
        RECT 278.930 99.690 279.845 99.990 ;
        RECT 279.105 99.660 279.845 99.690 ;
        RECT 276.580 99.330 277.255 99.490 ;
        RECT 277.715 99.410 277.885 99.500 ;
        RECT 276.580 99.320 277.545 99.330 ;
        RECT 276.220 99.150 276.390 99.290 ;
        RECT 272.965 98.350 273.215 98.810 ;
        RECT 273.385 98.520 273.635 98.850 ;
        RECT 273.850 98.520 274.530 98.850 ;
        RECT 274.700 98.950 275.775 99.120 ;
        RECT 276.220 98.980 276.780 99.150 ;
        RECT 277.085 99.030 277.545 99.320 ;
        RECT 277.715 99.240 278.935 99.410 ;
        RECT 274.700 98.610 274.870 98.950 ;
        RECT 275.105 98.350 275.435 98.780 ;
        RECT 275.605 98.610 275.775 98.950 ;
        RECT 276.070 98.350 276.440 98.810 ;
        RECT 276.610 98.520 276.780 98.980 ;
        RECT 277.715 98.860 277.885 99.240 ;
        RECT 279.105 99.070 279.275 99.660 ;
        RECT 280.015 99.540 280.225 100.190 ;
        RECT 280.490 100.350 280.660 100.730 ;
        RECT 280.840 100.520 281.170 100.900 ;
        RECT 280.490 100.180 281.155 100.350 ;
        RECT 281.350 100.225 281.610 100.730 ;
        RECT 280.420 99.630 280.750 100.000 ;
        RECT 280.985 99.925 281.155 100.180 ;
        RECT 277.015 98.520 277.885 98.860 ;
        RECT 278.475 98.900 279.275 99.070 ;
        RECT 278.055 98.350 278.305 98.810 ;
        RECT 278.475 98.610 278.645 98.900 ;
        RECT 278.825 98.350 279.155 98.730 ;
        RECT 279.495 98.350 279.800 99.490 ;
        RECT 279.970 98.660 280.225 99.540 ;
        RECT 280.985 99.595 281.270 99.925 ;
        RECT 280.985 99.450 281.155 99.595 ;
        RECT 280.490 99.280 281.155 99.450 ;
        RECT 281.440 99.425 281.610 100.225 ;
        RECT 281.785 100.350 282.040 100.640 ;
        RECT 282.210 100.520 282.540 100.900 ;
        RECT 281.785 100.180 282.535 100.350 ;
        RECT 280.490 98.520 280.660 99.280 ;
        RECT 280.840 98.350 281.170 99.110 ;
        RECT 281.340 98.520 281.610 99.425 ;
        RECT 281.785 99.360 282.135 100.010 ;
        RECT 282.305 99.190 282.535 100.180 ;
        RECT 281.785 99.020 282.535 99.190 ;
        RECT 281.785 98.520 282.040 99.020 ;
        RECT 282.210 98.350 282.540 98.850 ;
        RECT 282.710 98.520 282.880 100.640 ;
        RECT 283.240 100.540 283.570 100.900 ;
        RECT 283.740 100.510 284.235 100.680 ;
        RECT 284.440 100.510 285.295 100.680 ;
        RECT 283.110 99.320 283.570 100.370 ;
        RECT 283.050 98.535 283.375 99.320 ;
        RECT 283.740 99.150 283.910 100.510 ;
        RECT 284.080 99.600 284.430 100.220 ;
        RECT 284.600 100.000 284.955 100.220 ;
        RECT 284.600 99.410 284.770 100.000 ;
        RECT 285.125 99.800 285.295 100.510 ;
        RECT 286.170 100.440 286.500 100.900 ;
        RECT 286.710 100.540 287.060 100.710 ;
        RECT 285.500 99.970 286.290 100.220 ;
        RECT 286.710 100.150 286.970 100.540 ;
        RECT 287.280 100.450 288.230 100.730 ;
        RECT 288.400 100.460 288.590 100.900 ;
        RECT 288.760 100.520 289.830 100.690 ;
        RECT 286.460 99.800 286.630 99.980 ;
        RECT 283.740 98.980 284.135 99.150 ;
        RECT 284.305 99.020 284.770 99.410 ;
        RECT 284.940 99.630 286.630 99.800 ;
        RECT 283.965 98.850 284.135 98.980 ;
        RECT 284.940 98.850 285.110 99.630 ;
        RECT 286.800 99.460 286.970 100.150 ;
        RECT 285.470 99.290 286.970 99.460 ;
        RECT 287.160 99.490 287.370 100.280 ;
        RECT 287.540 99.660 287.890 100.280 ;
        RECT 288.060 99.670 288.230 100.450 ;
        RECT 288.760 100.290 288.930 100.520 ;
        RECT 288.400 100.120 288.930 100.290 ;
        RECT 288.400 99.840 288.620 100.120 ;
        RECT 289.100 99.950 289.340 100.350 ;
        RECT 288.060 99.500 288.465 99.670 ;
        RECT 288.800 99.580 289.340 99.950 ;
        RECT 289.510 100.165 289.830 100.520 ;
        RECT 290.075 100.440 290.380 100.900 ;
        RECT 290.550 100.190 290.805 100.720 ;
        RECT 289.510 99.990 289.835 100.165 ;
        RECT 289.510 99.690 290.425 99.990 ;
        RECT 289.685 99.660 290.425 99.690 ;
        RECT 287.160 99.330 287.835 99.490 ;
        RECT 288.295 99.410 288.465 99.500 ;
        RECT 287.160 99.320 288.125 99.330 ;
        RECT 286.800 99.150 286.970 99.290 ;
        RECT 283.545 98.350 283.795 98.810 ;
        RECT 283.965 98.520 284.215 98.850 ;
        RECT 284.430 98.520 285.110 98.850 ;
        RECT 285.280 98.950 286.355 99.120 ;
        RECT 286.800 98.980 287.360 99.150 ;
        RECT 287.665 99.030 288.125 99.320 ;
        RECT 288.295 99.240 289.515 99.410 ;
        RECT 285.280 98.610 285.450 98.950 ;
        RECT 285.685 98.350 286.015 98.780 ;
        RECT 286.185 98.610 286.355 98.950 ;
        RECT 286.650 98.350 287.020 98.810 ;
        RECT 287.190 98.520 287.360 98.980 ;
        RECT 288.295 98.860 288.465 99.240 ;
        RECT 289.685 99.070 289.855 99.660 ;
        RECT 290.595 99.540 290.805 100.190 ;
        RECT 290.980 100.175 291.270 100.900 ;
        RECT 292.365 100.350 292.620 100.640 ;
        RECT 292.790 100.520 293.120 100.900 ;
        RECT 292.365 100.180 293.115 100.350 ;
        RECT 287.595 98.520 288.465 98.860 ;
        RECT 289.055 98.900 289.855 99.070 ;
        RECT 288.635 98.350 288.885 98.810 ;
        RECT 289.055 98.610 289.225 98.900 ;
        RECT 289.405 98.350 289.735 98.730 ;
        RECT 290.075 98.350 290.380 99.490 ;
        RECT 290.550 98.660 290.805 99.540 ;
        RECT 290.980 98.350 291.270 99.515 ;
        RECT 292.365 99.360 292.715 100.010 ;
        RECT 292.885 99.190 293.115 100.180 ;
        RECT 292.365 99.020 293.115 99.190 ;
        RECT 292.365 98.520 292.620 99.020 ;
        RECT 292.790 98.350 293.120 98.850 ;
        RECT 293.290 98.520 293.460 100.640 ;
        RECT 293.820 100.540 294.150 100.900 ;
        RECT 294.320 100.510 294.815 100.680 ;
        RECT 295.020 100.510 295.875 100.680 ;
        RECT 293.690 99.320 294.150 100.370 ;
        RECT 293.630 98.535 293.955 99.320 ;
        RECT 294.320 99.150 294.490 100.510 ;
        RECT 294.660 99.600 295.010 100.220 ;
        RECT 295.180 100.000 295.535 100.220 ;
        RECT 295.180 99.410 295.350 100.000 ;
        RECT 295.705 99.800 295.875 100.510 ;
        RECT 296.750 100.440 297.080 100.900 ;
        RECT 297.290 100.540 297.640 100.710 ;
        RECT 296.080 99.970 296.870 100.220 ;
        RECT 297.290 100.150 297.550 100.540 ;
        RECT 297.860 100.450 298.810 100.730 ;
        RECT 298.980 100.460 299.170 100.900 ;
        RECT 299.340 100.520 300.410 100.690 ;
        RECT 297.040 99.800 297.210 99.980 ;
        RECT 294.320 98.980 294.715 99.150 ;
        RECT 294.885 99.020 295.350 99.410 ;
        RECT 295.520 99.630 297.210 99.800 ;
        RECT 294.545 98.850 294.715 98.980 ;
        RECT 295.520 98.850 295.690 99.630 ;
        RECT 297.380 99.460 297.550 100.150 ;
        RECT 296.050 99.290 297.550 99.460 ;
        RECT 297.740 99.490 297.950 100.280 ;
        RECT 298.120 99.660 298.470 100.280 ;
        RECT 298.640 99.670 298.810 100.450 ;
        RECT 299.340 100.290 299.510 100.520 ;
        RECT 298.980 100.120 299.510 100.290 ;
        RECT 298.980 99.840 299.200 100.120 ;
        RECT 299.680 99.950 299.920 100.350 ;
        RECT 298.640 99.500 299.045 99.670 ;
        RECT 299.380 99.580 299.920 99.950 ;
        RECT 300.090 100.165 300.410 100.520 ;
        RECT 300.655 100.440 300.960 100.900 ;
        RECT 301.130 100.190 301.380 100.720 ;
        RECT 300.090 99.990 300.415 100.165 ;
        RECT 300.090 99.690 301.005 99.990 ;
        RECT 300.265 99.660 301.005 99.690 ;
        RECT 297.740 99.330 298.415 99.490 ;
        RECT 298.875 99.410 299.045 99.500 ;
        RECT 297.740 99.320 298.705 99.330 ;
        RECT 297.380 99.150 297.550 99.290 ;
        RECT 294.125 98.350 294.375 98.810 ;
        RECT 294.545 98.520 294.795 98.850 ;
        RECT 295.010 98.520 295.690 98.850 ;
        RECT 295.860 98.950 296.935 99.120 ;
        RECT 297.380 98.980 297.940 99.150 ;
        RECT 298.245 99.030 298.705 99.320 ;
        RECT 298.875 99.240 300.095 99.410 ;
        RECT 295.860 98.610 296.030 98.950 ;
        RECT 296.265 98.350 296.595 98.780 ;
        RECT 296.765 98.610 296.935 98.950 ;
        RECT 297.230 98.350 297.600 98.810 ;
        RECT 297.770 98.520 297.940 98.980 ;
        RECT 298.875 98.860 299.045 99.240 ;
        RECT 300.265 99.070 300.435 99.660 ;
        RECT 301.175 99.540 301.380 100.190 ;
        RECT 301.550 100.145 301.800 100.900 ;
        RECT 302.025 100.160 302.280 100.730 ;
        RECT 302.450 100.500 302.780 100.900 ;
        RECT 303.205 100.365 303.735 100.730 ;
        RECT 303.925 100.560 304.200 100.730 ;
        RECT 303.920 100.390 304.200 100.560 ;
        RECT 303.205 100.330 303.380 100.365 ;
        RECT 302.450 100.160 303.380 100.330 ;
        RECT 298.175 98.520 299.045 98.860 ;
        RECT 299.635 98.900 300.435 99.070 ;
        RECT 299.215 98.350 299.465 98.810 ;
        RECT 299.635 98.610 299.805 98.900 ;
        RECT 299.985 98.350 300.315 98.730 ;
        RECT 300.655 98.350 300.960 99.490 ;
        RECT 301.130 98.660 301.380 99.540 ;
        RECT 302.025 99.490 302.195 100.160 ;
        RECT 302.450 99.990 302.620 100.160 ;
        RECT 302.365 99.660 302.620 99.990 ;
        RECT 302.845 99.660 303.040 99.990 ;
        RECT 301.550 98.350 301.800 99.490 ;
        RECT 302.025 98.520 302.360 99.490 ;
        RECT 302.530 98.350 302.700 99.490 ;
        RECT 302.870 98.690 303.040 99.660 ;
        RECT 303.210 99.030 303.380 100.160 ;
        RECT 303.550 99.370 303.720 100.170 ;
        RECT 303.925 99.570 304.200 100.390 ;
        RECT 304.370 99.370 304.560 100.730 ;
        RECT 304.740 100.365 305.250 100.900 ;
        RECT 305.470 100.090 305.715 100.695 ;
        RECT 306.250 100.350 306.420 100.730 ;
        RECT 306.635 100.520 306.965 100.900 ;
        RECT 306.250 100.180 306.965 100.350 ;
        RECT 304.760 99.920 305.990 100.090 ;
        RECT 303.550 99.200 304.560 99.370 ;
        RECT 304.730 99.355 305.480 99.545 ;
        RECT 303.210 98.860 304.335 99.030 ;
        RECT 304.730 98.690 304.900 99.355 ;
        RECT 305.650 99.110 305.990 99.920 ;
        RECT 306.160 99.630 306.515 100.000 ;
        RECT 306.795 99.990 306.965 100.180 ;
        RECT 307.135 100.155 307.390 100.730 ;
        RECT 306.795 99.660 307.050 99.990 ;
        RECT 306.795 99.450 306.965 99.660 ;
        RECT 302.870 98.520 304.900 98.690 ;
        RECT 305.070 98.350 305.240 99.110 ;
        RECT 305.475 98.700 305.990 99.110 ;
        RECT 306.250 99.280 306.965 99.450 ;
        RECT 307.220 99.425 307.390 100.155 ;
        RECT 307.565 100.060 307.825 100.900 ;
        RECT 308.090 100.350 308.260 100.730 ;
        RECT 308.475 100.520 308.805 100.900 ;
        RECT 308.090 100.180 308.805 100.350 ;
        RECT 308.000 99.630 308.355 100.000 ;
        RECT 308.635 99.990 308.805 100.180 ;
        RECT 308.975 100.155 309.230 100.730 ;
        RECT 308.635 99.660 308.890 99.990 ;
        RECT 306.250 98.520 306.420 99.280 ;
        RECT 306.635 98.350 306.965 99.110 ;
        RECT 307.135 98.520 307.390 99.425 ;
        RECT 307.565 98.350 307.825 99.500 ;
        RECT 308.635 99.450 308.805 99.660 ;
        RECT 308.090 99.280 308.805 99.450 ;
        RECT 309.060 99.425 309.230 100.155 ;
        RECT 309.405 100.060 309.665 100.900 ;
        RECT 309.840 100.150 311.050 100.900 ;
        RECT 308.090 98.520 308.260 99.280 ;
        RECT 308.475 98.350 308.805 99.110 ;
        RECT 308.975 98.520 309.230 99.425 ;
        RECT 309.405 98.350 309.665 99.500 ;
        RECT 309.840 99.440 310.360 99.980 ;
        RECT 310.530 99.610 311.050 100.150 ;
        RECT 309.840 98.350 311.050 99.440 ;
        RECT 162.095 98.180 311.135 98.350 ;
        RECT 162.180 97.090 163.390 98.180 ;
        RECT 163.560 97.745 168.905 98.180 ;
        RECT 162.180 96.380 162.700 96.920 ;
        RECT 162.870 96.550 163.390 97.090 ;
        RECT 162.180 95.630 163.390 96.380 ;
        RECT 165.145 96.175 165.485 97.005 ;
        RECT 166.965 96.495 167.315 97.745 ;
        RECT 170.000 97.105 170.270 98.010 ;
        RECT 170.440 97.420 170.770 98.180 ;
        RECT 170.950 97.250 171.120 98.010 ;
        RECT 170.000 96.305 170.170 97.105 ;
        RECT 170.455 97.080 171.120 97.250 ;
        RECT 171.380 97.105 171.650 98.010 ;
        RECT 171.820 97.420 172.150 98.180 ;
        RECT 172.330 97.250 172.500 98.010 ;
        RECT 170.455 96.935 170.625 97.080 ;
        RECT 170.340 96.605 170.625 96.935 ;
        RECT 170.455 96.350 170.625 96.605 ;
        RECT 170.860 96.530 171.190 96.900 ;
        RECT 163.560 95.630 168.905 96.175 ;
        RECT 170.000 95.800 170.260 96.305 ;
        RECT 170.455 96.180 171.120 96.350 ;
        RECT 170.440 95.630 170.770 96.010 ;
        RECT 170.950 95.800 171.120 96.180 ;
        RECT 171.380 96.305 171.550 97.105 ;
        RECT 171.835 97.080 172.500 97.250 ;
        RECT 172.760 97.105 173.030 98.010 ;
        RECT 173.200 97.420 173.530 98.180 ;
        RECT 173.710 97.250 173.880 98.010 ;
        RECT 171.835 96.935 172.005 97.080 ;
        RECT 171.720 96.605 172.005 96.935 ;
        RECT 171.835 96.350 172.005 96.605 ;
        RECT 172.240 96.530 172.570 96.900 ;
        RECT 171.380 95.800 171.640 96.305 ;
        RECT 171.835 96.180 172.500 96.350 ;
        RECT 171.820 95.630 172.150 96.010 ;
        RECT 172.330 95.800 172.500 96.180 ;
        RECT 172.760 96.305 172.930 97.105 ;
        RECT 173.215 97.080 173.880 97.250 ;
        RECT 173.215 96.935 173.385 97.080 ;
        RECT 175.060 97.015 175.350 98.180 ;
        RECT 175.525 97.040 175.860 98.010 ;
        RECT 176.030 97.040 176.200 98.180 ;
        RECT 176.370 97.840 178.400 98.010 ;
        RECT 173.100 96.605 173.385 96.935 ;
        RECT 173.215 96.350 173.385 96.605 ;
        RECT 173.620 96.530 173.950 96.900 ;
        RECT 175.525 96.370 175.695 97.040 ;
        RECT 176.370 96.870 176.540 97.840 ;
        RECT 175.865 96.540 176.120 96.870 ;
        RECT 176.345 96.540 176.540 96.870 ;
        RECT 176.710 97.500 177.835 97.670 ;
        RECT 175.950 96.370 176.120 96.540 ;
        RECT 176.710 96.370 176.880 97.500 ;
        RECT 172.760 95.800 173.020 96.305 ;
        RECT 173.215 96.180 173.880 96.350 ;
        RECT 173.200 95.630 173.530 96.010 ;
        RECT 173.710 95.800 173.880 96.180 ;
        RECT 175.060 95.630 175.350 96.355 ;
        RECT 175.525 95.800 175.780 96.370 ;
        RECT 175.950 96.200 176.880 96.370 ;
        RECT 177.050 97.160 178.060 97.330 ;
        RECT 177.050 96.360 177.220 97.160 ;
        RECT 177.425 96.820 177.700 96.960 ;
        RECT 177.420 96.650 177.700 96.820 ;
        RECT 176.705 96.165 176.880 96.200 ;
        RECT 175.950 95.630 176.280 96.030 ;
        RECT 176.705 95.800 177.235 96.165 ;
        RECT 177.425 95.800 177.700 96.650 ;
        RECT 177.870 95.800 178.060 97.160 ;
        RECT 178.230 97.175 178.400 97.840 ;
        RECT 178.570 97.420 178.740 98.180 ;
        RECT 178.975 97.420 179.490 97.830 ;
        RECT 178.230 96.985 178.980 97.175 ;
        RECT 179.150 96.610 179.490 97.420 ;
        RECT 179.660 97.090 183.170 98.180 ;
        RECT 183.345 97.510 183.600 98.010 ;
        RECT 183.770 97.680 184.100 98.180 ;
        RECT 183.345 97.340 184.095 97.510 ;
        RECT 178.260 96.440 179.490 96.610 ;
        RECT 178.240 95.630 178.750 96.165 ;
        RECT 178.970 95.835 179.215 96.440 ;
        RECT 179.660 96.400 181.310 96.920 ;
        RECT 181.480 96.570 183.170 97.090 ;
        RECT 183.345 96.520 183.695 97.170 ;
        RECT 179.660 95.630 183.170 96.400 ;
        RECT 183.865 96.350 184.095 97.340 ;
        RECT 183.345 96.180 184.095 96.350 ;
        RECT 183.345 95.890 183.600 96.180 ;
        RECT 183.770 95.630 184.100 96.010 ;
        RECT 184.270 95.890 184.440 98.010 ;
        RECT 184.610 97.210 184.935 97.995 ;
        RECT 185.105 97.720 185.355 98.180 ;
        RECT 185.525 97.680 185.775 98.010 ;
        RECT 185.990 97.680 186.670 98.010 ;
        RECT 185.525 97.550 185.695 97.680 ;
        RECT 185.300 97.380 185.695 97.550 ;
        RECT 184.670 96.160 185.130 97.210 ;
        RECT 185.300 96.020 185.470 97.380 ;
        RECT 185.865 97.120 186.330 97.510 ;
        RECT 185.640 96.310 185.990 96.930 ;
        RECT 186.160 96.530 186.330 97.120 ;
        RECT 186.500 96.900 186.670 97.680 ;
        RECT 186.840 97.580 187.010 97.920 ;
        RECT 187.245 97.750 187.575 98.180 ;
        RECT 187.745 97.580 187.915 97.920 ;
        RECT 188.210 97.720 188.580 98.180 ;
        RECT 186.840 97.410 187.915 97.580 ;
        RECT 188.750 97.550 188.920 98.010 ;
        RECT 189.155 97.670 190.025 98.010 ;
        RECT 190.195 97.720 190.445 98.180 ;
        RECT 188.360 97.380 188.920 97.550 ;
        RECT 188.360 97.240 188.530 97.380 ;
        RECT 187.030 97.070 188.530 97.240 ;
        RECT 189.225 97.210 189.685 97.500 ;
        RECT 186.500 96.730 188.190 96.900 ;
        RECT 186.160 96.310 186.515 96.530 ;
        RECT 186.685 96.020 186.855 96.730 ;
        RECT 187.060 96.310 187.850 96.560 ;
        RECT 188.020 96.550 188.190 96.730 ;
        RECT 188.360 96.380 188.530 97.070 ;
        RECT 184.800 95.630 185.130 95.990 ;
        RECT 185.300 95.850 185.795 96.020 ;
        RECT 186.000 95.850 186.855 96.020 ;
        RECT 187.730 95.630 188.060 96.090 ;
        RECT 188.270 95.990 188.530 96.380 ;
        RECT 188.720 97.200 189.685 97.210 ;
        RECT 189.855 97.290 190.025 97.670 ;
        RECT 190.615 97.630 190.785 97.920 ;
        RECT 190.965 97.800 191.295 98.180 ;
        RECT 190.615 97.460 191.415 97.630 ;
        RECT 188.720 97.040 189.395 97.200 ;
        RECT 189.855 97.120 191.075 97.290 ;
        RECT 188.720 96.250 188.930 97.040 ;
        RECT 189.855 97.030 190.025 97.120 ;
        RECT 189.100 96.250 189.450 96.870 ;
        RECT 189.620 96.860 190.025 97.030 ;
        RECT 189.620 96.080 189.790 96.860 ;
        RECT 189.960 96.410 190.180 96.690 ;
        RECT 190.360 96.580 190.900 96.950 ;
        RECT 191.245 96.870 191.415 97.460 ;
        RECT 191.635 97.040 191.940 98.180 ;
        RECT 192.110 96.990 192.360 97.870 ;
        RECT 192.530 97.040 192.780 98.180 ;
        RECT 193.000 97.105 193.270 98.010 ;
        RECT 193.440 97.420 193.770 98.180 ;
        RECT 193.950 97.250 194.120 98.010 ;
        RECT 191.245 96.840 191.985 96.870 ;
        RECT 189.960 96.240 190.490 96.410 ;
        RECT 188.270 95.820 188.620 95.990 ;
        RECT 188.840 95.800 189.790 96.080 ;
        RECT 189.960 95.630 190.150 96.070 ;
        RECT 190.320 96.010 190.490 96.240 ;
        RECT 190.660 96.180 190.900 96.580 ;
        RECT 191.070 96.540 191.985 96.840 ;
        RECT 191.070 96.365 191.395 96.540 ;
        RECT 191.070 96.010 191.390 96.365 ;
        RECT 192.155 96.340 192.360 96.990 ;
        RECT 190.320 95.840 191.390 96.010 ;
        RECT 191.635 95.630 191.940 96.090 ;
        RECT 192.110 95.810 192.360 96.340 ;
        RECT 192.530 95.630 192.780 96.385 ;
        RECT 193.000 96.305 193.170 97.105 ;
        RECT 193.455 97.080 194.120 97.250 ;
        RECT 194.380 97.090 195.590 98.180 ;
        RECT 193.455 96.935 193.625 97.080 ;
        RECT 193.340 96.605 193.625 96.935 ;
        RECT 193.455 96.350 193.625 96.605 ;
        RECT 193.860 96.530 194.190 96.900 ;
        RECT 194.380 96.380 194.900 96.920 ;
        RECT 195.070 96.550 195.590 97.090 ;
        RECT 195.765 97.040 196.100 98.010 ;
        RECT 196.270 97.040 196.440 98.180 ;
        RECT 196.610 97.840 198.640 98.010 ;
        RECT 193.000 95.800 193.260 96.305 ;
        RECT 193.455 96.180 194.120 96.350 ;
        RECT 193.440 95.630 193.770 96.010 ;
        RECT 193.950 95.800 194.120 96.180 ;
        RECT 194.380 95.630 195.590 96.380 ;
        RECT 195.765 96.370 195.935 97.040 ;
        RECT 196.610 96.870 196.780 97.840 ;
        RECT 196.105 96.540 196.360 96.870 ;
        RECT 196.585 96.540 196.780 96.870 ;
        RECT 196.950 97.500 198.075 97.670 ;
        RECT 196.190 96.370 196.360 96.540 ;
        RECT 196.950 96.370 197.120 97.500 ;
        RECT 195.765 95.800 196.020 96.370 ;
        RECT 196.190 96.200 197.120 96.370 ;
        RECT 197.290 97.160 198.300 97.330 ;
        RECT 197.290 96.360 197.460 97.160 ;
        RECT 197.665 96.480 197.940 96.960 ;
        RECT 197.660 96.310 197.940 96.480 ;
        RECT 196.945 96.165 197.120 96.200 ;
        RECT 196.190 95.630 196.520 96.030 ;
        RECT 196.945 95.800 197.475 96.165 ;
        RECT 197.665 95.800 197.940 96.310 ;
        RECT 198.110 95.800 198.300 97.160 ;
        RECT 198.470 97.175 198.640 97.840 ;
        RECT 198.810 97.420 198.980 98.180 ;
        RECT 199.215 97.420 199.730 97.830 ;
        RECT 198.470 96.985 199.220 97.175 ;
        RECT 199.390 96.610 199.730 97.420 ;
        RECT 200.820 97.015 201.110 98.180 ;
        RECT 198.500 96.440 199.730 96.610 ;
        RECT 201.280 96.575 201.560 98.010 ;
        RECT 201.730 97.405 202.440 98.180 ;
        RECT 202.610 97.235 202.940 98.010 ;
        RECT 201.790 97.020 202.940 97.235 ;
        RECT 198.480 95.630 198.990 96.165 ;
        RECT 199.210 95.835 199.455 96.440 ;
        RECT 200.820 95.630 201.110 96.355 ;
        RECT 201.280 95.800 201.620 96.575 ;
        RECT 201.790 96.450 202.075 97.020 ;
        RECT 202.260 96.620 202.730 96.850 ;
        RECT 203.135 96.820 203.350 97.935 ;
        RECT 203.530 97.460 203.860 98.180 ;
        RECT 204.500 97.420 205.015 97.830 ;
        RECT 205.250 97.420 205.420 98.180 ;
        RECT 205.590 97.840 207.620 98.010 ;
        RECT 203.640 96.820 203.870 97.160 ;
        RECT 202.900 96.640 203.350 96.820 ;
        RECT 202.900 96.620 203.230 96.640 ;
        RECT 203.540 96.620 203.870 96.820 ;
        RECT 204.500 96.610 204.840 97.420 ;
        RECT 205.590 97.175 205.760 97.840 ;
        RECT 206.155 97.500 207.280 97.670 ;
        RECT 205.010 96.985 205.760 97.175 ;
        RECT 205.930 97.160 206.940 97.330 ;
        RECT 201.790 96.260 202.500 96.450 ;
        RECT 202.200 96.120 202.500 96.260 ;
        RECT 202.690 96.260 203.870 96.450 ;
        RECT 204.500 96.440 205.730 96.610 ;
        RECT 202.690 96.180 203.020 96.260 ;
        RECT 202.200 96.110 202.515 96.120 ;
        RECT 202.200 96.100 202.525 96.110 ;
        RECT 202.200 96.095 202.535 96.100 ;
        RECT 201.790 95.630 201.960 96.090 ;
        RECT 202.200 96.085 202.540 96.095 ;
        RECT 202.200 96.080 202.545 96.085 ;
        RECT 202.200 96.070 202.550 96.080 ;
        RECT 202.200 96.065 202.555 96.070 ;
        RECT 202.200 95.800 202.560 96.065 ;
        RECT 203.190 95.630 203.360 96.090 ;
        RECT 203.530 95.800 203.870 96.260 ;
        RECT 204.775 95.835 205.020 96.440 ;
        RECT 205.240 95.630 205.750 96.165 ;
        RECT 205.930 95.800 206.120 97.160 ;
        RECT 206.290 96.480 206.565 96.960 ;
        RECT 206.290 96.310 206.570 96.480 ;
        RECT 206.770 96.360 206.940 97.160 ;
        RECT 207.110 96.370 207.280 97.500 ;
        RECT 207.450 96.870 207.620 97.840 ;
        RECT 207.790 97.040 207.960 98.180 ;
        RECT 208.130 97.040 208.465 98.010 ;
        RECT 207.450 96.540 207.645 96.870 ;
        RECT 207.870 96.540 208.125 96.870 ;
        RECT 207.870 96.370 208.040 96.540 ;
        RECT 208.295 96.370 208.465 97.040 ;
        RECT 206.290 95.800 206.565 96.310 ;
        RECT 207.110 96.200 208.040 96.370 ;
        RECT 207.110 96.165 207.285 96.200 ;
        RECT 206.755 95.800 207.285 96.165 ;
        RECT 207.710 95.630 208.040 96.030 ;
        RECT 208.210 95.800 208.465 96.370 ;
        RECT 208.640 96.575 208.920 98.010 ;
        RECT 209.090 97.405 209.800 98.180 ;
        RECT 209.970 97.235 210.300 98.010 ;
        RECT 209.150 97.020 210.300 97.235 ;
        RECT 208.640 95.800 208.980 96.575 ;
        RECT 209.150 96.450 209.435 97.020 ;
        RECT 209.620 96.620 210.090 96.850 ;
        RECT 210.495 96.820 210.710 97.935 ;
        RECT 210.890 97.460 211.220 98.180 ;
        RECT 211.000 96.820 211.230 97.160 ;
        RECT 211.400 97.090 214.910 98.180 ;
        RECT 210.260 96.640 210.710 96.820 ;
        RECT 210.260 96.620 210.590 96.640 ;
        RECT 210.900 96.620 211.230 96.820 ;
        RECT 209.150 96.260 209.860 96.450 ;
        RECT 209.560 96.120 209.860 96.260 ;
        RECT 210.050 96.260 211.230 96.450 ;
        RECT 210.050 96.180 210.380 96.260 ;
        RECT 209.560 96.110 209.875 96.120 ;
        RECT 209.560 96.100 209.885 96.110 ;
        RECT 209.560 96.095 209.895 96.100 ;
        RECT 209.150 95.630 209.320 96.090 ;
        RECT 209.560 96.085 209.900 96.095 ;
        RECT 209.560 96.080 209.905 96.085 ;
        RECT 209.560 96.070 209.910 96.080 ;
        RECT 209.560 96.065 209.915 96.070 ;
        RECT 209.560 95.800 209.920 96.065 ;
        RECT 210.550 95.630 210.720 96.090 ;
        RECT 210.890 95.800 211.230 96.260 ;
        RECT 211.400 96.400 213.050 96.920 ;
        RECT 213.220 96.570 214.910 97.090 ;
        RECT 216.090 97.250 216.260 98.010 ;
        RECT 216.440 97.420 216.770 98.180 ;
        RECT 216.090 97.080 216.755 97.250 ;
        RECT 216.940 97.105 217.210 98.010 ;
        RECT 216.585 96.935 216.755 97.080 ;
        RECT 216.020 96.530 216.350 96.900 ;
        RECT 216.585 96.605 216.870 96.935 ;
        RECT 211.400 95.630 214.910 96.400 ;
        RECT 216.585 96.350 216.755 96.605 ;
        RECT 216.090 96.180 216.755 96.350 ;
        RECT 217.040 96.305 217.210 97.105 ;
        RECT 218.305 97.790 218.640 98.010 ;
        RECT 219.645 97.800 220.000 98.180 ;
        RECT 218.305 97.170 218.560 97.790 ;
        RECT 218.810 97.630 219.040 97.670 ;
        RECT 220.170 97.630 220.420 98.010 ;
        RECT 218.810 97.430 220.420 97.630 ;
        RECT 218.810 97.340 218.995 97.430 ;
        RECT 219.585 97.420 220.420 97.430 ;
        RECT 220.670 97.400 220.920 98.180 ;
        RECT 221.090 97.330 221.350 98.010 ;
        RECT 219.150 97.230 219.480 97.260 ;
        RECT 219.150 97.170 220.950 97.230 ;
        RECT 218.305 97.060 221.010 97.170 ;
        RECT 218.305 97.000 219.480 97.060 ;
        RECT 220.810 97.025 221.010 97.060 ;
        RECT 218.300 96.620 218.790 96.820 ;
        RECT 218.980 96.620 219.455 96.830 ;
        RECT 216.090 95.800 216.260 96.180 ;
        RECT 216.440 95.630 216.770 96.010 ;
        RECT 216.950 95.800 217.210 96.305 ;
        RECT 218.305 95.630 218.760 96.395 ;
        RECT 219.235 96.220 219.455 96.620 ;
        RECT 219.700 96.620 220.030 96.830 ;
        RECT 219.700 96.220 219.910 96.620 ;
        RECT 220.200 96.585 220.610 96.890 ;
        RECT 220.840 96.450 221.010 97.025 ;
        RECT 220.740 96.330 221.010 96.450 ;
        RECT 220.165 96.285 221.010 96.330 ;
        RECT 220.165 96.160 220.920 96.285 ;
        RECT 220.165 96.010 220.335 96.160 ;
        RECT 221.180 96.130 221.350 97.330 ;
        RECT 219.035 95.800 220.335 96.010 ;
        RECT 220.590 95.630 220.920 95.990 ;
        RECT 221.090 95.800 221.350 96.130 ;
        RECT 221.520 97.330 221.780 98.010 ;
        RECT 221.950 97.400 222.200 98.180 ;
        RECT 222.450 97.630 222.700 98.010 ;
        RECT 222.870 97.800 223.225 98.180 ;
        RECT 224.230 97.790 224.565 98.010 ;
        RECT 223.830 97.630 224.060 97.670 ;
        RECT 222.450 97.430 224.060 97.630 ;
        RECT 222.450 97.420 223.285 97.430 ;
        RECT 223.875 97.340 224.060 97.430 ;
        RECT 221.520 96.140 221.690 97.330 ;
        RECT 223.390 97.230 223.720 97.260 ;
        RECT 221.920 97.170 223.720 97.230 ;
        RECT 224.310 97.170 224.565 97.790 ;
        RECT 221.860 97.060 224.565 97.170 ;
        RECT 224.740 97.090 226.410 98.180 ;
        RECT 221.860 97.025 222.060 97.060 ;
        RECT 221.860 96.450 222.030 97.025 ;
        RECT 223.390 97.000 224.565 97.060 ;
        RECT 222.260 96.585 222.670 96.890 ;
        RECT 222.840 96.620 223.170 96.830 ;
        RECT 221.860 96.330 222.130 96.450 ;
        RECT 221.860 96.285 222.705 96.330 ;
        RECT 221.950 96.160 222.705 96.285 ;
        RECT 222.960 96.220 223.170 96.620 ;
        RECT 223.415 96.620 223.890 96.830 ;
        RECT 224.080 96.620 224.570 96.820 ;
        RECT 223.415 96.220 223.635 96.620 ;
        RECT 224.740 96.400 225.490 96.920 ;
        RECT 225.660 96.570 226.410 97.090 ;
        RECT 226.580 97.015 226.870 98.180 ;
        RECT 227.045 97.790 227.380 98.010 ;
        RECT 228.385 97.800 228.740 98.180 ;
        RECT 227.045 97.170 227.300 97.790 ;
        RECT 227.550 97.630 227.780 97.670 ;
        RECT 228.910 97.630 229.160 98.010 ;
        RECT 227.550 97.430 229.160 97.630 ;
        RECT 227.550 97.340 227.735 97.430 ;
        RECT 228.325 97.420 229.160 97.430 ;
        RECT 229.410 97.400 229.660 98.180 ;
        RECT 229.830 97.330 230.090 98.010 ;
        RECT 227.890 97.230 228.220 97.260 ;
        RECT 227.890 97.170 229.690 97.230 ;
        RECT 227.045 97.060 229.750 97.170 ;
        RECT 227.045 97.000 228.220 97.060 ;
        RECT 229.550 97.025 229.750 97.060 ;
        RECT 227.040 96.620 227.530 96.820 ;
        RECT 227.720 96.620 228.195 96.830 ;
        RECT 221.520 96.130 221.750 96.140 ;
        RECT 221.520 95.800 221.780 96.130 ;
        RECT 222.535 96.010 222.705 96.160 ;
        RECT 221.950 95.630 222.280 95.990 ;
        RECT 222.535 95.800 223.835 96.010 ;
        RECT 224.110 95.630 224.565 96.395 ;
        RECT 224.740 95.630 226.410 96.400 ;
        RECT 226.580 95.630 226.870 96.355 ;
        RECT 227.045 95.630 227.500 96.395 ;
        RECT 227.975 96.220 228.195 96.620 ;
        RECT 228.440 96.620 228.770 96.830 ;
        RECT 228.440 96.220 228.650 96.620 ;
        RECT 228.940 96.585 229.350 96.890 ;
        RECT 229.580 96.450 229.750 97.025 ;
        RECT 229.480 96.330 229.750 96.450 ;
        RECT 228.905 96.285 229.750 96.330 ;
        RECT 228.905 96.160 229.660 96.285 ;
        RECT 228.905 96.010 229.075 96.160 ;
        RECT 229.920 96.140 230.090 97.330 ;
        RECT 230.260 97.090 233.770 98.180 ;
        RECT 229.860 96.130 230.090 96.140 ;
        RECT 227.775 95.800 229.075 96.010 ;
        RECT 229.330 95.630 229.660 95.990 ;
        RECT 229.830 95.800 230.090 96.130 ;
        RECT 230.260 96.400 231.910 96.920 ;
        RECT 232.080 96.570 233.770 97.090 ;
        RECT 234.865 97.790 235.200 98.010 ;
        RECT 236.205 97.800 236.560 98.180 ;
        RECT 234.865 97.170 235.120 97.790 ;
        RECT 235.370 97.630 235.600 97.670 ;
        RECT 236.730 97.630 236.980 98.010 ;
        RECT 235.370 97.430 236.980 97.630 ;
        RECT 235.370 97.340 235.555 97.430 ;
        RECT 236.145 97.420 236.980 97.430 ;
        RECT 237.230 97.400 237.480 98.180 ;
        RECT 237.650 97.330 237.910 98.010 ;
        RECT 235.710 97.230 236.040 97.260 ;
        RECT 235.710 97.170 237.510 97.230 ;
        RECT 234.865 97.060 237.570 97.170 ;
        RECT 234.865 97.000 236.040 97.060 ;
        RECT 237.370 97.025 237.570 97.060 ;
        RECT 234.860 96.620 235.350 96.820 ;
        RECT 235.540 96.620 236.015 96.830 ;
        RECT 230.260 95.630 233.770 96.400 ;
        RECT 234.865 95.630 235.320 96.395 ;
        RECT 235.795 96.220 236.015 96.620 ;
        RECT 236.260 96.620 236.590 96.830 ;
        RECT 236.260 96.220 236.470 96.620 ;
        RECT 236.760 96.585 237.170 96.890 ;
        RECT 237.400 96.450 237.570 97.025 ;
        RECT 237.300 96.330 237.570 96.450 ;
        RECT 236.725 96.285 237.570 96.330 ;
        RECT 236.725 96.160 237.480 96.285 ;
        RECT 236.725 96.010 236.895 96.160 ;
        RECT 237.740 96.130 237.910 97.330 ;
        RECT 238.170 97.170 238.340 98.010 ;
        RECT 238.510 97.840 239.680 98.010 ;
        RECT 238.510 97.340 238.840 97.840 ;
        RECT 239.350 97.800 239.680 97.840 ;
        RECT 239.870 97.760 240.225 98.180 ;
        RECT 239.010 97.580 239.240 97.670 ;
        RECT 240.395 97.580 240.645 98.010 ;
        RECT 239.010 97.340 240.645 97.580 ;
        RECT 240.815 97.420 241.145 98.180 ;
        RECT 241.315 97.340 241.570 98.010 ;
        RECT 241.760 97.745 247.105 98.180 ;
        RECT 238.170 97.000 241.230 97.170 ;
        RECT 238.085 96.620 238.435 96.830 ;
        RECT 238.605 96.620 239.050 96.820 ;
        RECT 239.220 96.620 239.695 96.820 ;
        RECT 235.595 95.800 236.895 96.010 ;
        RECT 237.150 95.630 237.480 95.990 ;
        RECT 237.650 95.800 237.910 96.130 ;
        RECT 238.170 96.280 239.235 96.450 ;
        RECT 238.170 95.800 238.340 96.280 ;
        RECT 238.510 95.630 238.840 96.110 ;
        RECT 239.065 96.050 239.235 96.280 ;
        RECT 239.415 96.220 239.695 96.620 ;
        RECT 239.965 96.620 240.295 96.820 ;
        RECT 240.465 96.620 240.830 96.820 ;
        RECT 239.965 96.220 240.250 96.620 ;
        RECT 241.060 96.450 241.230 97.000 ;
        RECT 240.430 96.280 241.230 96.450 ;
        RECT 240.430 96.050 240.600 96.280 ;
        RECT 241.400 96.210 241.570 97.340 ;
        RECT 241.385 96.140 241.570 96.210 ;
        RECT 243.345 96.175 243.685 97.005 ;
        RECT 245.165 96.495 245.515 97.745 ;
        RECT 247.280 97.090 250.790 98.180 ;
        RECT 250.960 97.090 252.170 98.180 ;
        RECT 247.280 96.400 248.930 96.920 ;
        RECT 249.100 96.570 250.790 97.090 ;
        RECT 241.360 96.130 241.570 96.140 ;
        RECT 239.065 95.800 240.600 96.050 ;
        RECT 240.770 95.630 241.100 96.110 ;
        RECT 241.315 95.800 241.570 96.130 ;
        RECT 241.760 95.630 247.105 96.175 ;
        RECT 247.280 95.630 250.790 96.400 ;
        RECT 250.960 96.380 251.480 96.920 ;
        RECT 251.650 96.550 252.170 97.090 ;
        RECT 252.340 97.015 252.630 98.180 ;
        RECT 252.800 97.090 254.470 98.180 ;
        RECT 252.800 96.400 253.550 96.920 ;
        RECT 253.720 96.570 254.470 97.090 ;
        RECT 254.645 97.790 254.980 98.010 ;
        RECT 255.985 97.800 256.340 98.180 ;
        RECT 254.645 97.170 254.900 97.790 ;
        RECT 255.150 97.630 255.380 97.670 ;
        RECT 256.510 97.630 256.760 98.010 ;
        RECT 255.150 97.430 256.760 97.630 ;
        RECT 255.150 97.340 255.335 97.430 ;
        RECT 255.925 97.420 256.760 97.430 ;
        RECT 257.010 97.400 257.260 98.180 ;
        RECT 257.430 97.330 257.690 98.010 ;
        RECT 255.490 97.230 255.820 97.260 ;
        RECT 255.490 97.170 257.290 97.230 ;
        RECT 254.645 97.060 257.350 97.170 ;
        RECT 254.645 97.000 255.820 97.060 ;
        RECT 257.150 97.025 257.350 97.060 ;
        RECT 254.640 96.620 255.130 96.820 ;
        RECT 255.320 96.620 255.795 96.830 ;
        RECT 250.960 95.630 252.170 96.380 ;
        RECT 252.340 95.630 252.630 96.355 ;
        RECT 252.800 95.630 254.470 96.400 ;
        RECT 254.645 95.630 255.100 96.395 ;
        RECT 255.575 96.220 255.795 96.620 ;
        RECT 256.040 96.620 256.370 96.830 ;
        RECT 256.040 96.220 256.250 96.620 ;
        RECT 256.540 96.585 256.950 96.890 ;
        RECT 257.180 96.450 257.350 97.025 ;
        RECT 257.080 96.330 257.350 96.450 ;
        RECT 256.505 96.285 257.350 96.330 ;
        RECT 256.505 96.160 257.260 96.285 ;
        RECT 256.505 96.010 256.675 96.160 ;
        RECT 257.520 96.130 257.690 97.330 ;
        RECT 257.950 97.170 258.120 98.010 ;
        RECT 258.290 97.840 259.460 98.010 ;
        RECT 258.290 97.340 258.620 97.840 ;
        RECT 259.130 97.800 259.460 97.840 ;
        RECT 259.650 97.760 260.005 98.180 ;
        RECT 258.790 97.580 259.020 97.670 ;
        RECT 260.175 97.580 260.425 98.010 ;
        RECT 258.790 97.340 260.425 97.580 ;
        RECT 260.595 97.420 260.925 98.180 ;
        RECT 261.095 97.340 261.350 98.010 ;
        RECT 257.950 97.000 261.010 97.170 ;
        RECT 257.865 96.620 258.215 96.830 ;
        RECT 258.385 96.620 258.830 96.820 ;
        RECT 259.000 96.620 259.475 96.820 ;
        RECT 255.375 95.800 256.675 96.010 ;
        RECT 256.930 95.630 257.260 95.990 ;
        RECT 257.430 95.800 257.690 96.130 ;
        RECT 257.950 96.280 259.015 96.450 ;
        RECT 257.950 95.800 258.120 96.280 ;
        RECT 258.290 95.630 258.620 96.110 ;
        RECT 258.845 96.050 259.015 96.280 ;
        RECT 259.195 96.220 259.475 96.620 ;
        RECT 259.745 96.620 260.075 96.820 ;
        RECT 260.245 96.620 260.610 96.820 ;
        RECT 259.745 96.220 260.030 96.620 ;
        RECT 260.840 96.450 261.010 97.000 ;
        RECT 260.210 96.280 261.010 96.450 ;
        RECT 260.210 96.050 260.380 96.280 ;
        RECT 261.180 96.210 261.350 97.340 ;
        RECT 261.545 97.790 261.880 98.010 ;
        RECT 262.885 97.800 263.240 98.180 ;
        RECT 261.545 97.170 261.800 97.790 ;
        RECT 262.050 97.630 262.280 97.670 ;
        RECT 263.410 97.630 263.660 98.010 ;
        RECT 262.050 97.430 263.660 97.630 ;
        RECT 262.050 97.340 262.235 97.430 ;
        RECT 262.825 97.420 263.660 97.430 ;
        RECT 263.910 97.400 264.160 98.180 ;
        RECT 264.330 97.330 264.590 98.010 ;
        RECT 264.765 97.670 266.420 97.960 ;
        RECT 262.390 97.230 262.720 97.260 ;
        RECT 262.390 97.170 264.190 97.230 ;
        RECT 261.545 97.060 264.250 97.170 ;
        RECT 261.545 97.000 262.720 97.060 ;
        RECT 264.050 97.025 264.250 97.060 ;
        RECT 261.540 96.620 262.030 96.820 ;
        RECT 262.220 96.620 262.695 96.830 ;
        RECT 261.165 96.140 261.350 96.210 ;
        RECT 261.140 96.130 261.350 96.140 ;
        RECT 258.845 95.800 260.380 96.050 ;
        RECT 260.550 95.630 260.880 96.110 ;
        RECT 261.095 95.800 261.350 96.130 ;
        RECT 261.545 95.630 262.000 96.395 ;
        RECT 262.475 96.220 262.695 96.620 ;
        RECT 262.940 96.620 263.270 96.830 ;
        RECT 262.940 96.220 263.150 96.620 ;
        RECT 263.440 96.585 263.850 96.890 ;
        RECT 264.080 96.450 264.250 97.025 ;
        RECT 263.980 96.330 264.250 96.450 ;
        RECT 263.405 96.285 264.250 96.330 ;
        RECT 263.405 96.160 264.160 96.285 ;
        RECT 263.405 96.010 263.575 96.160 ;
        RECT 264.420 96.130 264.590 97.330 ;
        RECT 264.765 97.330 266.355 97.500 ;
        RECT 266.590 97.380 266.870 98.180 ;
        RECT 264.765 97.040 265.085 97.330 ;
        RECT 266.185 97.210 266.355 97.330 ;
        RECT 265.280 96.990 265.995 97.160 ;
        RECT 266.185 97.040 266.910 97.210 ;
        RECT 267.080 97.040 267.350 98.010 ;
        RECT 267.520 97.745 272.865 98.180 ;
        RECT 264.765 96.300 265.115 96.870 ;
        RECT 265.285 96.540 265.995 96.990 ;
        RECT 266.740 96.870 266.910 97.040 ;
        RECT 266.165 96.540 266.570 96.870 ;
        RECT 266.740 96.540 267.010 96.870 ;
        RECT 266.740 96.370 266.910 96.540 ;
        RECT 265.300 96.200 266.910 96.370 ;
        RECT 267.180 96.305 267.350 97.040 ;
        RECT 262.275 95.800 263.575 96.010 ;
        RECT 263.830 95.630 264.160 95.990 ;
        RECT 264.330 95.800 264.590 96.130 ;
        RECT 264.770 95.630 265.100 96.130 ;
        RECT 265.300 95.850 265.470 96.200 ;
        RECT 265.670 95.630 266.000 96.030 ;
        RECT 266.170 95.850 266.340 96.200 ;
        RECT 266.510 95.630 266.890 96.030 ;
        RECT 267.080 95.960 267.350 96.305 ;
        RECT 269.105 96.175 269.445 97.005 ;
        RECT 270.925 96.495 271.275 97.745 ;
        RECT 273.500 97.105 273.770 98.010 ;
        RECT 273.940 97.420 274.270 98.180 ;
        RECT 274.450 97.250 274.620 98.010 ;
        RECT 273.500 96.305 273.670 97.105 ;
        RECT 273.955 97.080 274.620 97.250 ;
        RECT 274.880 97.090 277.470 98.180 ;
        RECT 273.955 96.935 274.125 97.080 ;
        RECT 273.840 96.605 274.125 96.935 ;
        RECT 273.955 96.350 274.125 96.605 ;
        RECT 274.360 96.530 274.690 96.900 ;
        RECT 274.880 96.400 276.090 96.920 ;
        RECT 276.260 96.570 277.470 97.090 ;
        RECT 278.100 97.015 278.390 98.180 ;
        RECT 278.565 97.040 278.900 98.010 ;
        RECT 279.070 97.040 279.240 98.180 ;
        RECT 279.410 97.840 281.440 98.010 ;
        RECT 267.520 95.630 272.865 96.175 ;
        RECT 273.500 95.800 273.760 96.305 ;
        RECT 273.955 96.180 274.620 96.350 ;
        RECT 273.940 95.630 274.270 96.010 ;
        RECT 274.450 95.800 274.620 96.180 ;
        RECT 274.880 95.630 277.470 96.400 ;
        RECT 278.565 96.370 278.735 97.040 ;
        RECT 279.410 96.870 279.580 97.840 ;
        RECT 278.905 96.540 279.160 96.870 ;
        RECT 279.385 96.540 279.580 96.870 ;
        RECT 279.750 97.500 280.875 97.670 ;
        RECT 278.990 96.370 279.160 96.540 ;
        RECT 279.750 96.370 279.920 97.500 ;
        RECT 278.100 95.630 278.390 96.355 ;
        RECT 278.565 95.800 278.820 96.370 ;
        RECT 278.990 96.200 279.920 96.370 ;
        RECT 280.090 97.160 281.100 97.330 ;
        RECT 280.090 96.360 280.260 97.160 ;
        RECT 280.465 96.820 280.740 96.960 ;
        RECT 280.460 96.650 280.740 96.820 ;
        RECT 279.745 96.165 279.920 96.200 ;
        RECT 278.990 95.630 279.320 96.030 ;
        RECT 279.745 95.800 280.275 96.165 ;
        RECT 280.465 95.800 280.740 96.650 ;
        RECT 280.910 95.800 281.100 97.160 ;
        RECT 281.270 97.175 281.440 97.840 ;
        RECT 281.610 97.420 281.780 98.180 ;
        RECT 282.015 97.420 282.530 97.830 ;
        RECT 281.270 96.985 282.020 97.175 ;
        RECT 282.190 96.610 282.530 97.420 ;
        RECT 281.300 96.440 282.530 96.610 ;
        RECT 282.705 97.040 283.040 98.010 ;
        RECT 283.210 97.040 283.380 98.180 ;
        RECT 283.550 97.840 285.580 98.010 ;
        RECT 281.280 95.630 281.790 96.165 ;
        RECT 282.010 95.835 282.255 96.440 ;
        RECT 282.705 96.370 282.875 97.040 ;
        RECT 283.550 96.870 283.720 97.840 ;
        RECT 283.045 96.540 283.300 96.870 ;
        RECT 283.525 96.540 283.720 96.870 ;
        RECT 283.890 97.500 285.015 97.670 ;
        RECT 283.130 96.370 283.300 96.540 ;
        RECT 283.890 96.370 284.060 97.500 ;
        RECT 282.705 95.800 282.960 96.370 ;
        RECT 283.130 96.200 284.060 96.370 ;
        RECT 284.230 97.160 285.240 97.330 ;
        RECT 284.230 96.360 284.400 97.160 ;
        RECT 284.605 96.820 284.880 96.960 ;
        RECT 284.600 96.650 284.880 96.820 ;
        RECT 283.885 96.165 284.060 96.200 ;
        RECT 283.130 95.630 283.460 96.030 ;
        RECT 283.885 95.800 284.415 96.165 ;
        RECT 284.605 95.800 284.880 96.650 ;
        RECT 285.050 95.800 285.240 97.160 ;
        RECT 285.410 97.175 285.580 97.840 ;
        RECT 285.750 97.420 285.920 98.180 ;
        RECT 286.155 97.420 286.670 97.830 ;
        RECT 285.410 96.985 286.160 97.175 ;
        RECT 286.330 96.610 286.670 97.420 ;
        RECT 285.440 96.440 286.670 96.610 ;
        RECT 286.845 97.040 287.180 98.010 ;
        RECT 287.350 97.040 287.520 98.180 ;
        RECT 287.690 97.840 289.720 98.010 ;
        RECT 285.420 95.630 285.930 96.165 ;
        RECT 286.150 95.835 286.395 96.440 ;
        RECT 286.845 96.370 287.015 97.040 ;
        RECT 287.690 96.870 287.860 97.840 ;
        RECT 287.185 96.540 287.440 96.870 ;
        RECT 287.665 96.540 287.860 96.870 ;
        RECT 288.030 97.500 289.155 97.670 ;
        RECT 287.270 96.370 287.440 96.540 ;
        RECT 288.030 96.370 288.200 97.500 ;
        RECT 286.845 95.800 287.100 96.370 ;
        RECT 287.270 96.200 288.200 96.370 ;
        RECT 288.370 97.160 289.380 97.330 ;
        RECT 288.370 96.360 288.540 97.160 ;
        RECT 288.745 96.820 289.020 96.960 ;
        RECT 288.740 96.650 289.020 96.820 ;
        RECT 288.025 96.165 288.200 96.200 ;
        RECT 287.270 95.630 287.600 96.030 ;
        RECT 288.025 95.800 288.555 96.165 ;
        RECT 288.745 95.800 289.020 96.650 ;
        RECT 289.190 95.800 289.380 97.160 ;
        RECT 289.550 97.175 289.720 97.840 ;
        RECT 289.890 97.420 290.060 98.180 ;
        RECT 290.295 97.420 290.810 97.830 ;
        RECT 289.550 96.985 290.300 97.175 ;
        RECT 290.470 96.610 290.810 97.420 ;
        RECT 289.580 96.440 290.810 96.610 ;
        RECT 291.905 97.040 292.240 98.010 ;
        RECT 292.410 97.040 292.580 98.180 ;
        RECT 292.750 97.840 294.780 98.010 ;
        RECT 289.560 95.630 290.070 96.165 ;
        RECT 290.290 95.835 290.535 96.440 ;
        RECT 291.905 96.370 292.075 97.040 ;
        RECT 292.750 96.870 292.920 97.840 ;
        RECT 292.245 96.540 292.500 96.870 ;
        RECT 292.725 96.540 292.920 96.870 ;
        RECT 293.090 97.500 294.215 97.670 ;
        RECT 292.330 96.370 292.500 96.540 ;
        RECT 293.090 96.370 293.260 97.500 ;
        RECT 291.905 95.800 292.160 96.370 ;
        RECT 292.330 96.200 293.260 96.370 ;
        RECT 293.430 97.160 294.440 97.330 ;
        RECT 293.430 96.360 293.600 97.160 ;
        RECT 293.805 96.820 294.080 96.960 ;
        RECT 293.800 96.650 294.080 96.820 ;
        RECT 293.085 96.165 293.260 96.200 ;
        RECT 292.330 95.630 292.660 96.030 ;
        RECT 293.085 95.800 293.615 96.165 ;
        RECT 293.805 95.800 294.080 96.650 ;
        RECT 294.250 95.800 294.440 97.160 ;
        RECT 294.610 97.175 294.780 97.840 ;
        RECT 294.950 97.420 295.120 98.180 ;
        RECT 295.355 97.420 295.870 97.830 ;
        RECT 294.610 96.985 295.360 97.175 ;
        RECT 295.530 96.610 295.870 97.420 ;
        RECT 294.640 96.440 295.870 96.610 ;
        RECT 296.500 97.420 297.015 97.830 ;
        RECT 297.250 97.420 297.420 98.180 ;
        RECT 297.590 97.840 299.620 98.010 ;
        RECT 296.500 96.610 296.840 97.420 ;
        RECT 297.590 97.175 297.760 97.840 ;
        RECT 298.155 97.500 299.280 97.670 ;
        RECT 297.010 96.985 297.760 97.175 ;
        RECT 297.930 97.160 298.940 97.330 ;
        RECT 296.500 96.440 297.730 96.610 ;
        RECT 294.620 95.630 295.130 96.165 ;
        RECT 295.350 95.835 295.595 96.440 ;
        RECT 296.775 95.835 297.020 96.440 ;
        RECT 297.240 95.630 297.750 96.165 ;
        RECT 297.930 95.800 298.120 97.160 ;
        RECT 298.290 96.140 298.565 96.960 ;
        RECT 298.770 96.360 298.940 97.160 ;
        RECT 299.110 96.370 299.280 97.500 ;
        RECT 299.450 96.870 299.620 97.840 ;
        RECT 299.790 97.040 299.960 98.180 ;
        RECT 300.130 97.040 300.465 98.010 ;
        RECT 300.730 97.250 300.900 98.010 ;
        RECT 301.080 97.420 301.410 98.180 ;
        RECT 300.730 97.080 301.395 97.250 ;
        RECT 301.580 97.105 301.850 98.010 ;
        RECT 299.450 96.540 299.645 96.870 ;
        RECT 299.870 96.540 300.125 96.870 ;
        RECT 299.870 96.370 300.040 96.540 ;
        RECT 300.295 96.370 300.465 97.040 ;
        RECT 301.225 96.935 301.395 97.080 ;
        RECT 300.660 96.530 300.990 96.900 ;
        RECT 301.225 96.605 301.510 96.935 ;
        RECT 299.110 96.200 300.040 96.370 ;
        RECT 299.110 96.165 299.285 96.200 ;
        RECT 298.290 95.970 298.570 96.140 ;
        RECT 298.290 95.800 298.565 95.970 ;
        RECT 298.755 95.800 299.285 96.165 ;
        RECT 299.710 95.630 300.040 96.030 ;
        RECT 300.210 95.800 300.465 96.370 ;
        RECT 301.225 96.350 301.395 96.605 ;
        RECT 300.730 96.180 301.395 96.350 ;
        RECT 301.680 96.305 301.850 97.105 ;
        RECT 300.730 95.800 300.900 96.180 ;
        RECT 301.080 95.630 301.410 96.010 ;
        RECT 301.590 95.800 301.850 96.305 ;
        RECT 302.020 97.105 302.290 98.010 ;
        RECT 302.460 97.420 302.790 98.180 ;
        RECT 302.970 97.250 303.140 98.010 ;
        RECT 302.020 96.305 302.190 97.105 ;
        RECT 302.475 97.080 303.140 97.250 ;
        RECT 302.475 96.935 302.645 97.080 ;
        RECT 303.860 97.015 304.150 98.180 ;
        RECT 304.320 97.090 307.830 98.180 ;
        RECT 302.360 96.605 302.645 96.935 ;
        RECT 302.475 96.350 302.645 96.605 ;
        RECT 302.880 96.530 303.210 96.900 ;
        RECT 304.320 96.400 305.970 96.920 ;
        RECT 306.140 96.570 307.830 97.090 ;
        RECT 308.090 97.250 308.260 98.010 ;
        RECT 308.475 97.420 308.805 98.180 ;
        RECT 308.090 97.080 308.805 97.250 ;
        RECT 308.975 97.105 309.230 98.010 ;
        RECT 308.000 96.530 308.355 96.900 ;
        RECT 308.635 96.870 308.805 97.080 ;
        RECT 308.635 96.540 308.890 96.870 ;
        RECT 302.020 95.800 302.280 96.305 ;
        RECT 302.475 96.180 303.140 96.350 ;
        RECT 302.460 95.630 302.790 96.010 ;
        RECT 302.970 95.800 303.140 96.180 ;
        RECT 303.860 95.630 304.150 96.355 ;
        RECT 304.320 95.630 307.830 96.400 ;
        RECT 308.635 96.350 308.805 96.540 ;
        RECT 309.060 96.375 309.230 97.105 ;
        RECT 309.405 97.030 309.665 98.180 ;
        RECT 309.840 97.090 311.050 98.180 ;
        RECT 309.840 96.550 310.360 97.090 ;
        RECT 308.090 96.180 308.805 96.350 ;
        RECT 308.090 95.800 308.260 96.180 ;
        RECT 308.475 95.630 308.805 96.010 ;
        RECT 308.975 95.800 309.230 96.375 ;
        RECT 309.405 95.630 309.665 96.470 ;
        RECT 310.530 96.380 311.050 96.920 ;
        RECT 309.840 95.630 311.050 96.380 ;
        RECT 162.095 95.460 311.135 95.630 ;
        RECT 162.180 94.710 163.390 95.460 ;
        RECT 163.620 94.980 163.900 95.460 ;
        RECT 164.070 94.810 164.330 95.200 ;
        RECT 164.505 94.980 164.760 95.460 ;
        RECT 164.930 94.810 165.225 95.200 ;
        RECT 165.405 94.980 165.680 95.460 ;
        RECT 165.850 94.960 166.150 95.290 ;
        RECT 162.180 94.170 162.700 94.710 ;
        RECT 163.575 94.640 165.225 94.810 ;
        RECT 162.870 94.000 163.390 94.540 ;
        RECT 162.180 92.910 163.390 94.000 ;
        RECT 163.575 94.130 163.980 94.640 ;
        RECT 164.150 94.300 165.290 94.470 ;
        RECT 163.575 93.960 164.330 94.130 ;
        RECT 163.615 92.910 163.900 93.780 ;
        RECT 164.070 93.710 164.330 93.960 ;
        RECT 165.120 94.050 165.290 94.300 ;
        RECT 165.460 94.220 165.810 94.790 ;
        RECT 165.980 94.050 166.150 94.960 ;
        RECT 166.320 94.690 167.990 95.460 ;
        RECT 168.625 94.910 168.880 95.200 ;
        RECT 169.050 95.080 169.380 95.460 ;
        RECT 168.625 94.740 169.375 94.910 ;
        RECT 166.320 94.170 167.070 94.690 ;
        RECT 165.120 93.880 166.150 94.050 ;
        RECT 167.240 94.000 167.990 94.520 ;
        RECT 164.070 93.540 165.190 93.710 ;
        RECT 164.070 93.080 164.330 93.540 ;
        RECT 164.505 92.910 164.760 93.370 ;
        RECT 164.930 93.080 165.190 93.540 ;
        RECT 165.360 92.910 165.670 93.710 ;
        RECT 165.840 93.080 166.150 93.880 ;
        RECT 166.320 92.910 167.990 94.000 ;
        RECT 168.625 93.920 168.975 94.570 ;
        RECT 169.145 93.750 169.375 94.740 ;
        RECT 168.625 93.580 169.375 93.750 ;
        RECT 168.625 93.080 168.880 93.580 ;
        RECT 169.050 92.910 169.380 93.410 ;
        RECT 169.550 93.080 169.720 95.200 ;
        RECT 170.080 95.100 170.410 95.460 ;
        RECT 170.580 95.070 171.075 95.240 ;
        RECT 171.280 95.070 172.135 95.240 ;
        RECT 169.950 93.880 170.410 94.930 ;
        RECT 169.890 93.095 170.215 93.880 ;
        RECT 170.580 93.710 170.750 95.070 ;
        RECT 170.920 94.160 171.270 94.780 ;
        RECT 171.440 94.560 171.795 94.780 ;
        RECT 171.440 93.970 171.610 94.560 ;
        RECT 171.965 94.360 172.135 95.070 ;
        RECT 173.010 95.000 173.340 95.460 ;
        RECT 173.550 95.100 173.900 95.270 ;
        RECT 172.340 94.530 173.130 94.780 ;
        RECT 173.550 94.710 173.810 95.100 ;
        RECT 174.120 95.010 175.070 95.290 ;
        RECT 175.240 95.020 175.430 95.460 ;
        RECT 175.600 95.080 176.670 95.250 ;
        RECT 173.300 94.360 173.470 94.540 ;
        RECT 170.580 93.540 170.975 93.710 ;
        RECT 171.145 93.580 171.610 93.970 ;
        RECT 171.780 94.190 173.470 94.360 ;
        RECT 170.805 93.410 170.975 93.540 ;
        RECT 171.780 93.410 171.950 94.190 ;
        RECT 173.640 94.020 173.810 94.710 ;
        RECT 172.310 93.850 173.810 94.020 ;
        RECT 174.000 94.050 174.210 94.840 ;
        RECT 174.380 94.220 174.730 94.840 ;
        RECT 174.900 94.230 175.070 95.010 ;
        RECT 175.600 94.850 175.770 95.080 ;
        RECT 175.240 94.680 175.770 94.850 ;
        RECT 175.240 94.400 175.460 94.680 ;
        RECT 175.940 94.510 176.180 94.910 ;
        RECT 174.900 94.060 175.305 94.230 ;
        RECT 175.640 94.140 176.180 94.510 ;
        RECT 176.350 94.725 176.670 95.080 ;
        RECT 176.915 95.000 177.220 95.460 ;
        RECT 177.390 94.750 177.645 95.280 ;
        RECT 177.820 94.915 183.165 95.460 ;
        RECT 176.350 94.550 176.675 94.725 ;
        RECT 176.350 94.250 177.265 94.550 ;
        RECT 176.525 94.220 177.265 94.250 ;
        RECT 174.000 93.890 174.675 94.050 ;
        RECT 175.135 93.970 175.305 94.060 ;
        RECT 174.000 93.880 174.965 93.890 ;
        RECT 173.640 93.710 173.810 93.850 ;
        RECT 170.385 92.910 170.635 93.370 ;
        RECT 170.805 93.080 171.055 93.410 ;
        RECT 171.270 93.080 171.950 93.410 ;
        RECT 172.120 93.510 173.195 93.680 ;
        RECT 173.640 93.540 174.200 93.710 ;
        RECT 174.505 93.590 174.965 93.880 ;
        RECT 175.135 93.800 176.355 93.970 ;
        RECT 172.120 93.170 172.290 93.510 ;
        RECT 172.525 92.910 172.855 93.340 ;
        RECT 173.025 93.170 173.195 93.510 ;
        RECT 173.490 92.910 173.860 93.370 ;
        RECT 174.030 93.080 174.200 93.540 ;
        RECT 175.135 93.420 175.305 93.800 ;
        RECT 176.525 93.630 176.695 94.220 ;
        RECT 177.435 94.100 177.645 94.750 ;
        RECT 174.435 93.080 175.305 93.420 ;
        RECT 175.895 93.460 176.695 93.630 ;
        RECT 175.475 92.910 175.725 93.370 ;
        RECT 175.895 93.170 176.065 93.460 ;
        RECT 176.245 92.910 176.575 93.290 ;
        RECT 176.915 92.910 177.220 94.050 ;
        RECT 177.390 93.220 177.645 94.100 ;
        RECT 179.405 94.085 179.745 94.915 ;
        RECT 183.340 94.690 185.930 95.460 ;
        RECT 186.100 94.785 186.360 95.290 ;
        RECT 186.540 95.080 186.870 95.460 ;
        RECT 187.050 94.910 187.220 95.290 ;
        RECT 181.225 93.345 181.575 94.595 ;
        RECT 183.340 94.170 184.550 94.690 ;
        RECT 184.720 94.000 185.930 94.520 ;
        RECT 177.820 92.910 183.165 93.345 ;
        RECT 183.340 92.910 185.930 94.000 ;
        RECT 186.100 93.985 186.270 94.785 ;
        RECT 186.555 94.740 187.220 94.910 ;
        RECT 186.555 94.485 186.725 94.740 ;
        RECT 187.940 94.735 188.230 95.460 ;
        RECT 188.405 94.720 188.660 95.290 ;
        RECT 188.830 95.060 189.160 95.460 ;
        RECT 189.585 94.925 190.115 95.290 ;
        RECT 190.305 95.120 190.580 95.290 ;
        RECT 190.300 94.950 190.580 95.120 ;
        RECT 189.585 94.890 189.760 94.925 ;
        RECT 188.830 94.720 189.760 94.890 ;
        RECT 186.440 94.155 186.725 94.485 ;
        RECT 186.960 94.190 187.290 94.560 ;
        RECT 186.555 94.010 186.725 94.155 ;
        RECT 186.100 93.080 186.370 93.985 ;
        RECT 186.555 93.840 187.220 94.010 ;
        RECT 186.540 92.910 186.870 93.670 ;
        RECT 187.050 93.080 187.220 93.840 ;
        RECT 187.940 92.910 188.230 94.075 ;
        RECT 188.405 94.050 188.575 94.720 ;
        RECT 188.830 94.550 189.000 94.720 ;
        RECT 188.745 94.220 189.000 94.550 ;
        RECT 189.225 94.220 189.420 94.550 ;
        RECT 188.405 93.080 188.740 94.050 ;
        RECT 188.910 92.910 189.080 94.050 ;
        RECT 189.250 93.250 189.420 94.220 ;
        RECT 189.590 93.590 189.760 94.720 ;
        RECT 189.930 93.930 190.100 94.730 ;
        RECT 190.305 94.130 190.580 94.950 ;
        RECT 190.750 93.930 190.940 95.290 ;
        RECT 191.120 94.925 191.630 95.460 ;
        RECT 191.850 94.650 192.095 95.255 ;
        RECT 192.540 94.785 192.800 95.290 ;
        RECT 192.980 95.080 193.310 95.460 ;
        RECT 193.490 94.910 193.660 95.290 ;
        RECT 193.920 94.915 199.265 95.460 ;
        RECT 191.140 94.480 192.370 94.650 ;
        RECT 189.930 93.760 190.940 93.930 ;
        RECT 191.110 93.915 191.860 94.105 ;
        RECT 189.590 93.420 190.715 93.590 ;
        RECT 191.110 93.250 191.280 93.915 ;
        RECT 192.030 93.670 192.370 94.480 ;
        RECT 189.250 93.080 191.280 93.250 ;
        RECT 191.450 92.910 191.620 93.670 ;
        RECT 191.855 93.260 192.370 93.670 ;
        RECT 192.540 93.985 192.710 94.785 ;
        RECT 192.995 94.740 193.660 94.910 ;
        RECT 192.995 94.485 193.165 94.740 ;
        RECT 192.880 94.155 193.165 94.485 ;
        RECT 193.400 94.190 193.730 94.560 ;
        RECT 192.995 94.010 193.165 94.155 ;
        RECT 195.505 94.085 195.845 94.915 ;
        RECT 199.440 94.690 201.110 95.460 ;
        RECT 201.280 94.785 201.540 95.290 ;
        RECT 201.720 95.080 202.050 95.460 ;
        RECT 202.230 94.910 202.400 95.290 ;
        RECT 202.660 94.915 208.005 95.460 ;
        RECT 208.180 94.915 213.525 95.460 ;
        RECT 192.540 93.080 192.810 93.985 ;
        RECT 192.995 93.840 193.660 94.010 ;
        RECT 192.980 92.910 193.310 93.670 ;
        RECT 193.490 93.080 193.660 93.840 ;
        RECT 197.325 93.345 197.675 94.595 ;
        RECT 199.440 94.170 200.190 94.690 ;
        RECT 200.360 94.000 201.110 94.520 ;
        RECT 193.920 92.910 199.265 93.345 ;
        RECT 199.440 92.910 201.110 94.000 ;
        RECT 201.280 93.985 201.450 94.785 ;
        RECT 201.735 94.740 202.400 94.910 ;
        RECT 201.735 94.485 201.905 94.740 ;
        RECT 201.620 94.155 201.905 94.485 ;
        RECT 202.140 94.190 202.470 94.560 ;
        RECT 201.735 94.010 201.905 94.155 ;
        RECT 204.245 94.085 204.585 94.915 ;
        RECT 201.280 93.080 201.550 93.985 ;
        RECT 201.735 93.840 202.400 94.010 ;
        RECT 201.720 92.910 202.050 93.670 ;
        RECT 202.230 93.080 202.400 93.840 ;
        RECT 206.065 93.345 206.415 94.595 ;
        RECT 209.765 94.085 210.105 94.915 ;
        RECT 213.700 94.735 213.990 95.460 ;
        RECT 214.160 94.690 216.750 95.460 ;
        RECT 217.010 94.810 217.180 95.290 ;
        RECT 217.350 94.980 217.680 95.460 ;
        RECT 217.905 95.040 219.440 95.290 ;
        RECT 217.905 94.810 218.075 95.040 ;
        RECT 211.585 93.345 211.935 94.595 ;
        RECT 214.160 94.170 215.370 94.690 ;
        RECT 217.010 94.640 218.075 94.810 ;
        RECT 202.660 92.910 208.005 93.345 ;
        RECT 208.180 92.910 213.525 93.345 ;
        RECT 213.700 92.910 213.990 94.075 ;
        RECT 215.540 94.000 216.750 94.520 ;
        RECT 218.255 94.470 218.535 94.870 ;
        RECT 216.925 94.260 217.275 94.470 ;
        RECT 217.445 94.270 217.890 94.470 ;
        RECT 218.060 94.270 218.535 94.470 ;
        RECT 218.805 94.470 219.090 94.870 ;
        RECT 219.270 94.810 219.440 95.040 ;
        RECT 219.610 94.980 219.940 95.460 ;
        RECT 220.155 94.960 220.410 95.290 ;
        RECT 220.200 94.950 220.410 94.960 ;
        RECT 220.225 94.880 220.410 94.950 ;
        RECT 219.270 94.640 220.070 94.810 ;
        RECT 218.805 94.270 219.135 94.470 ;
        RECT 219.305 94.440 219.670 94.470 ;
        RECT 219.305 94.270 219.680 94.440 ;
        RECT 219.900 94.090 220.070 94.640 ;
        RECT 214.160 92.910 216.750 94.000 ;
        RECT 217.010 93.920 220.070 94.090 ;
        RECT 217.010 93.080 217.180 93.920 ;
        RECT 220.240 93.750 220.410 94.880 ;
        RECT 220.615 94.890 220.870 95.240 ;
        RECT 221.040 95.060 221.370 95.460 ;
        RECT 221.540 94.890 221.710 95.240 ;
        RECT 221.880 95.060 222.260 95.460 ;
        RECT 220.615 94.720 222.280 94.890 ;
        RECT 222.450 94.785 222.725 95.130 ;
        RECT 222.110 94.550 222.280 94.720 ;
        RECT 220.600 94.220 220.945 94.550 ;
        RECT 221.115 94.220 221.940 94.550 ;
        RECT 222.110 94.220 222.385 94.550 ;
        RECT 217.350 93.250 217.680 93.750 ;
        RECT 217.850 93.510 219.485 93.750 ;
        RECT 217.850 93.420 218.080 93.510 ;
        RECT 218.190 93.250 218.520 93.290 ;
        RECT 217.350 93.080 218.520 93.250 ;
        RECT 218.710 92.910 219.065 93.330 ;
        RECT 219.235 93.080 219.485 93.510 ;
        RECT 219.655 92.910 219.985 93.670 ;
        RECT 220.155 93.080 220.410 93.750 ;
        RECT 220.620 93.760 220.945 94.050 ;
        RECT 221.115 93.930 221.310 94.220 ;
        RECT 222.110 94.050 222.280 94.220 ;
        RECT 222.555 94.050 222.725 94.785 ;
        RECT 222.910 94.740 223.240 95.460 ;
        RECT 223.785 95.060 225.400 95.230 ;
        RECT 225.570 95.060 225.900 95.460 ;
        RECT 225.230 94.890 225.400 95.060 ;
        RECT 226.070 94.985 226.405 95.245 ;
        RECT 222.965 94.220 223.315 94.550 ;
        RECT 223.625 94.220 224.045 94.885 ;
        RECT 224.215 94.440 224.505 94.880 ;
        RECT 224.695 94.440 224.965 94.880 ;
        RECT 225.230 94.720 225.790 94.890 ;
        RECT 225.620 94.550 225.790 94.720 ;
        RECT 225.175 94.440 225.425 94.550 ;
        RECT 224.215 94.270 224.510 94.440 ;
        RECT 224.695 94.270 224.970 94.440 ;
        RECT 225.175 94.270 225.430 94.440 ;
        RECT 224.215 94.220 224.505 94.270 ;
        RECT 224.695 94.220 224.965 94.270 ;
        RECT 225.175 94.220 225.425 94.270 ;
        RECT 225.620 94.220 225.925 94.550 ;
        RECT 222.965 94.100 223.170 94.220 ;
        RECT 221.620 93.880 222.280 94.050 ;
        RECT 221.620 93.760 221.790 93.880 ;
        RECT 220.620 93.590 221.790 93.760 ;
        RECT 220.600 93.130 221.790 93.420 ;
        RECT 221.960 92.910 222.240 93.710 ;
        RECT 222.450 93.080 222.725 94.050 ;
        RECT 222.960 93.930 223.170 94.100 ;
        RECT 225.620 94.050 225.790 94.220 ;
        RECT 223.420 93.880 225.790 94.050 ;
        RECT 222.990 93.250 223.160 93.750 ;
        RECT 223.420 93.420 223.590 93.880 ;
        RECT 223.820 93.500 225.245 93.670 ;
        RECT 223.820 93.250 224.150 93.500 ;
        RECT 222.990 93.080 224.150 93.250 ;
        RECT 224.375 92.910 224.705 93.330 ;
        RECT 224.960 93.080 225.245 93.500 ;
        RECT 225.490 92.910 225.820 93.710 ;
        RECT 226.150 93.630 226.405 94.985 ;
        RECT 226.590 94.960 226.920 95.460 ;
        RECT 227.120 94.890 227.290 95.240 ;
        RECT 227.490 95.060 227.820 95.460 ;
        RECT 227.990 94.890 228.160 95.240 ;
        RECT 228.330 95.060 228.710 95.460 ;
        RECT 226.585 94.220 226.935 94.790 ;
        RECT 227.120 94.720 228.730 94.890 ;
        RECT 228.900 94.785 229.170 95.130 ;
        RECT 229.340 94.915 234.685 95.460 ;
        RECT 228.560 94.550 228.730 94.720 ;
        RECT 226.070 93.120 226.405 93.630 ;
        RECT 226.585 93.760 226.905 94.050 ;
        RECT 227.105 93.930 227.815 94.550 ;
        RECT 227.985 94.220 228.390 94.550 ;
        RECT 228.560 94.220 228.830 94.550 ;
        RECT 228.560 94.050 228.730 94.220 ;
        RECT 229.000 94.050 229.170 94.785 ;
        RECT 230.925 94.085 231.265 94.915 ;
        RECT 235.870 94.810 236.040 95.290 ;
        RECT 236.210 94.980 236.540 95.460 ;
        RECT 236.765 95.040 238.300 95.290 ;
        RECT 236.765 94.810 236.935 95.040 ;
        RECT 235.870 94.640 236.935 94.810 ;
        RECT 228.005 93.880 228.730 94.050 ;
        RECT 228.005 93.760 228.175 93.880 ;
        RECT 226.585 93.590 228.175 93.760 ;
        RECT 226.585 93.130 228.240 93.420 ;
        RECT 228.410 92.910 228.690 93.710 ;
        RECT 228.900 93.080 229.170 94.050 ;
        RECT 232.745 93.345 233.095 94.595 ;
        RECT 237.115 94.470 237.395 94.870 ;
        RECT 235.785 94.260 236.135 94.470 ;
        RECT 236.305 94.270 236.750 94.470 ;
        RECT 236.920 94.270 237.395 94.470 ;
        RECT 237.665 94.470 237.950 94.870 ;
        RECT 238.130 94.810 238.300 95.040 ;
        RECT 238.470 94.980 238.800 95.460 ;
        RECT 239.015 94.960 239.270 95.290 ;
        RECT 239.085 94.880 239.270 94.960 ;
        RECT 238.130 94.640 238.930 94.810 ;
        RECT 237.665 94.270 237.995 94.470 ;
        RECT 238.165 94.270 238.530 94.470 ;
        RECT 238.760 94.090 238.930 94.640 ;
        RECT 235.870 93.920 238.930 94.090 ;
        RECT 229.340 92.910 234.685 93.345 ;
        RECT 235.870 93.080 236.040 93.920 ;
        RECT 239.100 93.750 239.270 94.880 ;
        RECT 239.460 94.735 239.750 95.460 ;
        RECT 240.010 94.810 240.180 95.290 ;
        RECT 240.350 94.980 240.680 95.460 ;
        RECT 240.905 95.040 242.440 95.290 ;
        RECT 240.905 94.810 241.075 95.040 ;
        RECT 240.010 94.640 241.075 94.810 ;
        RECT 241.255 94.470 241.535 94.870 ;
        RECT 239.925 94.260 240.275 94.470 ;
        RECT 240.445 94.270 240.890 94.470 ;
        RECT 241.060 94.270 241.535 94.470 ;
        RECT 241.805 94.470 242.090 94.870 ;
        RECT 242.270 94.810 242.440 95.040 ;
        RECT 242.610 94.980 242.940 95.460 ;
        RECT 243.155 94.960 243.410 95.290 ;
        RECT 243.200 94.950 243.410 94.960 ;
        RECT 243.225 94.880 243.410 94.950 ;
        RECT 242.270 94.640 243.070 94.810 ;
        RECT 241.805 94.270 242.135 94.470 ;
        RECT 242.305 94.270 242.670 94.470 ;
        RECT 242.900 94.090 243.070 94.640 ;
        RECT 236.210 93.250 236.540 93.750 ;
        RECT 236.710 93.510 238.345 93.750 ;
        RECT 236.710 93.420 236.940 93.510 ;
        RECT 237.050 93.250 237.380 93.290 ;
        RECT 236.210 93.080 237.380 93.250 ;
        RECT 237.570 92.910 237.925 93.330 ;
        RECT 238.095 93.080 238.345 93.510 ;
        RECT 238.515 92.910 238.845 93.670 ;
        RECT 239.015 93.080 239.270 93.750 ;
        RECT 239.460 92.910 239.750 94.075 ;
        RECT 240.010 93.920 243.070 94.090 ;
        RECT 240.010 93.080 240.180 93.920 ;
        RECT 243.240 93.750 243.410 94.880 ;
        RECT 240.350 93.250 240.680 93.750 ;
        RECT 240.850 93.510 242.485 93.750 ;
        RECT 240.850 93.420 241.080 93.510 ;
        RECT 241.190 93.250 241.520 93.290 ;
        RECT 240.350 93.080 241.520 93.250 ;
        RECT 241.710 92.910 242.065 93.330 ;
        RECT 242.235 93.080 242.485 93.510 ;
        RECT 242.655 92.910 242.985 93.670 ;
        RECT 243.155 93.080 243.410 93.750 ;
        RECT 243.600 94.960 243.860 95.290 ;
        RECT 244.030 95.100 244.360 95.460 ;
        RECT 244.615 95.080 245.915 95.290 ;
        RECT 243.600 93.760 243.770 94.960 ;
        RECT 244.615 94.930 244.785 95.080 ;
        RECT 244.030 94.805 244.785 94.930 ;
        RECT 243.940 94.760 244.785 94.805 ;
        RECT 243.940 94.640 244.210 94.760 ;
        RECT 243.940 94.065 244.110 94.640 ;
        RECT 244.340 94.200 244.750 94.505 ;
        RECT 245.040 94.470 245.250 94.870 ;
        RECT 244.920 94.260 245.250 94.470 ;
        RECT 245.495 94.470 245.715 94.870 ;
        RECT 246.190 94.695 246.645 95.460 ;
        RECT 246.820 94.915 252.165 95.460 ;
        RECT 252.340 94.915 257.685 95.460 ;
        RECT 245.495 94.260 245.970 94.470 ;
        RECT 246.160 94.270 246.650 94.470 ;
        RECT 243.940 94.030 244.140 94.065 ;
        RECT 245.470 94.030 246.645 94.090 ;
        RECT 248.405 94.085 248.745 94.915 ;
        RECT 243.940 93.920 246.645 94.030 ;
        RECT 244.000 93.860 245.800 93.920 ;
        RECT 245.470 93.830 245.800 93.860 ;
        RECT 243.600 93.080 243.860 93.760 ;
        RECT 244.030 92.910 244.280 93.690 ;
        RECT 244.530 93.660 245.365 93.670 ;
        RECT 245.955 93.660 246.140 93.750 ;
        RECT 244.530 93.460 246.140 93.660 ;
        RECT 244.530 93.080 244.780 93.460 ;
        RECT 245.910 93.420 246.140 93.460 ;
        RECT 246.390 93.300 246.645 93.920 ;
        RECT 250.225 93.345 250.575 94.595 ;
        RECT 253.925 94.085 254.265 94.915 ;
        RECT 257.950 94.810 258.120 95.290 ;
        RECT 258.290 94.980 258.620 95.460 ;
        RECT 258.845 95.040 260.380 95.290 ;
        RECT 258.845 94.810 259.015 95.040 ;
        RECT 257.950 94.640 259.015 94.810 ;
        RECT 255.745 93.345 256.095 94.595 ;
        RECT 259.195 94.470 259.475 94.870 ;
        RECT 257.865 94.260 258.215 94.470 ;
        RECT 258.385 94.270 258.830 94.470 ;
        RECT 259.000 94.270 259.475 94.470 ;
        RECT 259.745 94.470 260.030 94.870 ;
        RECT 260.210 94.810 260.380 95.040 ;
        RECT 260.550 94.980 260.880 95.460 ;
        RECT 261.095 94.960 261.350 95.290 ;
        RECT 261.140 94.950 261.350 94.960 ;
        RECT 261.165 94.880 261.350 94.950 ;
        RECT 260.210 94.640 261.010 94.810 ;
        RECT 259.745 94.270 260.075 94.470 ;
        RECT 260.245 94.270 260.610 94.470 ;
        RECT 260.840 94.090 261.010 94.640 ;
        RECT 257.950 93.920 261.010 94.090 ;
        RECT 244.950 92.910 245.305 93.290 ;
        RECT 246.310 93.080 246.645 93.300 ;
        RECT 246.820 92.910 252.165 93.345 ;
        RECT 252.340 92.910 257.685 93.345 ;
        RECT 257.950 93.080 258.120 93.920 ;
        RECT 261.180 93.750 261.350 94.880 ;
        RECT 261.545 94.695 262.000 95.460 ;
        RECT 262.275 95.080 263.575 95.290 ;
        RECT 263.830 95.100 264.160 95.460 ;
        RECT 263.405 94.930 263.575 95.080 ;
        RECT 264.330 94.960 264.590 95.290 ;
        RECT 262.475 94.470 262.695 94.870 ;
        RECT 261.540 94.270 262.030 94.470 ;
        RECT 262.220 94.260 262.695 94.470 ;
        RECT 262.940 94.470 263.150 94.870 ;
        RECT 263.405 94.805 264.160 94.930 ;
        RECT 263.405 94.760 264.250 94.805 ;
        RECT 263.980 94.640 264.250 94.760 ;
        RECT 262.940 94.260 263.270 94.470 ;
        RECT 263.440 94.200 263.850 94.505 ;
        RECT 258.290 93.250 258.620 93.750 ;
        RECT 258.790 93.510 260.425 93.750 ;
        RECT 258.790 93.420 259.020 93.510 ;
        RECT 259.130 93.250 259.460 93.290 ;
        RECT 258.290 93.080 259.460 93.250 ;
        RECT 259.650 92.910 260.005 93.330 ;
        RECT 260.175 93.080 260.425 93.510 ;
        RECT 260.595 92.910 260.925 93.670 ;
        RECT 261.095 93.080 261.350 93.750 ;
        RECT 261.545 94.030 262.720 94.090 ;
        RECT 264.080 94.065 264.250 94.640 ;
        RECT 264.050 94.030 264.250 94.065 ;
        RECT 261.545 93.920 264.250 94.030 ;
        RECT 261.545 93.300 261.800 93.920 ;
        RECT 262.390 93.860 264.190 93.920 ;
        RECT 262.390 93.830 262.720 93.860 ;
        RECT 264.420 93.760 264.590 94.960 ;
        RECT 265.220 94.735 265.510 95.460 ;
        RECT 265.680 94.915 271.025 95.460 ;
        RECT 271.200 94.915 276.545 95.460 ;
        RECT 267.265 94.085 267.605 94.915 ;
        RECT 262.050 93.660 262.235 93.750 ;
        RECT 262.825 93.660 263.660 93.670 ;
        RECT 262.050 93.460 263.660 93.660 ;
        RECT 262.050 93.420 262.280 93.460 ;
        RECT 261.545 93.080 261.880 93.300 ;
        RECT 262.885 92.910 263.240 93.290 ;
        RECT 263.410 93.080 263.660 93.460 ;
        RECT 263.910 92.910 264.160 93.690 ;
        RECT 264.330 93.080 264.590 93.760 ;
        RECT 265.220 92.910 265.510 94.075 ;
        RECT 269.085 93.345 269.435 94.595 ;
        RECT 272.785 94.085 273.125 94.915 ;
        RECT 277.640 94.830 277.980 95.290 ;
        RECT 278.150 95.000 278.320 95.460 ;
        RECT 278.950 95.025 279.310 95.290 ;
        RECT 278.955 95.020 279.310 95.025 ;
        RECT 278.960 95.010 279.310 95.020 ;
        RECT 278.965 95.005 279.310 95.010 ;
        RECT 278.970 94.995 279.310 95.005 ;
        RECT 279.550 95.000 279.720 95.460 ;
        RECT 278.975 94.990 279.310 94.995 ;
        RECT 278.985 94.980 279.310 94.990 ;
        RECT 278.995 94.970 279.310 94.980 ;
        RECT 278.490 94.830 278.820 94.910 ;
        RECT 277.640 94.640 278.820 94.830 ;
        RECT 279.010 94.830 279.310 94.970 ;
        RECT 279.010 94.640 279.720 94.830 ;
        RECT 274.605 93.345 274.955 94.595 ;
        RECT 277.640 94.270 277.970 94.470 ;
        RECT 278.280 94.450 278.610 94.470 ;
        RECT 278.160 94.270 278.610 94.450 ;
        RECT 277.640 93.930 277.870 94.270 ;
        RECT 265.680 92.910 271.025 93.345 ;
        RECT 271.200 92.910 276.545 93.345 ;
        RECT 277.650 92.910 277.980 93.630 ;
        RECT 278.160 93.155 278.375 94.270 ;
        RECT 278.780 94.240 279.250 94.470 ;
        RECT 279.435 94.070 279.720 94.640 ;
        RECT 279.890 94.515 280.230 95.290 ;
        RECT 280.400 94.830 280.740 95.290 ;
        RECT 280.910 95.000 281.080 95.460 ;
        RECT 281.710 95.025 282.070 95.290 ;
        RECT 281.715 95.020 282.070 95.025 ;
        RECT 281.720 95.010 282.070 95.020 ;
        RECT 281.725 95.005 282.070 95.010 ;
        RECT 281.730 94.995 282.070 95.005 ;
        RECT 282.310 95.000 282.480 95.460 ;
        RECT 281.735 94.990 282.070 94.995 ;
        RECT 281.745 94.980 282.070 94.990 ;
        RECT 281.755 94.970 282.070 94.980 ;
        RECT 281.250 94.830 281.580 94.910 ;
        RECT 280.400 94.640 281.580 94.830 ;
        RECT 281.770 94.830 282.070 94.970 ;
        RECT 281.770 94.640 282.480 94.830 ;
        RECT 278.570 93.855 279.720 94.070 ;
        RECT 278.570 93.080 278.900 93.855 ;
        RECT 279.070 92.910 279.780 93.685 ;
        RECT 279.950 93.080 280.230 94.515 ;
        RECT 280.400 94.270 280.730 94.470 ;
        RECT 281.040 94.450 281.370 94.470 ;
        RECT 280.920 94.270 281.370 94.450 ;
        RECT 280.400 93.930 280.630 94.270 ;
        RECT 280.410 92.910 280.740 93.630 ;
        RECT 280.920 93.155 281.135 94.270 ;
        RECT 281.540 94.240 282.010 94.470 ;
        RECT 282.195 94.070 282.480 94.640 ;
        RECT 282.650 94.515 282.990 95.290 ;
        RECT 281.330 93.855 282.480 94.070 ;
        RECT 281.330 93.080 281.660 93.855 ;
        RECT 281.830 92.910 282.540 93.685 ;
        RECT 282.710 93.080 282.990 94.515 ;
        RECT 283.160 94.785 283.420 95.290 ;
        RECT 283.600 95.080 283.930 95.460 ;
        RECT 284.110 94.910 284.280 95.290 ;
        RECT 283.160 93.985 283.330 94.785 ;
        RECT 283.615 94.740 284.280 94.910 ;
        RECT 283.615 94.485 283.785 94.740 ;
        RECT 284.540 94.690 288.050 95.460 ;
        RECT 288.220 94.710 289.430 95.460 ;
        RECT 289.690 94.910 289.860 95.290 ;
        RECT 290.040 95.080 290.370 95.460 ;
        RECT 289.690 94.740 290.355 94.910 ;
        RECT 290.550 94.785 290.810 95.290 ;
        RECT 283.500 94.155 283.785 94.485 ;
        RECT 284.020 94.190 284.350 94.560 ;
        RECT 284.540 94.170 286.190 94.690 ;
        RECT 283.615 94.010 283.785 94.155 ;
        RECT 283.160 93.080 283.430 93.985 ;
        RECT 283.615 93.840 284.280 94.010 ;
        RECT 286.360 94.000 288.050 94.520 ;
        RECT 288.220 94.170 288.740 94.710 ;
        RECT 288.910 94.000 289.430 94.540 ;
        RECT 289.620 94.190 289.950 94.560 ;
        RECT 290.185 94.485 290.355 94.740 ;
        RECT 290.185 94.155 290.470 94.485 ;
        RECT 290.185 94.010 290.355 94.155 ;
        RECT 283.600 92.910 283.930 93.670 ;
        RECT 284.110 93.080 284.280 93.840 ;
        RECT 284.540 92.910 288.050 94.000 ;
        RECT 288.220 92.910 289.430 94.000 ;
        RECT 289.690 93.840 290.355 94.010 ;
        RECT 290.640 93.985 290.810 94.785 ;
        RECT 290.980 94.735 291.270 95.460 ;
        RECT 291.445 94.750 291.700 95.280 ;
        RECT 291.870 95.000 292.175 95.460 ;
        RECT 292.420 95.080 293.490 95.250 ;
        RECT 291.445 94.100 291.655 94.750 ;
        RECT 292.420 94.725 292.740 95.080 ;
        RECT 292.415 94.550 292.740 94.725 ;
        RECT 291.825 94.250 292.740 94.550 ;
        RECT 292.910 94.510 293.150 94.910 ;
        RECT 293.320 94.850 293.490 95.080 ;
        RECT 293.660 95.020 293.850 95.460 ;
        RECT 294.020 95.010 294.970 95.290 ;
        RECT 295.190 95.100 295.540 95.270 ;
        RECT 293.320 94.680 293.850 94.850 ;
        RECT 291.825 94.220 292.565 94.250 ;
        RECT 289.690 93.080 289.860 93.840 ;
        RECT 290.040 92.910 290.370 93.670 ;
        RECT 290.540 93.080 290.810 93.985 ;
        RECT 290.980 92.910 291.270 94.075 ;
        RECT 291.445 93.220 291.700 94.100 ;
        RECT 291.870 92.910 292.175 94.050 ;
        RECT 292.395 93.630 292.565 94.220 ;
        RECT 292.910 94.140 293.450 94.510 ;
        RECT 293.630 94.400 293.850 94.680 ;
        RECT 294.020 94.230 294.190 95.010 ;
        RECT 293.785 94.060 294.190 94.230 ;
        RECT 294.360 94.220 294.710 94.840 ;
        RECT 293.785 93.970 293.955 94.060 ;
        RECT 294.880 94.050 295.090 94.840 ;
        RECT 292.735 93.800 293.955 93.970 ;
        RECT 294.415 93.890 295.090 94.050 ;
        RECT 292.395 93.460 293.195 93.630 ;
        RECT 292.515 92.910 292.845 93.290 ;
        RECT 293.025 93.170 293.195 93.460 ;
        RECT 293.785 93.420 293.955 93.800 ;
        RECT 294.125 93.880 295.090 93.890 ;
        RECT 295.280 94.710 295.540 95.100 ;
        RECT 295.750 95.000 296.080 95.460 ;
        RECT 296.955 95.070 297.810 95.240 ;
        RECT 298.015 95.070 298.510 95.240 ;
        RECT 298.680 95.100 299.010 95.460 ;
        RECT 295.280 94.020 295.450 94.710 ;
        RECT 295.620 94.360 295.790 94.540 ;
        RECT 295.960 94.530 296.750 94.780 ;
        RECT 296.955 94.360 297.125 95.070 ;
        RECT 297.295 94.560 297.650 94.780 ;
        RECT 295.620 94.190 297.310 94.360 ;
        RECT 294.125 93.590 294.585 93.880 ;
        RECT 295.280 93.850 296.780 94.020 ;
        RECT 295.280 93.710 295.450 93.850 ;
        RECT 294.890 93.540 295.450 93.710 ;
        RECT 293.365 92.910 293.615 93.370 ;
        RECT 293.785 93.080 294.655 93.420 ;
        RECT 294.890 93.080 295.060 93.540 ;
        RECT 295.895 93.510 296.970 93.680 ;
        RECT 295.230 92.910 295.600 93.370 ;
        RECT 295.895 93.170 296.065 93.510 ;
        RECT 296.235 92.910 296.565 93.340 ;
        RECT 296.800 93.170 296.970 93.510 ;
        RECT 297.140 93.410 297.310 94.190 ;
        RECT 297.480 93.970 297.650 94.560 ;
        RECT 297.820 94.160 298.170 94.780 ;
        RECT 297.480 93.580 297.945 93.970 ;
        RECT 298.340 93.710 298.510 95.070 ;
        RECT 298.680 93.880 299.140 94.930 ;
        RECT 298.115 93.540 298.510 93.710 ;
        RECT 298.115 93.410 298.285 93.540 ;
        RECT 297.140 93.080 297.820 93.410 ;
        RECT 298.035 93.080 298.285 93.410 ;
        RECT 298.455 92.910 298.705 93.370 ;
        RECT 298.875 93.095 299.200 93.880 ;
        RECT 299.370 93.080 299.540 95.200 ;
        RECT 299.710 95.080 300.040 95.460 ;
        RECT 300.210 94.910 300.465 95.200 ;
        RECT 299.715 94.740 300.465 94.910 ;
        RECT 300.645 94.910 300.900 95.200 ;
        RECT 301.070 95.080 301.400 95.460 ;
        RECT 300.645 94.740 301.395 94.910 ;
        RECT 299.715 93.750 299.945 94.740 ;
        RECT 300.115 93.920 300.465 94.570 ;
        RECT 300.645 93.920 300.995 94.570 ;
        RECT 301.165 93.750 301.395 94.740 ;
        RECT 299.715 93.580 300.465 93.750 ;
        RECT 299.710 92.910 300.040 93.410 ;
        RECT 300.210 93.080 300.465 93.580 ;
        RECT 300.645 93.580 301.395 93.750 ;
        RECT 300.645 93.080 300.900 93.580 ;
        RECT 301.070 92.910 301.400 93.410 ;
        RECT 301.570 93.080 301.740 95.200 ;
        RECT 302.100 95.100 302.430 95.460 ;
        RECT 302.600 95.070 303.095 95.240 ;
        RECT 303.300 95.070 304.155 95.240 ;
        RECT 301.970 93.880 302.430 94.930 ;
        RECT 301.910 93.095 302.235 93.880 ;
        RECT 302.600 93.710 302.770 95.070 ;
        RECT 302.940 94.160 303.290 94.780 ;
        RECT 303.460 94.560 303.815 94.780 ;
        RECT 303.460 93.970 303.630 94.560 ;
        RECT 303.985 94.360 304.155 95.070 ;
        RECT 305.030 95.000 305.360 95.460 ;
        RECT 305.570 95.100 305.920 95.270 ;
        RECT 304.360 94.530 305.150 94.780 ;
        RECT 305.570 94.710 305.830 95.100 ;
        RECT 306.140 95.010 307.090 95.290 ;
        RECT 307.260 95.020 307.450 95.460 ;
        RECT 307.620 95.080 308.690 95.250 ;
        RECT 305.320 94.360 305.490 94.540 ;
        RECT 302.600 93.540 302.995 93.710 ;
        RECT 303.165 93.580 303.630 93.970 ;
        RECT 303.800 94.190 305.490 94.360 ;
        RECT 302.825 93.410 302.995 93.540 ;
        RECT 303.800 93.410 303.970 94.190 ;
        RECT 305.660 94.020 305.830 94.710 ;
        RECT 304.330 93.850 305.830 94.020 ;
        RECT 306.020 94.050 306.230 94.840 ;
        RECT 306.400 94.220 306.750 94.840 ;
        RECT 306.920 94.230 307.090 95.010 ;
        RECT 307.620 94.850 307.790 95.080 ;
        RECT 307.260 94.680 307.790 94.850 ;
        RECT 307.260 94.400 307.480 94.680 ;
        RECT 307.960 94.510 308.200 94.910 ;
        RECT 306.920 94.060 307.325 94.230 ;
        RECT 307.660 94.140 308.200 94.510 ;
        RECT 308.370 94.725 308.690 95.080 ;
        RECT 308.935 95.000 309.240 95.460 ;
        RECT 309.410 94.750 309.665 95.280 ;
        RECT 308.370 94.550 308.695 94.725 ;
        RECT 308.370 94.250 309.285 94.550 ;
        RECT 308.545 94.220 309.285 94.250 ;
        RECT 306.020 93.890 306.695 94.050 ;
        RECT 307.155 93.970 307.325 94.060 ;
        RECT 306.020 93.880 306.985 93.890 ;
        RECT 305.660 93.710 305.830 93.850 ;
        RECT 302.405 92.910 302.655 93.370 ;
        RECT 302.825 93.080 303.075 93.410 ;
        RECT 303.290 93.080 303.970 93.410 ;
        RECT 304.140 93.510 305.215 93.680 ;
        RECT 305.660 93.540 306.220 93.710 ;
        RECT 306.525 93.590 306.985 93.880 ;
        RECT 307.155 93.800 308.375 93.970 ;
        RECT 304.140 93.170 304.310 93.510 ;
        RECT 304.545 92.910 304.875 93.340 ;
        RECT 305.045 93.170 305.215 93.510 ;
        RECT 305.510 92.910 305.880 93.370 ;
        RECT 306.050 93.080 306.220 93.540 ;
        RECT 307.155 93.420 307.325 93.800 ;
        RECT 308.545 93.630 308.715 94.220 ;
        RECT 309.455 94.100 309.665 94.750 ;
        RECT 309.840 94.710 311.050 95.460 ;
        RECT 306.455 93.080 307.325 93.420 ;
        RECT 307.915 93.460 308.715 93.630 ;
        RECT 307.495 92.910 307.745 93.370 ;
        RECT 307.915 93.170 308.085 93.460 ;
        RECT 308.265 92.910 308.595 93.290 ;
        RECT 308.935 92.910 309.240 94.050 ;
        RECT 309.410 93.220 309.665 94.100 ;
        RECT 309.840 94.000 310.360 94.540 ;
        RECT 310.530 94.170 311.050 94.710 ;
        RECT 309.840 92.910 311.050 94.000 ;
        RECT 162.095 92.740 311.135 92.910 ;
        RECT 162.180 91.650 163.390 92.740 ;
        RECT 163.560 91.650 165.230 92.740 ;
        RECT 165.405 92.070 165.660 92.570 ;
        RECT 165.830 92.240 166.160 92.740 ;
        RECT 165.405 91.900 166.155 92.070 ;
        RECT 162.180 90.940 162.700 91.480 ;
        RECT 162.870 91.110 163.390 91.650 ;
        RECT 163.560 90.960 164.310 91.480 ;
        RECT 164.480 91.130 165.230 91.650 ;
        RECT 165.405 91.080 165.755 91.730 ;
        RECT 162.180 90.190 163.390 90.940 ;
        RECT 163.560 90.190 165.230 90.960 ;
        RECT 165.925 90.910 166.155 91.900 ;
        RECT 165.405 90.740 166.155 90.910 ;
        RECT 165.405 90.450 165.660 90.740 ;
        RECT 165.830 90.190 166.160 90.570 ;
        RECT 166.330 90.450 166.500 92.570 ;
        RECT 166.670 91.770 166.995 92.555 ;
        RECT 167.165 92.280 167.415 92.740 ;
        RECT 167.585 92.240 167.835 92.570 ;
        RECT 168.050 92.240 168.730 92.570 ;
        RECT 167.585 92.110 167.755 92.240 ;
        RECT 167.360 91.940 167.755 92.110 ;
        RECT 166.730 90.720 167.190 91.770 ;
        RECT 167.360 90.580 167.530 91.940 ;
        RECT 167.925 91.680 168.390 92.070 ;
        RECT 167.700 90.870 168.050 91.490 ;
        RECT 168.220 91.090 168.390 91.680 ;
        RECT 168.560 91.460 168.730 92.240 ;
        RECT 168.900 92.140 169.070 92.480 ;
        RECT 169.305 92.310 169.635 92.740 ;
        RECT 169.805 92.140 169.975 92.480 ;
        RECT 170.270 92.280 170.640 92.740 ;
        RECT 168.900 91.970 169.975 92.140 ;
        RECT 170.810 92.110 170.980 92.570 ;
        RECT 171.215 92.230 172.085 92.570 ;
        RECT 172.255 92.280 172.505 92.740 ;
        RECT 170.420 91.940 170.980 92.110 ;
        RECT 170.420 91.800 170.590 91.940 ;
        RECT 169.090 91.630 170.590 91.800 ;
        RECT 171.285 91.770 171.745 92.060 ;
        RECT 168.560 91.290 170.250 91.460 ;
        RECT 168.220 90.870 168.575 91.090 ;
        RECT 168.745 90.580 168.915 91.290 ;
        RECT 169.120 90.870 169.910 91.120 ;
        RECT 170.080 91.110 170.250 91.290 ;
        RECT 170.420 90.940 170.590 91.630 ;
        RECT 166.860 90.190 167.190 90.550 ;
        RECT 167.360 90.410 167.855 90.580 ;
        RECT 168.060 90.410 168.915 90.580 ;
        RECT 169.790 90.190 170.120 90.650 ;
        RECT 170.330 90.550 170.590 90.940 ;
        RECT 170.780 91.760 171.745 91.770 ;
        RECT 171.915 91.850 172.085 92.230 ;
        RECT 172.675 92.190 172.845 92.480 ;
        RECT 173.025 92.360 173.355 92.740 ;
        RECT 172.675 92.020 173.475 92.190 ;
        RECT 170.780 91.600 171.455 91.760 ;
        RECT 171.915 91.680 173.135 91.850 ;
        RECT 170.780 90.810 170.990 91.600 ;
        RECT 171.915 91.590 172.085 91.680 ;
        RECT 171.160 90.810 171.510 91.430 ;
        RECT 171.680 91.420 172.085 91.590 ;
        RECT 171.680 90.640 171.850 91.420 ;
        RECT 172.020 90.970 172.240 91.250 ;
        RECT 172.420 91.140 172.960 91.510 ;
        RECT 173.305 91.430 173.475 92.020 ;
        RECT 173.695 91.600 174.000 92.740 ;
        RECT 174.170 91.550 174.420 92.430 ;
        RECT 174.590 91.600 174.840 92.740 ;
        RECT 175.060 91.575 175.350 92.740 ;
        RECT 175.525 91.600 175.860 92.570 ;
        RECT 176.030 91.600 176.200 92.740 ;
        RECT 176.370 92.400 178.400 92.570 ;
        RECT 173.305 91.400 174.045 91.430 ;
        RECT 172.020 90.800 172.550 90.970 ;
        RECT 170.330 90.380 170.680 90.550 ;
        RECT 170.900 90.360 171.850 90.640 ;
        RECT 172.020 90.190 172.210 90.630 ;
        RECT 172.380 90.570 172.550 90.800 ;
        RECT 172.720 90.740 172.960 91.140 ;
        RECT 173.130 91.100 174.045 91.400 ;
        RECT 173.130 90.925 173.455 91.100 ;
        RECT 173.130 90.570 173.450 90.925 ;
        RECT 174.215 90.900 174.420 91.550 ;
        RECT 172.380 90.400 173.450 90.570 ;
        RECT 173.695 90.190 174.000 90.650 ;
        RECT 174.170 90.370 174.420 90.900 ;
        RECT 174.590 90.190 174.840 90.945 ;
        RECT 175.525 90.930 175.695 91.600 ;
        RECT 176.370 91.430 176.540 92.400 ;
        RECT 175.865 91.100 176.120 91.430 ;
        RECT 176.345 91.100 176.540 91.430 ;
        RECT 176.710 92.060 177.835 92.230 ;
        RECT 175.950 90.930 176.120 91.100 ;
        RECT 176.710 90.930 176.880 92.060 ;
        RECT 175.060 90.190 175.350 90.915 ;
        RECT 175.525 90.360 175.780 90.930 ;
        RECT 175.950 90.760 176.880 90.930 ;
        RECT 177.050 91.720 178.060 91.890 ;
        RECT 177.050 90.920 177.220 91.720 ;
        RECT 177.425 91.040 177.700 91.520 ;
        RECT 177.420 90.870 177.700 91.040 ;
        RECT 176.705 90.725 176.880 90.760 ;
        RECT 175.950 90.190 176.280 90.590 ;
        RECT 176.705 90.360 177.235 90.725 ;
        RECT 177.425 90.360 177.700 90.870 ;
        RECT 177.870 90.360 178.060 91.720 ;
        RECT 178.230 91.735 178.400 92.400 ;
        RECT 178.570 91.980 178.740 92.740 ;
        RECT 178.975 91.980 179.490 92.390 ;
        RECT 178.230 91.545 178.980 91.735 ;
        RECT 179.150 91.170 179.490 91.980 ;
        RECT 179.660 91.650 183.170 92.740 ;
        RECT 178.260 91.000 179.490 91.170 ;
        RECT 178.240 90.190 178.750 90.725 ;
        RECT 178.970 90.395 179.215 91.000 ;
        RECT 179.660 90.960 181.310 91.480 ;
        RECT 181.480 91.130 183.170 91.650 ;
        RECT 183.800 91.980 184.315 92.390 ;
        RECT 184.550 91.980 184.720 92.740 ;
        RECT 184.890 92.400 186.920 92.570 ;
        RECT 183.800 91.170 184.140 91.980 ;
        RECT 184.890 91.735 185.060 92.400 ;
        RECT 185.455 92.060 186.580 92.230 ;
        RECT 184.310 91.545 185.060 91.735 ;
        RECT 185.230 91.720 186.240 91.890 ;
        RECT 183.800 91.000 185.030 91.170 ;
        RECT 179.660 90.190 183.170 90.960 ;
        RECT 184.075 90.395 184.320 91.000 ;
        RECT 184.540 90.190 185.050 90.725 ;
        RECT 185.230 90.360 185.420 91.720 ;
        RECT 185.590 90.700 185.865 91.520 ;
        RECT 186.070 90.920 186.240 91.720 ;
        RECT 186.410 90.930 186.580 92.060 ;
        RECT 186.750 91.430 186.920 92.400 ;
        RECT 187.090 91.600 187.260 92.740 ;
        RECT 187.430 91.600 187.765 92.570 ;
        RECT 186.750 91.100 186.945 91.430 ;
        RECT 187.170 91.100 187.425 91.430 ;
        RECT 187.170 90.930 187.340 91.100 ;
        RECT 187.595 90.930 187.765 91.600 ;
        RECT 186.410 90.760 187.340 90.930 ;
        RECT 186.410 90.725 186.585 90.760 ;
        RECT 185.590 90.530 185.870 90.700 ;
        RECT 185.590 90.360 185.865 90.530 ;
        RECT 186.055 90.360 186.585 90.725 ;
        RECT 187.010 90.190 187.340 90.590 ;
        RECT 187.510 90.360 187.765 90.930 ;
        RECT 188.865 91.600 189.200 92.570 ;
        RECT 189.370 91.600 189.540 92.740 ;
        RECT 189.710 92.400 191.740 92.570 ;
        RECT 188.865 90.930 189.035 91.600 ;
        RECT 189.710 91.430 189.880 92.400 ;
        RECT 189.205 91.100 189.460 91.430 ;
        RECT 189.685 91.100 189.880 91.430 ;
        RECT 190.050 92.060 191.175 92.230 ;
        RECT 189.290 90.930 189.460 91.100 ;
        RECT 190.050 90.930 190.220 92.060 ;
        RECT 188.865 90.360 189.120 90.930 ;
        RECT 189.290 90.760 190.220 90.930 ;
        RECT 190.390 91.720 191.400 91.890 ;
        RECT 190.390 90.920 190.560 91.720 ;
        RECT 190.765 91.040 191.040 91.520 ;
        RECT 190.760 90.870 191.040 91.040 ;
        RECT 190.045 90.725 190.220 90.760 ;
        RECT 189.290 90.190 189.620 90.590 ;
        RECT 190.045 90.360 190.575 90.725 ;
        RECT 190.765 90.360 191.040 90.870 ;
        RECT 191.210 90.360 191.400 91.720 ;
        RECT 191.570 91.735 191.740 92.400 ;
        RECT 191.910 91.980 192.080 92.740 ;
        RECT 192.315 91.980 192.830 92.390 ;
        RECT 191.570 91.545 192.320 91.735 ;
        RECT 192.490 91.170 192.830 91.980 ;
        RECT 191.600 91.000 192.830 91.170 ;
        RECT 193.925 91.600 194.260 92.570 ;
        RECT 194.430 91.600 194.600 92.740 ;
        RECT 194.770 92.400 196.800 92.570 ;
        RECT 191.580 90.190 192.090 90.725 ;
        RECT 192.310 90.395 192.555 91.000 ;
        RECT 193.925 90.930 194.095 91.600 ;
        RECT 194.770 91.430 194.940 92.400 ;
        RECT 194.265 91.100 194.520 91.430 ;
        RECT 194.745 91.100 194.940 91.430 ;
        RECT 195.110 92.060 196.235 92.230 ;
        RECT 194.350 90.930 194.520 91.100 ;
        RECT 195.110 90.930 195.280 92.060 ;
        RECT 193.925 90.360 194.180 90.930 ;
        RECT 194.350 90.760 195.280 90.930 ;
        RECT 195.450 91.720 196.460 91.890 ;
        RECT 195.450 90.920 195.620 91.720 ;
        RECT 195.105 90.725 195.280 90.760 ;
        RECT 194.350 90.190 194.680 90.590 ;
        RECT 195.105 90.360 195.635 90.725 ;
        RECT 195.825 90.700 196.100 91.520 ;
        RECT 195.820 90.530 196.100 90.700 ;
        RECT 195.825 90.360 196.100 90.530 ;
        RECT 196.270 90.360 196.460 91.720 ;
        RECT 196.630 91.735 196.800 92.400 ;
        RECT 196.970 91.980 197.140 92.740 ;
        RECT 197.375 91.980 197.890 92.390 ;
        RECT 196.630 91.545 197.380 91.735 ;
        RECT 197.550 91.170 197.890 91.980 ;
        RECT 198.115 91.870 198.400 92.740 ;
        RECT 198.570 92.110 198.830 92.570 ;
        RECT 199.005 92.280 199.260 92.740 ;
        RECT 199.430 92.110 199.690 92.570 ;
        RECT 198.570 91.940 199.690 92.110 ;
        RECT 199.860 91.940 200.170 92.740 ;
        RECT 198.570 91.690 198.830 91.940 ;
        RECT 200.340 91.770 200.650 92.570 ;
        RECT 196.660 91.000 197.890 91.170 ;
        RECT 198.075 91.520 198.830 91.690 ;
        RECT 199.620 91.600 200.650 91.770 ;
        RECT 198.075 91.010 198.480 91.520 ;
        RECT 199.620 91.350 199.790 91.600 ;
        RECT 198.650 91.180 199.790 91.350 ;
        RECT 196.640 90.190 197.150 90.725 ;
        RECT 197.370 90.395 197.615 91.000 ;
        RECT 198.075 90.840 199.725 91.010 ;
        RECT 199.960 90.860 200.310 91.430 ;
        RECT 198.120 90.190 198.400 90.670 ;
        RECT 198.570 90.450 198.830 90.840 ;
        RECT 199.005 90.190 199.260 90.670 ;
        RECT 199.430 90.450 199.725 90.840 ;
        RECT 200.480 90.690 200.650 91.600 ;
        RECT 200.820 91.575 201.110 92.740 ;
        RECT 201.280 91.650 202.490 92.740 ;
        RECT 201.280 90.940 201.800 91.480 ;
        RECT 201.970 91.110 202.490 91.650 ;
        RECT 202.665 91.600 203.000 92.570 ;
        RECT 203.170 91.600 203.340 92.740 ;
        RECT 203.510 92.400 205.540 92.570 ;
        RECT 199.905 90.190 200.180 90.670 ;
        RECT 200.350 90.360 200.650 90.690 ;
        RECT 200.820 90.190 201.110 90.915 ;
        RECT 201.280 90.190 202.490 90.940 ;
        RECT 202.665 90.930 202.835 91.600 ;
        RECT 203.510 91.430 203.680 92.400 ;
        RECT 203.005 91.100 203.260 91.430 ;
        RECT 203.485 91.100 203.680 91.430 ;
        RECT 203.850 92.060 204.975 92.230 ;
        RECT 203.090 90.930 203.260 91.100 ;
        RECT 203.850 90.930 204.020 92.060 ;
        RECT 202.665 90.360 202.920 90.930 ;
        RECT 203.090 90.760 204.020 90.930 ;
        RECT 204.190 91.720 205.200 91.890 ;
        RECT 204.190 90.920 204.360 91.720 ;
        RECT 204.565 91.380 204.840 91.520 ;
        RECT 204.560 91.210 204.840 91.380 ;
        RECT 203.845 90.725 204.020 90.760 ;
        RECT 203.090 90.190 203.420 90.590 ;
        RECT 203.845 90.360 204.375 90.725 ;
        RECT 204.565 90.360 204.840 91.210 ;
        RECT 205.010 90.360 205.200 91.720 ;
        RECT 205.370 91.735 205.540 92.400 ;
        RECT 205.710 91.980 205.880 92.740 ;
        RECT 206.115 91.980 206.630 92.390 ;
        RECT 205.370 91.545 206.120 91.735 ;
        RECT 206.290 91.170 206.630 91.980 ;
        RECT 205.400 91.000 206.630 91.170 ;
        RECT 206.800 91.135 207.080 92.570 ;
        RECT 207.250 91.965 207.960 92.740 ;
        RECT 208.130 91.795 208.460 92.570 ;
        RECT 207.310 91.580 208.460 91.795 ;
        RECT 205.380 90.190 205.890 90.725 ;
        RECT 206.110 90.395 206.355 91.000 ;
        RECT 206.800 90.360 207.140 91.135 ;
        RECT 207.310 91.010 207.595 91.580 ;
        RECT 207.780 91.180 208.250 91.410 ;
        RECT 208.655 91.380 208.870 92.495 ;
        RECT 209.050 92.020 209.380 92.740 ;
        RECT 209.160 91.380 209.390 91.720 ;
        RECT 209.560 91.650 212.150 92.740 ;
        RECT 208.420 91.200 208.870 91.380 ;
        RECT 208.420 91.180 208.750 91.200 ;
        RECT 209.060 91.180 209.390 91.380 ;
        RECT 207.310 90.820 208.020 91.010 ;
        RECT 207.720 90.680 208.020 90.820 ;
        RECT 208.210 90.820 209.390 91.010 ;
        RECT 208.210 90.740 208.540 90.820 ;
        RECT 207.720 90.670 208.035 90.680 ;
        RECT 207.720 90.660 208.045 90.670 ;
        RECT 207.720 90.655 208.055 90.660 ;
        RECT 207.310 90.190 207.480 90.650 ;
        RECT 207.720 90.645 208.060 90.655 ;
        RECT 207.720 90.640 208.065 90.645 ;
        RECT 207.720 90.630 208.070 90.640 ;
        RECT 207.720 90.625 208.075 90.630 ;
        RECT 207.720 90.360 208.080 90.625 ;
        RECT 208.710 90.190 208.880 90.650 ;
        RECT 209.050 90.360 209.390 90.820 ;
        RECT 209.560 90.960 210.770 91.480 ;
        RECT 210.940 91.130 212.150 91.650 ;
        RECT 209.560 90.190 212.150 90.960 ;
        RECT 212.780 90.360 213.530 92.570 ;
        RECT 214.625 92.360 214.960 92.740 ;
        RECT 214.620 90.870 214.860 92.180 ;
        RECT 215.130 91.770 215.380 92.570 ;
        RECT 215.600 92.020 215.930 92.740 ;
        RECT 216.115 91.770 216.365 92.570 ;
        RECT 216.830 91.940 217.160 92.740 ;
        RECT 217.330 92.310 217.670 92.570 ;
        RECT 215.030 91.600 217.220 91.770 ;
        RECT 215.030 90.690 215.200 91.600 ;
        RECT 216.905 91.430 217.220 91.600 ;
        RECT 214.705 90.360 215.200 90.690 ;
        RECT 215.420 90.465 215.770 91.430 ;
        RECT 215.950 90.460 216.250 91.430 ;
        RECT 216.430 90.460 216.710 91.430 ;
        RECT 216.905 91.180 217.235 91.430 ;
        RECT 216.890 90.190 217.160 90.990 ;
        RECT 217.410 90.910 217.670 92.310 ;
        RECT 217.840 91.650 219.510 92.740 ;
        RECT 217.330 90.400 217.670 90.910 ;
        RECT 217.840 90.960 218.590 91.480 ;
        RECT 218.760 91.130 219.510 91.650 ;
        RECT 219.680 92.310 220.020 92.570 ;
        RECT 217.840 90.190 219.510 90.960 ;
        RECT 219.680 90.910 219.940 92.310 ;
        RECT 220.190 91.940 220.520 92.740 ;
        RECT 220.985 91.770 221.235 92.570 ;
        RECT 221.420 92.020 221.750 92.740 ;
        RECT 221.970 91.770 222.220 92.570 ;
        RECT 222.390 92.360 222.725 92.740 ;
        RECT 220.130 91.600 222.320 91.770 ;
        RECT 220.130 91.430 220.445 91.600 ;
        RECT 220.115 91.180 220.445 91.430 ;
        RECT 219.680 90.400 220.020 90.910 ;
        RECT 220.190 90.190 220.460 90.990 ;
        RECT 220.640 90.460 220.920 91.430 ;
        RECT 221.100 90.460 221.400 91.430 ;
        RECT 221.580 90.465 221.930 91.430 ;
        RECT 222.150 90.690 222.320 91.600 ;
        RECT 222.490 90.870 222.730 92.180 ;
        RECT 222.150 90.360 222.645 90.690 ;
        RECT 223.820 90.360 224.570 92.570 ;
        RECT 224.740 91.650 226.410 92.740 ;
        RECT 224.740 90.960 225.490 91.480 ;
        RECT 225.660 91.130 226.410 91.650 ;
        RECT 226.580 91.575 226.870 92.740 ;
        RECT 227.040 91.870 227.315 92.570 ;
        RECT 227.525 92.195 227.740 92.740 ;
        RECT 227.910 92.230 228.385 92.570 ;
        RECT 228.555 92.235 229.170 92.740 ;
        RECT 228.555 92.060 228.750 92.235 ;
        RECT 224.740 90.190 226.410 90.960 ;
        RECT 226.580 90.190 226.870 90.915 ;
        RECT 227.040 90.840 227.210 91.870 ;
        RECT 227.485 91.700 228.200 91.995 ;
        RECT 228.420 91.870 228.750 92.060 ;
        RECT 228.920 91.700 229.170 92.065 ;
        RECT 227.380 91.530 229.170 91.700 ;
        RECT 227.380 91.100 227.610 91.530 ;
        RECT 227.040 90.360 227.300 90.840 ;
        RECT 227.780 90.830 228.190 91.350 ;
        RECT 227.470 90.190 227.800 90.650 ;
        RECT 227.990 90.410 228.190 90.830 ;
        RECT 228.360 90.675 228.615 91.530 ;
        RECT 229.410 91.350 229.580 92.570 ;
        RECT 229.830 92.230 230.090 92.740 ;
        RECT 230.260 92.305 235.605 92.740 ;
        RECT 228.785 91.100 229.580 91.350 ;
        RECT 229.750 91.180 230.090 92.060 ;
        RECT 229.330 91.010 229.580 91.100 ;
        RECT 228.360 90.410 229.150 90.675 ;
        RECT 229.330 90.590 229.660 91.010 ;
        RECT 229.830 90.190 230.090 91.010 ;
        RECT 231.845 90.735 232.185 91.565 ;
        RECT 233.665 91.055 234.015 92.305 ;
        RECT 235.780 91.650 237.450 92.740 ;
        RECT 238.165 92.120 238.340 92.570 ;
        RECT 238.510 92.300 238.840 92.740 ;
        RECT 239.145 92.150 239.315 92.570 ;
        RECT 239.550 92.330 240.220 92.740 ;
        RECT 240.435 92.150 240.605 92.570 ;
        RECT 240.805 92.330 241.135 92.740 ;
        RECT 238.165 91.950 238.795 92.120 ;
        RECT 235.780 90.960 236.530 91.480 ;
        RECT 236.700 91.130 237.450 91.650 ;
        RECT 238.080 91.100 238.445 91.780 ;
        RECT 238.625 91.430 238.795 91.950 ;
        RECT 239.145 91.980 241.160 92.150 ;
        RECT 238.625 91.100 238.975 91.430 ;
        RECT 230.260 90.190 235.605 90.735 ;
        RECT 235.780 90.190 237.450 90.960 ;
        RECT 238.625 90.930 238.795 91.100 ;
        RECT 238.165 90.760 238.795 90.930 ;
        RECT 238.165 90.360 238.340 90.760 ;
        RECT 239.145 90.690 239.315 91.980 ;
        RECT 238.510 90.190 238.840 90.570 ;
        RECT 239.085 90.360 239.315 90.690 ;
        RECT 239.515 90.525 239.795 91.800 ;
        RECT 240.020 91.720 240.290 91.800 ;
        RECT 239.980 91.550 240.290 91.720 ;
        RECT 240.020 90.525 240.290 91.550 ;
        RECT 240.480 90.770 240.820 91.800 ;
        RECT 240.990 91.430 241.160 91.980 ;
        RECT 241.330 91.600 241.590 92.570 ;
        RECT 241.760 92.230 242.950 92.520 ;
        RECT 241.780 91.890 242.950 92.060 ;
        RECT 243.120 91.940 243.400 92.740 ;
        RECT 241.780 91.600 242.105 91.890 ;
        RECT 242.780 91.770 242.950 91.890 ;
        RECT 240.990 91.100 241.250 91.430 ;
        RECT 241.420 90.910 241.590 91.600 ;
        RECT 242.275 91.430 242.470 91.720 ;
        RECT 242.780 91.600 243.440 91.770 ;
        RECT 243.610 91.600 243.885 92.570 ;
        RECT 244.060 92.305 249.405 92.740 ;
        RECT 243.270 91.430 243.440 91.600 ;
        RECT 241.760 91.100 242.105 91.430 ;
        RECT 242.275 91.100 243.100 91.430 ;
        RECT 243.270 91.100 243.545 91.430 ;
        RECT 243.270 90.930 243.440 91.100 ;
        RECT 240.750 90.190 241.080 90.570 ;
        RECT 241.250 90.445 241.590 90.910 ;
        RECT 241.775 90.760 243.440 90.930 ;
        RECT 243.715 90.865 243.885 91.600 ;
        RECT 241.250 90.400 241.585 90.445 ;
        RECT 241.775 90.410 242.030 90.760 ;
        RECT 242.200 90.190 242.530 90.590 ;
        RECT 242.700 90.410 242.870 90.760 ;
        RECT 243.040 90.190 243.420 90.590 ;
        RECT 243.610 90.520 243.885 90.865 ;
        RECT 245.645 90.735 245.985 91.565 ;
        RECT 247.465 91.055 247.815 92.305 ;
        RECT 249.580 91.650 252.170 92.740 ;
        RECT 249.580 90.960 250.790 91.480 ;
        RECT 250.960 91.130 252.170 91.650 ;
        RECT 252.340 91.575 252.630 92.740 ;
        RECT 252.800 92.305 258.145 92.740 ;
        RECT 244.060 90.190 249.405 90.735 ;
        RECT 249.580 90.190 252.170 90.960 ;
        RECT 252.340 90.190 252.630 90.915 ;
        RECT 254.385 90.735 254.725 91.565 ;
        RECT 256.205 91.055 256.555 92.305 ;
        RECT 258.785 91.790 259.050 92.560 ;
        RECT 259.220 92.020 259.550 92.740 ;
        RECT 259.740 92.200 260.000 92.560 ;
        RECT 260.170 92.370 260.500 92.740 ;
        RECT 260.670 92.200 260.930 92.560 ;
        RECT 259.740 91.970 260.930 92.200 ;
        RECT 261.500 91.790 261.790 92.560 ;
        RECT 262.000 92.305 267.345 92.740 ;
        RECT 267.520 92.305 272.865 92.740 ;
        RECT 252.800 90.190 258.145 90.735 ;
        RECT 258.785 90.370 259.120 91.790 ;
        RECT 259.295 91.610 261.790 91.790 ;
        RECT 259.295 90.920 259.520 91.610 ;
        RECT 259.720 91.100 260.000 91.430 ;
        RECT 260.180 91.100 260.755 91.430 ;
        RECT 260.935 91.100 261.370 91.430 ;
        RECT 261.550 91.100 261.820 91.430 ;
        RECT 259.295 90.730 261.780 90.920 ;
        RECT 263.585 90.735 263.925 91.565 ;
        RECT 265.405 91.055 265.755 92.305 ;
        RECT 269.105 90.735 269.445 91.565 ;
        RECT 270.925 91.055 271.275 92.305 ;
        RECT 273.040 91.650 276.550 92.740 ;
        RECT 273.040 90.960 274.690 91.480 ;
        RECT 274.860 91.130 276.550 91.650 ;
        RECT 276.720 91.665 276.990 92.570 ;
        RECT 277.160 91.980 277.490 92.740 ;
        RECT 277.670 91.810 277.840 92.570 ;
        RECT 259.300 90.190 260.045 90.560 ;
        RECT 260.610 90.370 260.865 90.730 ;
        RECT 261.045 90.190 261.375 90.560 ;
        RECT 261.555 90.370 261.780 90.730 ;
        RECT 262.000 90.190 267.345 90.735 ;
        RECT 267.520 90.190 272.865 90.735 ;
        RECT 273.040 90.190 276.550 90.960 ;
        RECT 276.720 90.865 276.890 91.665 ;
        RECT 277.175 91.640 277.840 91.810 ;
        RECT 277.175 91.495 277.345 91.640 ;
        RECT 278.100 91.575 278.390 92.740 ;
        RECT 278.565 91.600 278.900 92.570 ;
        RECT 279.070 91.600 279.240 92.740 ;
        RECT 279.410 92.400 281.440 92.570 ;
        RECT 277.060 91.165 277.345 91.495 ;
        RECT 277.175 90.910 277.345 91.165 ;
        RECT 277.580 91.090 277.910 91.460 ;
        RECT 278.565 90.930 278.735 91.600 ;
        RECT 279.410 91.430 279.580 92.400 ;
        RECT 278.905 91.100 279.160 91.430 ;
        RECT 279.385 91.100 279.580 91.430 ;
        RECT 279.750 92.060 280.875 92.230 ;
        RECT 278.990 90.930 279.160 91.100 ;
        RECT 279.750 90.930 279.920 92.060 ;
        RECT 276.720 90.360 276.980 90.865 ;
        RECT 277.175 90.740 277.840 90.910 ;
        RECT 277.160 90.190 277.490 90.570 ;
        RECT 277.670 90.360 277.840 90.740 ;
        RECT 278.100 90.190 278.390 90.915 ;
        RECT 278.565 90.360 278.820 90.930 ;
        RECT 278.990 90.760 279.920 90.930 ;
        RECT 280.090 91.720 281.100 91.890 ;
        RECT 280.090 90.920 280.260 91.720 ;
        RECT 280.465 91.040 280.740 91.520 ;
        RECT 280.460 90.870 280.740 91.040 ;
        RECT 279.745 90.725 279.920 90.760 ;
        RECT 278.990 90.190 279.320 90.590 ;
        RECT 279.745 90.360 280.275 90.725 ;
        RECT 280.465 90.360 280.740 90.870 ;
        RECT 280.910 90.360 281.100 91.720 ;
        RECT 281.270 91.735 281.440 92.400 ;
        RECT 281.610 91.980 281.780 92.740 ;
        RECT 282.015 91.980 282.530 92.390 ;
        RECT 281.270 91.545 282.020 91.735 ;
        RECT 282.190 91.170 282.530 91.980 ;
        RECT 282.790 91.810 282.960 92.570 ;
        RECT 283.140 91.980 283.470 92.740 ;
        RECT 282.790 91.640 283.455 91.810 ;
        RECT 283.640 91.665 283.910 92.570 ;
        RECT 284.080 92.305 289.425 92.740 ;
        RECT 283.285 91.495 283.455 91.640 ;
        RECT 281.300 91.000 282.530 91.170 ;
        RECT 282.720 91.090 283.050 91.460 ;
        RECT 283.285 91.165 283.570 91.495 ;
        RECT 281.280 90.190 281.790 90.725 ;
        RECT 282.010 90.395 282.255 91.000 ;
        RECT 283.285 90.910 283.455 91.165 ;
        RECT 282.790 90.740 283.455 90.910 ;
        RECT 283.740 90.865 283.910 91.665 ;
        RECT 282.790 90.360 282.960 90.740 ;
        RECT 283.140 90.190 283.470 90.570 ;
        RECT 283.650 90.360 283.910 90.865 ;
        RECT 285.665 90.735 286.005 91.565 ;
        RECT 287.485 91.055 287.835 92.305 ;
        RECT 290.065 91.600 290.400 92.570 ;
        RECT 290.570 91.600 290.740 92.740 ;
        RECT 290.910 92.400 292.940 92.570 ;
        RECT 290.065 90.930 290.235 91.600 ;
        RECT 290.910 91.430 291.080 92.400 ;
        RECT 290.405 91.100 290.660 91.430 ;
        RECT 290.885 91.100 291.080 91.430 ;
        RECT 291.250 92.060 292.375 92.230 ;
        RECT 290.490 90.930 290.660 91.100 ;
        RECT 291.250 90.930 291.420 92.060 ;
        RECT 284.080 90.190 289.425 90.735 ;
        RECT 290.065 90.360 290.320 90.930 ;
        RECT 290.490 90.760 291.420 90.930 ;
        RECT 291.590 91.720 292.600 91.890 ;
        RECT 291.590 90.920 291.760 91.720 ;
        RECT 291.965 91.040 292.240 91.520 ;
        RECT 291.960 90.870 292.240 91.040 ;
        RECT 291.245 90.725 291.420 90.760 ;
        RECT 290.490 90.190 290.820 90.590 ;
        RECT 291.245 90.360 291.775 90.725 ;
        RECT 291.965 90.360 292.240 90.870 ;
        RECT 292.410 90.360 292.600 91.720 ;
        RECT 292.770 91.735 292.940 92.400 ;
        RECT 293.110 91.980 293.280 92.740 ;
        RECT 293.515 91.980 294.030 92.390 ;
        RECT 292.770 91.545 293.520 91.735 ;
        RECT 293.690 91.170 294.030 91.980 ;
        RECT 294.200 91.650 295.870 92.740 ;
        RECT 292.800 91.000 294.030 91.170 ;
        RECT 292.780 90.190 293.290 90.725 ;
        RECT 293.510 90.395 293.755 91.000 ;
        RECT 294.200 90.960 294.950 91.480 ;
        RECT 295.120 91.130 295.870 91.650 ;
        RECT 296.040 91.980 296.555 92.390 ;
        RECT 296.790 91.980 296.960 92.740 ;
        RECT 297.130 92.400 299.160 92.570 ;
        RECT 296.040 91.170 296.380 91.980 ;
        RECT 297.130 91.735 297.300 92.400 ;
        RECT 297.695 92.060 298.820 92.230 ;
        RECT 296.550 91.545 297.300 91.735 ;
        RECT 297.470 91.720 298.480 91.890 ;
        RECT 296.040 91.000 297.270 91.170 ;
        RECT 294.200 90.190 295.870 90.960 ;
        RECT 296.315 90.395 296.560 91.000 ;
        RECT 296.780 90.190 297.290 90.725 ;
        RECT 297.470 90.360 297.660 91.720 ;
        RECT 297.830 90.700 298.105 91.520 ;
        RECT 298.310 90.920 298.480 91.720 ;
        RECT 298.650 90.930 298.820 92.060 ;
        RECT 298.990 91.430 299.160 92.400 ;
        RECT 299.330 91.600 299.500 92.740 ;
        RECT 299.670 91.600 300.005 92.570 ;
        RECT 300.270 91.810 300.440 92.570 ;
        RECT 300.620 91.980 300.950 92.740 ;
        RECT 300.270 91.640 300.935 91.810 ;
        RECT 301.120 91.665 301.390 92.570 ;
        RECT 298.990 91.100 299.185 91.430 ;
        RECT 299.410 91.100 299.665 91.430 ;
        RECT 299.410 90.930 299.580 91.100 ;
        RECT 299.835 90.930 300.005 91.600 ;
        RECT 300.765 91.495 300.935 91.640 ;
        RECT 300.200 91.090 300.530 91.460 ;
        RECT 300.765 91.165 301.050 91.495 ;
        RECT 298.650 90.760 299.580 90.930 ;
        RECT 298.650 90.725 298.825 90.760 ;
        RECT 297.830 90.530 298.110 90.700 ;
        RECT 297.830 90.360 298.105 90.530 ;
        RECT 298.295 90.360 298.825 90.725 ;
        RECT 299.250 90.190 299.580 90.590 ;
        RECT 299.750 90.360 300.005 90.930 ;
        RECT 300.765 90.910 300.935 91.165 ;
        RECT 300.270 90.740 300.935 90.910 ;
        RECT 301.220 90.865 301.390 91.665 ;
        RECT 301.560 91.650 303.230 92.740 ;
        RECT 300.270 90.360 300.440 90.740 ;
        RECT 300.620 90.190 300.950 90.570 ;
        RECT 301.130 90.360 301.390 90.865 ;
        RECT 301.560 90.960 302.310 91.480 ;
        RECT 302.480 91.130 303.230 91.650 ;
        RECT 303.860 91.575 304.150 92.740 ;
        RECT 304.320 92.305 309.665 92.740 ;
        RECT 301.560 90.190 303.230 90.960 ;
        RECT 303.860 90.190 304.150 90.915 ;
        RECT 305.905 90.735 306.245 91.565 ;
        RECT 307.725 91.055 308.075 92.305 ;
        RECT 309.840 91.650 311.050 92.740 ;
        RECT 309.840 91.110 310.360 91.650 ;
        RECT 310.530 90.940 311.050 91.480 ;
        RECT 304.320 90.190 309.665 90.735 ;
        RECT 309.840 90.190 311.050 90.940 ;
        RECT 162.095 90.020 311.135 90.190 ;
        RECT 162.180 89.270 163.390 90.020 ;
        RECT 163.560 89.270 164.770 90.020 ;
        RECT 165.030 89.470 165.200 89.850 ;
        RECT 165.380 89.640 165.710 90.020 ;
        RECT 165.030 89.300 165.695 89.470 ;
        RECT 165.890 89.345 166.150 89.850 ;
        RECT 162.180 88.730 162.700 89.270 ;
        RECT 162.870 88.560 163.390 89.100 ;
        RECT 163.560 88.730 164.080 89.270 ;
        RECT 164.250 88.560 164.770 89.100 ;
        RECT 164.960 88.750 165.290 89.120 ;
        RECT 165.525 89.045 165.695 89.300 ;
        RECT 165.525 88.715 165.810 89.045 ;
        RECT 165.525 88.570 165.695 88.715 ;
        RECT 162.180 87.470 163.390 88.560 ;
        RECT 163.560 87.470 164.770 88.560 ;
        RECT 165.030 88.400 165.695 88.570 ;
        RECT 165.980 88.545 166.150 89.345 ;
        RECT 166.325 89.470 166.580 89.760 ;
        RECT 166.750 89.640 167.080 90.020 ;
        RECT 166.325 89.300 167.075 89.470 ;
        RECT 165.030 87.640 165.200 88.400 ;
        RECT 165.380 87.470 165.710 88.230 ;
        RECT 165.880 87.640 166.150 88.545 ;
        RECT 166.325 88.480 166.675 89.130 ;
        RECT 166.845 88.310 167.075 89.300 ;
        RECT 166.325 88.140 167.075 88.310 ;
        RECT 166.325 87.640 166.580 88.140 ;
        RECT 166.750 87.470 167.080 87.970 ;
        RECT 167.250 87.640 167.420 89.760 ;
        RECT 167.780 89.660 168.110 90.020 ;
        RECT 168.280 89.630 168.775 89.800 ;
        RECT 168.980 89.630 169.835 89.800 ;
        RECT 167.650 88.440 168.110 89.490 ;
        RECT 167.590 87.655 167.915 88.440 ;
        RECT 168.280 88.270 168.450 89.630 ;
        RECT 168.620 88.720 168.970 89.340 ;
        RECT 169.140 89.120 169.495 89.340 ;
        RECT 169.140 88.530 169.310 89.120 ;
        RECT 169.665 88.920 169.835 89.630 ;
        RECT 170.710 89.560 171.040 90.020 ;
        RECT 171.250 89.660 171.600 89.830 ;
        RECT 170.040 89.090 170.830 89.340 ;
        RECT 171.250 89.270 171.510 89.660 ;
        RECT 171.820 89.570 172.770 89.850 ;
        RECT 172.940 89.580 173.130 90.020 ;
        RECT 173.300 89.640 174.370 89.810 ;
        RECT 171.000 88.920 171.170 89.100 ;
        RECT 168.280 88.100 168.675 88.270 ;
        RECT 168.845 88.140 169.310 88.530 ;
        RECT 169.480 88.750 171.170 88.920 ;
        RECT 168.505 87.970 168.675 88.100 ;
        RECT 169.480 87.970 169.650 88.750 ;
        RECT 171.340 88.580 171.510 89.270 ;
        RECT 170.010 88.410 171.510 88.580 ;
        RECT 171.700 88.610 171.910 89.400 ;
        RECT 172.080 88.780 172.430 89.400 ;
        RECT 172.600 88.790 172.770 89.570 ;
        RECT 173.300 89.410 173.470 89.640 ;
        RECT 172.940 89.240 173.470 89.410 ;
        RECT 172.940 88.960 173.160 89.240 ;
        RECT 173.640 89.070 173.880 89.470 ;
        RECT 172.600 88.620 173.005 88.790 ;
        RECT 173.340 88.700 173.880 89.070 ;
        RECT 174.050 89.285 174.370 89.640 ;
        RECT 174.615 89.560 174.920 90.020 ;
        RECT 175.090 89.310 175.340 89.840 ;
        RECT 174.050 89.110 174.375 89.285 ;
        RECT 174.050 88.810 174.965 89.110 ;
        RECT 174.225 88.780 174.965 88.810 ;
        RECT 171.700 88.450 172.375 88.610 ;
        RECT 172.835 88.530 173.005 88.620 ;
        RECT 171.700 88.440 172.665 88.450 ;
        RECT 171.340 88.270 171.510 88.410 ;
        RECT 168.085 87.470 168.335 87.930 ;
        RECT 168.505 87.640 168.755 87.970 ;
        RECT 168.970 87.640 169.650 87.970 ;
        RECT 169.820 88.070 170.895 88.240 ;
        RECT 171.340 88.100 171.900 88.270 ;
        RECT 172.205 88.150 172.665 88.440 ;
        RECT 172.835 88.360 174.055 88.530 ;
        RECT 169.820 87.730 169.990 88.070 ;
        RECT 170.225 87.470 170.555 87.900 ;
        RECT 170.725 87.730 170.895 88.070 ;
        RECT 171.190 87.470 171.560 87.930 ;
        RECT 171.730 87.640 171.900 88.100 ;
        RECT 172.835 87.980 173.005 88.360 ;
        RECT 174.225 88.190 174.395 88.780 ;
        RECT 175.135 88.660 175.340 89.310 ;
        RECT 175.510 89.265 175.760 90.020 ;
        RECT 175.985 89.470 176.240 89.760 ;
        RECT 176.410 89.640 176.740 90.020 ;
        RECT 175.985 89.300 176.735 89.470 ;
        RECT 172.135 87.640 173.005 87.980 ;
        RECT 173.595 88.020 174.395 88.190 ;
        RECT 173.175 87.470 173.425 87.930 ;
        RECT 173.595 87.730 173.765 88.020 ;
        RECT 173.945 87.470 174.275 87.850 ;
        RECT 174.615 87.470 174.920 88.610 ;
        RECT 175.090 87.780 175.340 88.660 ;
        RECT 175.510 87.470 175.760 88.610 ;
        RECT 175.985 88.480 176.335 89.130 ;
        RECT 176.505 88.310 176.735 89.300 ;
        RECT 175.985 88.140 176.735 88.310 ;
        RECT 175.985 87.640 176.240 88.140 ;
        RECT 176.410 87.470 176.740 87.970 ;
        RECT 176.910 87.640 177.080 89.760 ;
        RECT 177.440 89.660 177.770 90.020 ;
        RECT 177.940 89.630 178.435 89.800 ;
        RECT 178.640 89.630 179.495 89.800 ;
        RECT 177.310 88.440 177.770 89.490 ;
        RECT 177.250 87.655 177.575 88.440 ;
        RECT 177.940 88.270 178.110 89.630 ;
        RECT 178.280 88.720 178.630 89.340 ;
        RECT 178.800 89.120 179.155 89.340 ;
        RECT 178.800 88.530 178.970 89.120 ;
        RECT 179.325 88.920 179.495 89.630 ;
        RECT 180.370 89.560 180.700 90.020 ;
        RECT 180.910 89.660 181.260 89.830 ;
        RECT 179.700 89.090 180.490 89.340 ;
        RECT 180.910 89.270 181.170 89.660 ;
        RECT 181.480 89.570 182.430 89.850 ;
        RECT 182.600 89.580 182.790 90.020 ;
        RECT 182.960 89.640 184.030 89.810 ;
        RECT 180.660 88.920 180.830 89.100 ;
        RECT 177.940 88.100 178.335 88.270 ;
        RECT 178.505 88.140 178.970 88.530 ;
        RECT 179.140 88.750 180.830 88.920 ;
        RECT 178.165 87.970 178.335 88.100 ;
        RECT 179.140 87.970 179.310 88.750 ;
        RECT 181.000 88.580 181.170 89.270 ;
        RECT 179.670 88.410 181.170 88.580 ;
        RECT 181.360 88.610 181.570 89.400 ;
        RECT 181.740 88.780 182.090 89.400 ;
        RECT 182.260 88.790 182.430 89.570 ;
        RECT 182.960 89.410 183.130 89.640 ;
        RECT 182.600 89.240 183.130 89.410 ;
        RECT 182.600 88.960 182.820 89.240 ;
        RECT 183.300 89.070 183.540 89.470 ;
        RECT 182.260 88.620 182.665 88.790 ;
        RECT 183.000 88.700 183.540 89.070 ;
        RECT 183.710 89.285 184.030 89.640 ;
        RECT 184.275 89.560 184.580 90.020 ;
        RECT 184.750 89.310 185.000 89.840 ;
        RECT 183.710 89.110 184.035 89.285 ;
        RECT 183.710 88.810 184.625 89.110 ;
        RECT 183.885 88.780 184.625 88.810 ;
        RECT 181.360 88.450 182.035 88.610 ;
        RECT 182.495 88.530 182.665 88.620 ;
        RECT 181.360 88.440 182.325 88.450 ;
        RECT 181.000 88.270 181.170 88.410 ;
        RECT 177.745 87.470 177.995 87.930 ;
        RECT 178.165 87.640 178.415 87.970 ;
        RECT 178.630 87.640 179.310 87.970 ;
        RECT 179.480 88.070 180.555 88.240 ;
        RECT 181.000 88.100 181.560 88.270 ;
        RECT 181.865 88.150 182.325 88.440 ;
        RECT 182.495 88.360 183.715 88.530 ;
        RECT 179.480 87.730 179.650 88.070 ;
        RECT 179.885 87.470 180.215 87.900 ;
        RECT 180.385 87.730 180.555 88.070 ;
        RECT 180.850 87.470 181.220 87.930 ;
        RECT 181.390 87.640 181.560 88.100 ;
        RECT 182.495 87.980 182.665 88.360 ;
        RECT 183.885 88.190 184.055 88.780 ;
        RECT 184.795 88.660 185.000 89.310 ;
        RECT 185.170 89.265 185.420 90.020 ;
        RECT 186.560 89.345 186.820 89.850 ;
        RECT 187.000 89.640 187.330 90.020 ;
        RECT 187.510 89.470 187.680 89.850 ;
        RECT 181.795 87.640 182.665 87.980 ;
        RECT 183.255 88.020 184.055 88.190 ;
        RECT 182.835 87.470 183.085 87.930 ;
        RECT 183.255 87.730 183.425 88.020 ;
        RECT 183.605 87.470 183.935 87.850 ;
        RECT 184.275 87.470 184.580 88.610 ;
        RECT 184.750 87.780 185.000 88.660 ;
        RECT 185.170 87.470 185.420 88.610 ;
        RECT 186.560 88.545 186.730 89.345 ;
        RECT 187.015 89.300 187.680 89.470 ;
        RECT 187.015 89.045 187.185 89.300 ;
        RECT 187.940 89.295 188.230 90.020 ;
        RECT 188.400 89.345 188.660 89.850 ;
        RECT 188.840 89.640 189.170 90.020 ;
        RECT 189.350 89.470 189.520 89.850 ;
        RECT 186.900 88.715 187.185 89.045 ;
        RECT 187.420 88.750 187.750 89.120 ;
        RECT 187.015 88.570 187.185 88.715 ;
        RECT 186.560 87.640 186.830 88.545 ;
        RECT 187.015 88.400 187.680 88.570 ;
        RECT 187.000 87.470 187.330 88.230 ;
        RECT 187.510 87.640 187.680 88.400 ;
        RECT 187.940 87.470 188.230 88.635 ;
        RECT 188.400 88.545 188.570 89.345 ;
        RECT 188.855 89.300 189.520 89.470 ;
        RECT 189.785 89.470 190.040 89.760 ;
        RECT 190.210 89.640 190.540 90.020 ;
        RECT 189.785 89.300 190.535 89.470 ;
        RECT 188.855 89.045 189.025 89.300 ;
        RECT 188.740 88.715 189.025 89.045 ;
        RECT 189.260 88.750 189.590 89.120 ;
        RECT 188.855 88.570 189.025 88.715 ;
        RECT 188.400 87.640 188.670 88.545 ;
        RECT 188.855 88.400 189.520 88.570 ;
        RECT 189.785 88.480 190.135 89.130 ;
        RECT 188.840 87.470 189.170 88.230 ;
        RECT 189.350 87.640 189.520 88.400 ;
        RECT 190.305 88.310 190.535 89.300 ;
        RECT 189.785 88.140 190.535 88.310 ;
        RECT 189.785 87.640 190.040 88.140 ;
        RECT 190.210 87.470 190.540 87.970 ;
        RECT 190.710 87.640 190.880 89.760 ;
        RECT 191.240 89.660 191.570 90.020 ;
        RECT 191.740 89.630 192.235 89.800 ;
        RECT 192.440 89.630 193.295 89.800 ;
        RECT 191.110 88.440 191.570 89.490 ;
        RECT 191.050 87.655 191.375 88.440 ;
        RECT 191.740 88.270 191.910 89.630 ;
        RECT 192.080 88.720 192.430 89.340 ;
        RECT 192.600 89.120 192.955 89.340 ;
        RECT 192.600 88.530 192.770 89.120 ;
        RECT 193.125 88.920 193.295 89.630 ;
        RECT 194.170 89.560 194.500 90.020 ;
        RECT 194.710 89.660 195.060 89.830 ;
        RECT 193.500 89.090 194.290 89.340 ;
        RECT 194.710 89.270 194.970 89.660 ;
        RECT 195.280 89.570 196.230 89.850 ;
        RECT 196.400 89.580 196.590 90.020 ;
        RECT 196.760 89.640 197.830 89.810 ;
        RECT 194.460 88.920 194.630 89.100 ;
        RECT 191.740 88.100 192.135 88.270 ;
        RECT 192.305 88.140 192.770 88.530 ;
        RECT 192.940 88.750 194.630 88.920 ;
        RECT 191.965 87.970 192.135 88.100 ;
        RECT 192.940 87.970 193.110 88.750 ;
        RECT 194.800 88.580 194.970 89.270 ;
        RECT 193.470 88.410 194.970 88.580 ;
        RECT 195.160 88.610 195.370 89.400 ;
        RECT 195.540 88.780 195.890 89.400 ;
        RECT 196.060 88.790 196.230 89.570 ;
        RECT 196.760 89.410 196.930 89.640 ;
        RECT 196.400 89.240 196.930 89.410 ;
        RECT 196.400 88.960 196.620 89.240 ;
        RECT 197.100 89.070 197.340 89.470 ;
        RECT 196.060 88.620 196.465 88.790 ;
        RECT 196.800 88.700 197.340 89.070 ;
        RECT 197.510 89.285 197.830 89.640 ;
        RECT 198.075 89.560 198.380 90.020 ;
        RECT 198.550 89.310 198.805 89.840 ;
        RECT 197.510 89.110 197.835 89.285 ;
        RECT 197.510 88.810 198.425 89.110 ;
        RECT 197.685 88.780 198.425 88.810 ;
        RECT 195.160 88.450 195.835 88.610 ;
        RECT 196.295 88.530 196.465 88.620 ;
        RECT 195.160 88.440 196.125 88.450 ;
        RECT 194.800 88.270 194.970 88.410 ;
        RECT 191.545 87.470 191.795 87.930 ;
        RECT 191.965 87.640 192.215 87.970 ;
        RECT 192.430 87.640 193.110 87.970 ;
        RECT 193.280 88.070 194.355 88.240 ;
        RECT 194.800 88.100 195.360 88.270 ;
        RECT 195.665 88.150 196.125 88.440 ;
        RECT 196.295 88.360 197.515 88.530 ;
        RECT 193.280 87.730 193.450 88.070 ;
        RECT 193.685 87.470 194.015 87.900 ;
        RECT 194.185 87.730 194.355 88.070 ;
        RECT 194.650 87.470 195.020 87.930 ;
        RECT 195.190 87.640 195.360 88.100 ;
        RECT 196.295 87.980 196.465 88.360 ;
        RECT 197.685 88.190 197.855 88.780 ;
        RECT 198.595 88.660 198.805 89.310 ;
        RECT 199.990 89.470 200.160 89.850 ;
        RECT 200.340 89.640 200.670 90.020 ;
        RECT 199.990 89.300 200.655 89.470 ;
        RECT 200.850 89.345 201.110 89.850 ;
        RECT 199.920 88.750 200.250 89.120 ;
        RECT 200.485 89.045 200.655 89.300 ;
        RECT 195.595 87.640 196.465 87.980 ;
        RECT 197.055 88.020 197.855 88.190 ;
        RECT 196.635 87.470 196.885 87.930 ;
        RECT 197.055 87.730 197.225 88.020 ;
        RECT 197.405 87.470 197.735 87.850 ;
        RECT 198.075 87.470 198.380 88.610 ;
        RECT 198.550 87.780 198.805 88.660 ;
        RECT 200.485 88.715 200.770 89.045 ;
        RECT 200.485 88.570 200.655 88.715 ;
        RECT 199.990 88.400 200.655 88.570 ;
        RECT 200.940 88.545 201.110 89.345 ;
        RECT 201.285 89.470 201.540 89.760 ;
        RECT 201.710 89.640 202.040 90.020 ;
        RECT 201.285 89.300 202.035 89.470 ;
        RECT 199.990 87.640 200.160 88.400 ;
        RECT 200.340 87.470 200.670 88.230 ;
        RECT 200.840 87.640 201.110 88.545 ;
        RECT 201.285 88.480 201.635 89.130 ;
        RECT 201.805 88.310 202.035 89.300 ;
        RECT 201.285 88.140 202.035 88.310 ;
        RECT 201.285 87.640 201.540 88.140 ;
        RECT 201.710 87.470 202.040 87.970 ;
        RECT 202.210 87.640 202.380 89.760 ;
        RECT 202.740 89.660 203.070 90.020 ;
        RECT 203.240 89.630 203.735 89.800 ;
        RECT 203.940 89.630 204.795 89.800 ;
        RECT 202.610 88.440 203.070 89.490 ;
        RECT 202.550 87.655 202.875 88.440 ;
        RECT 203.240 88.270 203.410 89.630 ;
        RECT 203.580 88.720 203.930 89.340 ;
        RECT 204.100 89.120 204.455 89.340 ;
        RECT 204.100 88.530 204.270 89.120 ;
        RECT 204.625 88.920 204.795 89.630 ;
        RECT 205.670 89.560 206.000 90.020 ;
        RECT 206.210 89.660 206.560 89.830 ;
        RECT 205.000 89.090 205.790 89.340 ;
        RECT 206.210 89.270 206.470 89.660 ;
        RECT 206.780 89.570 207.730 89.850 ;
        RECT 207.900 89.580 208.090 90.020 ;
        RECT 208.260 89.640 209.330 89.810 ;
        RECT 205.960 88.920 206.130 89.100 ;
        RECT 203.240 88.100 203.635 88.270 ;
        RECT 203.805 88.140 204.270 88.530 ;
        RECT 204.440 88.750 206.130 88.920 ;
        RECT 203.465 87.970 203.635 88.100 ;
        RECT 204.440 87.970 204.610 88.750 ;
        RECT 206.300 88.580 206.470 89.270 ;
        RECT 204.970 88.410 206.470 88.580 ;
        RECT 206.660 88.610 206.870 89.400 ;
        RECT 207.040 88.780 207.390 89.400 ;
        RECT 207.560 88.790 207.730 89.570 ;
        RECT 208.260 89.410 208.430 89.640 ;
        RECT 207.900 89.240 208.430 89.410 ;
        RECT 207.900 88.960 208.120 89.240 ;
        RECT 208.600 89.070 208.840 89.470 ;
        RECT 207.560 88.620 207.965 88.790 ;
        RECT 208.300 88.700 208.840 89.070 ;
        RECT 209.010 89.285 209.330 89.640 ;
        RECT 209.575 89.560 209.880 90.020 ;
        RECT 210.050 89.310 210.300 89.840 ;
        RECT 209.010 89.110 209.335 89.285 ;
        RECT 209.010 88.810 209.925 89.110 ;
        RECT 209.185 88.780 209.925 88.810 ;
        RECT 206.660 88.450 207.335 88.610 ;
        RECT 207.795 88.530 207.965 88.620 ;
        RECT 206.660 88.440 207.625 88.450 ;
        RECT 206.300 88.270 206.470 88.410 ;
        RECT 203.045 87.470 203.295 87.930 ;
        RECT 203.465 87.640 203.715 87.970 ;
        RECT 203.930 87.640 204.610 87.970 ;
        RECT 204.780 88.070 205.855 88.240 ;
        RECT 206.300 88.100 206.860 88.270 ;
        RECT 207.165 88.150 207.625 88.440 ;
        RECT 207.795 88.360 209.015 88.530 ;
        RECT 204.780 87.730 204.950 88.070 ;
        RECT 205.185 87.470 205.515 87.900 ;
        RECT 205.685 87.730 205.855 88.070 ;
        RECT 206.150 87.470 206.520 87.930 ;
        RECT 206.690 87.640 206.860 88.100 ;
        RECT 207.795 87.980 207.965 88.360 ;
        RECT 209.185 88.190 209.355 88.780 ;
        RECT 210.095 88.660 210.300 89.310 ;
        RECT 210.470 89.265 210.720 90.020 ;
        RECT 211.030 89.470 211.200 89.850 ;
        RECT 211.415 89.640 211.745 90.020 ;
        RECT 211.030 89.300 211.745 89.470 ;
        RECT 210.940 88.750 211.295 89.120 ;
        RECT 211.575 89.110 211.745 89.300 ;
        RECT 211.915 89.275 212.170 89.850 ;
        RECT 211.575 88.780 211.830 89.110 ;
        RECT 207.095 87.640 207.965 87.980 ;
        RECT 208.555 88.020 209.355 88.190 ;
        RECT 208.135 87.470 208.385 87.930 ;
        RECT 208.555 87.730 208.725 88.020 ;
        RECT 208.905 87.470 209.235 87.850 ;
        RECT 209.575 87.470 209.880 88.610 ;
        RECT 210.050 87.780 210.300 88.660 ;
        RECT 210.470 87.470 210.720 88.610 ;
        RECT 211.575 88.570 211.745 88.780 ;
        RECT 211.030 88.400 211.745 88.570 ;
        RECT 212.000 88.545 212.170 89.275 ;
        RECT 212.345 89.180 212.605 90.020 ;
        RECT 213.700 89.295 213.990 90.020 ;
        RECT 214.160 89.250 217.670 90.020 ;
        RECT 218.860 89.345 219.100 90.020 ;
        RECT 219.275 89.260 219.830 89.820 ;
        RECT 220.010 89.450 220.215 89.845 ;
        RECT 220.385 89.620 220.730 90.020 ;
        RECT 220.900 89.455 221.230 89.845 ;
        RECT 221.505 89.635 222.180 90.020 ;
        RECT 220.900 89.450 222.120 89.455 ;
        RECT 220.010 89.280 222.120 89.450 ;
        RECT 214.160 88.730 215.810 89.250 ;
        RECT 219.525 89.110 219.830 89.260 ;
        RECT 211.030 87.640 211.200 88.400 ;
        RECT 211.415 87.470 211.745 88.230 ;
        RECT 211.915 87.640 212.170 88.545 ;
        RECT 212.345 87.470 212.605 88.620 ;
        RECT 213.700 87.470 213.990 88.635 ;
        RECT 215.980 88.560 217.670 89.080 ;
        RECT 218.805 88.815 219.305 89.080 ;
        RECT 219.525 88.780 219.910 89.110 ;
        RECT 214.160 87.470 217.670 88.560 ;
        RECT 218.825 88.440 219.955 88.610 ;
        RECT 218.825 87.645 219.095 88.440 ;
        RECT 219.275 87.470 219.490 88.270 ;
        RECT 219.670 87.645 219.955 88.440 ;
        RECT 220.135 87.640 220.415 89.110 ;
        RECT 220.595 87.640 220.925 89.055 ;
        RECT 221.095 88.815 221.525 89.055 ;
        RECT 221.095 87.640 221.300 88.815 ;
        RECT 221.900 88.640 222.120 89.280 ;
        RECT 221.470 88.460 222.120 88.640 ;
        RECT 222.350 88.485 222.680 89.850 ;
        RECT 221.470 87.645 221.680 88.460 ;
        RECT 221.920 87.470 222.250 88.290 ;
        RECT 222.425 87.645 222.680 88.485 ;
        RECT 222.900 87.640 223.160 89.850 ;
        RECT 223.330 89.640 223.660 90.020 ;
        RECT 223.870 89.110 224.065 89.685 ;
        RECT 224.335 89.110 224.520 89.690 ;
        RECT 223.330 88.190 223.500 89.110 ;
        RECT 223.810 88.780 224.065 89.110 ;
        RECT 224.290 88.780 224.520 89.110 ;
        RECT 224.770 89.680 226.250 89.850 ;
        RECT 224.770 88.780 224.940 89.680 ;
        RECT 225.110 89.180 225.660 89.510 ;
        RECT 225.850 89.350 226.250 89.680 ;
        RECT 226.430 89.640 226.760 90.020 ;
        RECT 227.070 89.520 227.330 89.850 ;
        RECT 223.870 88.470 224.065 88.780 ;
        RECT 224.335 88.470 224.520 88.780 ;
        RECT 225.110 88.190 225.280 89.180 ;
        RECT 225.850 88.870 226.020 89.350 ;
        RECT 226.600 89.160 226.810 89.340 ;
        RECT 226.190 88.990 226.810 89.160 ;
        RECT 223.330 88.020 225.280 88.190 ;
        RECT 225.450 88.700 226.020 88.870 ;
        RECT 227.160 88.820 227.330 89.520 ;
        RECT 227.500 89.475 232.845 90.020 ;
        RECT 225.450 88.190 225.620 88.700 ;
        RECT 226.200 88.650 227.330 88.820 ;
        RECT 226.200 88.530 226.370 88.650 ;
        RECT 225.790 88.360 226.370 88.530 ;
        RECT 225.450 88.020 226.190 88.190 ;
        RECT 226.640 88.150 226.990 88.480 ;
        RECT 223.330 87.470 223.660 87.850 ;
        RECT 224.085 87.640 224.255 88.020 ;
        RECT 224.515 87.470 224.845 87.850 ;
        RECT 225.040 87.640 225.210 88.020 ;
        RECT 225.420 87.470 225.750 87.850 ;
        RECT 226.000 87.640 226.190 88.020 ;
        RECT 227.160 87.970 227.330 88.650 ;
        RECT 229.085 88.645 229.425 89.475 ;
        RECT 233.020 89.250 235.610 90.020 ;
        RECT 236.290 89.480 236.515 89.840 ;
        RECT 236.695 89.650 237.025 90.020 ;
        RECT 237.205 89.480 237.460 89.840 ;
        RECT 238.025 89.650 238.770 90.020 ;
        RECT 236.290 89.290 238.775 89.480 ;
        RECT 226.430 87.470 226.760 87.850 ;
        RECT 227.070 87.640 227.330 87.970 ;
        RECT 230.905 87.905 231.255 89.155 ;
        RECT 233.020 88.730 234.230 89.250 ;
        RECT 234.400 88.560 235.610 89.080 ;
        RECT 236.250 88.780 236.520 89.110 ;
        RECT 236.700 88.780 237.135 89.110 ;
        RECT 237.315 88.780 237.890 89.110 ;
        RECT 238.070 88.780 238.350 89.110 ;
        RECT 238.550 88.600 238.775 89.290 ;
        RECT 227.500 87.470 232.845 87.905 ;
        RECT 233.020 87.470 235.610 88.560 ;
        RECT 236.280 88.420 238.775 88.600 ;
        RECT 238.950 88.420 239.285 89.840 ;
        RECT 239.460 89.295 239.750 90.020 ;
        RECT 240.080 89.460 240.410 89.850 ;
        RECT 240.580 89.630 241.765 89.800 ;
        RECT 242.025 89.550 242.195 90.020 ;
        RECT 240.080 89.280 240.590 89.460 ;
        RECT 239.920 88.820 240.250 89.110 ;
        RECT 240.420 88.650 240.590 89.280 ;
        RECT 240.995 89.370 241.380 89.460 ;
        RECT 242.365 89.370 242.695 89.835 ;
        RECT 240.995 89.200 242.695 89.370 ;
        RECT 242.865 89.200 243.035 90.020 ;
        RECT 243.205 89.200 243.890 89.840 ;
        RECT 244.060 89.475 249.405 90.020 ;
        RECT 240.760 88.820 241.090 89.030 ;
        RECT 241.270 88.780 241.650 89.030 ;
        RECT 241.840 89.000 242.325 89.030 ;
        RECT 241.820 88.830 242.325 89.000 ;
        RECT 236.280 87.650 236.570 88.420 ;
        RECT 237.140 88.010 238.330 88.240 ;
        RECT 237.140 87.650 237.400 88.010 ;
        RECT 237.570 87.470 237.900 87.840 ;
        RECT 238.070 87.650 238.330 88.010 ;
        RECT 238.520 87.470 238.850 88.190 ;
        RECT 239.020 87.650 239.285 88.420 ;
        RECT 239.460 87.470 239.750 88.635 ;
        RECT 240.075 88.480 241.160 88.650 ;
        RECT 240.075 87.640 240.375 88.480 ;
        RECT 240.570 87.470 240.820 88.310 ;
        RECT 240.990 88.230 241.160 88.480 ;
        RECT 241.330 88.400 241.650 88.780 ;
        RECT 241.840 88.820 242.325 88.830 ;
        RECT 242.515 88.820 242.965 89.030 ;
        RECT 243.135 88.820 243.470 89.030 ;
        RECT 241.840 88.400 242.215 88.820 ;
        RECT 243.135 88.650 243.305 88.820 ;
        RECT 242.385 88.480 243.305 88.650 ;
        RECT 242.385 88.230 242.555 88.480 ;
        RECT 240.990 88.060 242.555 88.230 ;
        RECT 241.410 87.640 242.215 88.060 ;
        RECT 242.725 87.470 243.055 88.310 ;
        RECT 243.640 88.230 243.890 89.200 ;
        RECT 245.645 88.645 245.985 89.475 ;
        RECT 249.580 89.250 253.090 90.020 ;
        RECT 253.770 89.480 253.995 89.840 ;
        RECT 254.175 89.650 254.505 90.020 ;
        RECT 254.685 89.480 254.940 89.840 ;
        RECT 255.505 89.650 256.250 90.020 ;
        RECT 253.770 89.290 256.255 89.480 ;
        RECT 243.225 87.640 243.890 88.230 ;
        RECT 247.465 87.905 247.815 89.155 ;
        RECT 249.580 88.730 251.230 89.250 ;
        RECT 251.400 88.560 253.090 89.080 ;
        RECT 253.730 88.780 254.000 89.110 ;
        RECT 254.180 88.780 254.615 89.110 ;
        RECT 254.795 88.780 255.370 89.110 ;
        RECT 255.550 88.780 255.830 89.110 ;
        RECT 256.030 88.600 256.255 89.290 ;
        RECT 244.060 87.470 249.405 87.905 ;
        RECT 249.580 87.470 253.090 88.560 ;
        RECT 253.760 88.420 256.255 88.600 ;
        RECT 256.430 88.420 256.765 89.840 ;
        RECT 253.760 87.650 254.050 88.420 ;
        RECT 254.620 88.010 255.810 88.240 ;
        RECT 254.620 87.650 254.880 88.010 ;
        RECT 255.050 87.470 255.380 87.840 ;
        RECT 255.550 87.650 255.810 88.010 ;
        RECT 256.000 87.470 256.330 88.190 ;
        RECT 256.500 87.650 256.765 88.420 ;
        RECT 256.945 89.545 257.280 89.805 ;
        RECT 257.450 89.620 257.780 90.020 ;
        RECT 257.950 89.620 259.565 89.790 ;
        RECT 256.945 88.190 257.200 89.545 ;
        RECT 257.950 89.450 258.120 89.620 ;
        RECT 257.560 89.280 258.120 89.450 ;
        RECT 258.385 89.340 258.655 89.440 ;
        RECT 257.560 89.110 257.730 89.280 ;
        RECT 258.380 89.170 258.655 89.340 ;
        RECT 257.425 88.780 257.730 89.110 ;
        RECT 257.925 89.000 258.175 89.110 ;
        RECT 257.920 88.830 258.175 89.000 ;
        RECT 257.925 88.780 258.175 88.830 ;
        RECT 258.385 88.780 258.655 89.170 ;
        RECT 258.845 88.780 259.135 89.440 ;
        RECT 259.305 88.780 259.725 89.445 ;
        RECT 260.110 89.300 260.440 90.020 ;
        RECT 260.625 89.545 260.960 89.805 ;
        RECT 261.130 89.620 261.460 90.020 ;
        RECT 261.630 89.620 263.245 89.790 ;
        RECT 260.035 89.000 260.385 89.110 ;
        RECT 260.035 88.830 260.390 89.000 ;
        RECT 260.035 88.780 260.385 88.830 ;
        RECT 257.560 88.610 257.730 88.780 ;
        RECT 257.560 88.440 259.930 88.610 ;
        RECT 260.180 88.490 260.385 88.780 ;
        RECT 256.945 87.680 257.280 88.190 ;
        RECT 257.530 87.470 257.860 88.270 ;
        RECT 258.105 88.060 259.530 88.230 ;
        RECT 258.105 87.640 258.390 88.060 ;
        RECT 258.645 87.470 258.975 87.890 ;
        RECT 259.200 87.810 259.530 88.060 ;
        RECT 259.760 87.980 259.930 88.440 ;
        RECT 260.190 87.810 260.360 88.310 ;
        RECT 259.200 87.640 260.360 87.810 ;
        RECT 260.625 88.190 260.880 89.545 ;
        RECT 261.630 89.450 261.800 89.620 ;
        RECT 261.240 89.280 261.800 89.450 ;
        RECT 262.065 89.340 262.335 89.440 ;
        RECT 261.240 89.110 261.410 89.280 ;
        RECT 262.060 89.170 262.335 89.340 ;
        RECT 261.105 88.780 261.410 89.110 ;
        RECT 261.605 89.000 261.855 89.110 ;
        RECT 261.600 88.830 261.855 89.000 ;
        RECT 261.605 88.780 261.855 88.830 ;
        RECT 262.065 88.780 262.335 89.170 ;
        RECT 262.525 89.000 262.815 89.440 ;
        RECT 262.520 88.830 262.815 89.000 ;
        RECT 262.525 88.780 262.815 88.830 ;
        RECT 262.985 88.780 263.405 89.445 ;
        RECT 263.790 89.300 264.120 90.020 ;
        RECT 265.220 89.295 265.510 90.020 ;
        RECT 265.845 89.510 266.085 90.020 ;
        RECT 266.265 89.510 266.545 89.840 ;
        RECT 266.775 89.510 266.990 90.020 ;
        RECT 263.715 89.000 264.065 89.110 ;
        RECT 263.715 88.830 264.070 89.000 ;
        RECT 263.715 88.780 264.065 88.830 ;
        RECT 265.740 88.780 266.095 89.340 ;
        RECT 261.240 88.610 261.410 88.780 ;
        RECT 261.240 88.440 263.610 88.610 ;
        RECT 263.860 88.490 264.065 88.780 ;
        RECT 260.625 87.680 260.960 88.190 ;
        RECT 261.210 87.470 261.540 88.270 ;
        RECT 261.785 88.060 263.210 88.230 ;
        RECT 261.785 87.640 262.070 88.060 ;
        RECT 262.325 87.470 262.655 87.890 ;
        RECT 262.880 87.810 263.210 88.060 ;
        RECT 263.440 87.980 263.610 88.440 ;
        RECT 263.870 87.810 264.040 88.310 ;
        RECT 262.880 87.640 264.040 87.810 ;
        RECT 265.220 87.470 265.510 88.635 ;
        RECT 266.265 88.610 266.435 89.510 ;
        RECT 266.605 88.780 266.870 89.340 ;
        RECT 267.160 89.280 267.775 89.850 ;
        RECT 267.120 88.610 267.290 89.110 ;
        RECT 265.865 88.440 267.290 88.610 ;
        RECT 265.865 88.265 266.255 88.440 ;
        RECT 266.740 87.470 267.070 88.270 ;
        RECT 267.460 88.260 267.775 89.280 ;
        RECT 267.980 89.250 269.650 90.020 ;
        RECT 270.065 89.540 270.365 90.020 ;
        RECT 270.535 89.370 270.795 89.825 ;
        RECT 270.965 89.540 271.225 90.020 ;
        RECT 271.395 89.370 271.655 89.825 ;
        RECT 271.825 89.540 272.085 90.020 ;
        RECT 272.255 89.370 272.515 89.825 ;
        RECT 272.685 89.540 272.945 90.020 ;
        RECT 273.115 89.370 273.375 89.825 ;
        RECT 273.545 89.495 273.805 90.020 ;
        RECT 267.980 88.730 268.730 89.250 ;
        RECT 270.065 89.200 273.375 89.370 ;
        RECT 268.900 88.560 269.650 89.080 ;
        RECT 267.240 87.640 267.775 88.260 ;
        RECT 267.980 87.470 269.650 88.560 ;
        RECT 270.065 88.610 271.035 89.200 ;
        RECT 273.975 89.030 274.225 89.840 ;
        RECT 274.405 89.560 274.650 90.020 ;
        RECT 274.885 89.470 275.140 89.760 ;
        RECT 275.310 89.640 275.640 90.020 ;
        RECT 271.205 88.780 274.225 89.030 ;
        RECT 274.395 88.780 274.710 89.390 ;
        RECT 274.885 89.300 275.635 89.470 ;
        RECT 270.065 88.370 273.375 88.610 ;
        RECT 270.070 87.470 270.365 88.200 ;
        RECT 270.535 87.645 270.795 88.370 ;
        RECT 270.965 87.470 271.225 88.200 ;
        RECT 271.395 87.645 271.655 88.370 ;
        RECT 271.825 87.470 272.085 88.200 ;
        RECT 272.255 87.645 272.515 88.370 ;
        RECT 272.685 87.470 272.945 88.200 ;
        RECT 273.115 87.645 273.375 88.370 ;
        RECT 273.545 87.470 273.805 88.580 ;
        RECT 273.975 87.645 274.225 88.780 ;
        RECT 274.405 87.470 274.700 88.580 ;
        RECT 274.885 88.480 275.235 89.130 ;
        RECT 275.405 88.310 275.635 89.300 ;
        RECT 274.885 88.140 275.635 88.310 ;
        RECT 274.885 87.640 275.140 88.140 ;
        RECT 275.310 87.470 275.640 87.970 ;
        RECT 275.810 87.640 275.980 89.760 ;
        RECT 276.340 89.660 276.670 90.020 ;
        RECT 276.840 89.630 277.335 89.800 ;
        RECT 277.540 89.630 278.395 89.800 ;
        RECT 276.210 88.440 276.670 89.490 ;
        RECT 276.150 87.655 276.475 88.440 ;
        RECT 276.840 88.270 277.010 89.630 ;
        RECT 277.180 88.720 277.530 89.340 ;
        RECT 277.700 89.120 278.055 89.340 ;
        RECT 277.700 88.530 277.870 89.120 ;
        RECT 278.225 88.920 278.395 89.630 ;
        RECT 279.270 89.560 279.600 90.020 ;
        RECT 279.810 89.660 280.160 89.830 ;
        RECT 278.600 89.090 279.390 89.340 ;
        RECT 279.810 89.270 280.070 89.660 ;
        RECT 280.380 89.570 281.330 89.850 ;
        RECT 281.500 89.580 281.690 90.020 ;
        RECT 281.860 89.640 282.930 89.810 ;
        RECT 279.560 88.920 279.730 89.100 ;
        RECT 276.840 88.100 277.235 88.270 ;
        RECT 277.405 88.140 277.870 88.530 ;
        RECT 278.040 88.750 279.730 88.920 ;
        RECT 277.065 87.970 277.235 88.100 ;
        RECT 278.040 87.970 278.210 88.750 ;
        RECT 279.900 88.580 280.070 89.270 ;
        RECT 278.570 88.410 280.070 88.580 ;
        RECT 280.260 88.610 280.470 89.400 ;
        RECT 280.640 88.780 280.990 89.400 ;
        RECT 281.160 88.790 281.330 89.570 ;
        RECT 281.860 89.410 282.030 89.640 ;
        RECT 281.500 89.240 282.030 89.410 ;
        RECT 281.500 88.960 281.720 89.240 ;
        RECT 282.200 89.070 282.440 89.470 ;
        RECT 281.160 88.620 281.565 88.790 ;
        RECT 281.900 88.700 282.440 89.070 ;
        RECT 282.610 89.285 282.930 89.640 ;
        RECT 283.175 89.560 283.480 90.020 ;
        RECT 283.650 89.310 283.905 89.840 ;
        RECT 282.610 89.110 282.935 89.285 ;
        RECT 282.610 88.810 283.525 89.110 ;
        RECT 282.785 88.780 283.525 88.810 ;
        RECT 280.260 88.450 280.935 88.610 ;
        RECT 281.395 88.530 281.565 88.620 ;
        RECT 280.260 88.440 281.225 88.450 ;
        RECT 279.900 88.270 280.070 88.410 ;
        RECT 276.645 87.470 276.895 87.930 ;
        RECT 277.065 87.640 277.315 87.970 ;
        RECT 277.530 87.640 278.210 87.970 ;
        RECT 278.380 88.070 279.455 88.240 ;
        RECT 279.900 88.100 280.460 88.270 ;
        RECT 280.765 88.150 281.225 88.440 ;
        RECT 281.395 88.360 282.615 88.530 ;
        RECT 278.380 87.730 278.550 88.070 ;
        RECT 278.785 87.470 279.115 87.900 ;
        RECT 279.285 87.730 279.455 88.070 ;
        RECT 279.750 87.470 280.120 87.930 ;
        RECT 280.290 87.640 280.460 88.100 ;
        RECT 281.395 87.980 281.565 88.360 ;
        RECT 282.785 88.190 282.955 88.780 ;
        RECT 283.695 88.660 283.905 89.310 ;
        RECT 280.695 87.640 281.565 87.980 ;
        RECT 282.155 88.020 282.955 88.190 ;
        RECT 281.735 87.470 281.985 87.930 ;
        RECT 282.155 87.730 282.325 88.020 ;
        RECT 282.505 87.470 282.835 87.850 ;
        RECT 283.175 87.470 283.480 88.610 ;
        RECT 283.650 87.780 283.905 88.660 ;
        RECT 284.085 89.280 284.340 89.850 ;
        RECT 284.510 89.620 284.840 90.020 ;
        RECT 285.265 89.485 285.795 89.850 ;
        RECT 285.265 89.450 285.440 89.485 ;
        RECT 284.510 89.280 285.440 89.450 ;
        RECT 284.085 88.610 284.255 89.280 ;
        RECT 284.510 89.110 284.680 89.280 ;
        RECT 284.425 88.780 284.680 89.110 ;
        RECT 284.905 88.780 285.100 89.110 ;
        RECT 284.085 87.640 284.420 88.610 ;
        RECT 284.590 87.470 284.760 88.610 ;
        RECT 284.930 87.810 285.100 88.780 ;
        RECT 285.270 88.150 285.440 89.280 ;
        RECT 285.610 88.490 285.780 89.290 ;
        RECT 285.985 89.000 286.260 89.850 ;
        RECT 285.980 88.830 286.260 89.000 ;
        RECT 285.985 88.690 286.260 88.830 ;
        RECT 286.430 88.490 286.620 89.850 ;
        RECT 286.800 89.485 287.310 90.020 ;
        RECT 287.530 89.210 287.775 89.815 ;
        RECT 288.220 89.270 289.430 90.020 ;
        RECT 289.690 89.470 289.860 89.850 ;
        RECT 290.040 89.640 290.370 90.020 ;
        RECT 289.690 89.300 290.355 89.470 ;
        RECT 290.550 89.345 290.810 89.850 ;
        RECT 286.820 89.040 288.050 89.210 ;
        RECT 285.610 88.320 286.620 88.490 ;
        RECT 286.790 88.475 287.540 88.665 ;
        RECT 285.270 87.980 286.395 88.150 ;
        RECT 286.790 87.810 286.960 88.475 ;
        RECT 287.710 88.230 288.050 89.040 ;
        RECT 288.220 88.730 288.740 89.270 ;
        RECT 288.910 88.560 289.430 89.100 ;
        RECT 289.620 88.750 289.950 89.120 ;
        RECT 290.185 89.045 290.355 89.300 ;
        RECT 290.185 88.715 290.470 89.045 ;
        RECT 290.185 88.570 290.355 88.715 ;
        RECT 284.930 87.640 286.960 87.810 ;
        RECT 287.130 87.470 287.300 88.230 ;
        RECT 287.535 87.820 288.050 88.230 ;
        RECT 288.220 87.470 289.430 88.560 ;
        RECT 289.690 88.400 290.355 88.570 ;
        RECT 290.640 88.545 290.810 89.345 ;
        RECT 290.980 89.295 291.270 90.020 ;
        RECT 291.445 89.470 291.700 89.760 ;
        RECT 291.870 89.640 292.200 90.020 ;
        RECT 291.445 89.300 292.195 89.470 ;
        RECT 289.690 87.640 289.860 88.400 ;
        RECT 290.040 87.470 290.370 88.230 ;
        RECT 290.540 87.640 290.810 88.545 ;
        RECT 290.980 87.470 291.270 88.635 ;
        RECT 291.445 88.480 291.795 89.130 ;
        RECT 291.965 88.310 292.195 89.300 ;
        RECT 291.445 88.140 292.195 88.310 ;
        RECT 291.445 87.640 291.700 88.140 ;
        RECT 291.870 87.470 292.200 87.970 ;
        RECT 292.370 87.640 292.540 89.760 ;
        RECT 292.900 89.660 293.230 90.020 ;
        RECT 293.400 89.630 293.895 89.800 ;
        RECT 294.100 89.630 294.955 89.800 ;
        RECT 292.770 88.440 293.230 89.490 ;
        RECT 292.710 87.655 293.035 88.440 ;
        RECT 293.400 88.270 293.570 89.630 ;
        RECT 293.740 88.720 294.090 89.340 ;
        RECT 294.260 89.120 294.615 89.340 ;
        RECT 294.260 88.530 294.430 89.120 ;
        RECT 294.785 88.920 294.955 89.630 ;
        RECT 295.830 89.560 296.160 90.020 ;
        RECT 296.370 89.660 296.720 89.830 ;
        RECT 295.160 89.090 295.950 89.340 ;
        RECT 296.370 89.270 296.630 89.660 ;
        RECT 296.940 89.570 297.890 89.850 ;
        RECT 298.060 89.580 298.250 90.020 ;
        RECT 298.420 89.640 299.490 89.810 ;
        RECT 296.120 88.920 296.290 89.100 ;
        RECT 293.400 88.100 293.795 88.270 ;
        RECT 293.965 88.140 294.430 88.530 ;
        RECT 294.600 88.750 296.290 88.920 ;
        RECT 293.625 87.970 293.795 88.100 ;
        RECT 294.600 87.970 294.770 88.750 ;
        RECT 296.460 88.580 296.630 89.270 ;
        RECT 295.130 88.410 296.630 88.580 ;
        RECT 296.820 88.610 297.030 89.400 ;
        RECT 297.200 88.780 297.550 89.400 ;
        RECT 297.720 88.790 297.890 89.570 ;
        RECT 298.420 89.410 298.590 89.640 ;
        RECT 298.060 89.240 298.590 89.410 ;
        RECT 298.060 88.960 298.280 89.240 ;
        RECT 298.760 89.070 299.000 89.470 ;
        RECT 297.720 88.620 298.125 88.790 ;
        RECT 298.460 88.700 299.000 89.070 ;
        RECT 299.170 89.285 299.490 89.640 ;
        RECT 299.735 89.560 300.040 90.020 ;
        RECT 300.210 89.310 300.465 89.840 ;
        RECT 299.170 89.110 299.495 89.285 ;
        RECT 299.170 88.810 300.085 89.110 ;
        RECT 299.345 88.780 300.085 88.810 ;
        RECT 296.820 88.450 297.495 88.610 ;
        RECT 297.955 88.530 298.125 88.620 ;
        RECT 296.820 88.440 297.785 88.450 ;
        RECT 296.460 88.270 296.630 88.410 ;
        RECT 293.205 87.470 293.455 87.930 ;
        RECT 293.625 87.640 293.875 87.970 ;
        RECT 294.090 87.640 294.770 87.970 ;
        RECT 294.940 88.070 296.015 88.240 ;
        RECT 296.460 88.100 297.020 88.270 ;
        RECT 297.325 88.150 297.785 88.440 ;
        RECT 297.955 88.360 299.175 88.530 ;
        RECT 294.940 87.730 295.110 88.070 ;
        RECT 295.345 87.470 295.675 87.900 ;
        RECT 295.845 87.730 296.015 88.070 ;
        RECT 296.310 87.470 296.680 87.930 ;
        RECT 296.850 87.640 297.020 88.100 ;
        RECT 297.955 87.980 298.125 88.360 ;
        RECT 299.345 88.190 299.515 88.780 ;
        RECT 300.255 88.660 300.465 89.310 ;
        RECT 300.645 89.470 300.900 89.760 ;
        RECT 301.070 89.640 301.400 90.020 ;
        RECT 300.645 89.300 301.395 89.470 ;
        RECT 297.255 87.640 298.125 87.980 ;
        RECT 298.715 88.020 299.515 88.190 ;
        RECT 298.295 87.470 298.545 87.930 ;
        RECT 298.715 87.730 298.885 88.020 ;
        RECT 299.065 87.470 299.395 87.850 ;
        RECT 299.735 87.470 300.040 88.610 ;
        RECT 300.210 87.780 300.465 88.660 ;
        RECT 300.645 88.480 300.995 89.130 ;
        RECT 301.165 88.310 301.395 89.300 ;
        RECT 300.645 88.140 301.395 88.310 ;
        RECT 300.645 87.640 300.900 88.140 ;
        RECT 301.070 87.470 301.400 87.970 ;
        RECT 301.570 87.640 301.740 89.760 ;
        RECT 302.100 89.660 302.430 90.020 ;
        RECT 302.600 89.630 303.095 89.800 ;
        RECT 303.300 89.630 304.155 89.800 ;
        RECT 301.970 88.440 302.430 89.490 ;
        RECT 301.910 87.655 302.235 88.440 ;
        RECT 302.600 88.270 302.770 89.630 ;
        RECT 302.940 88.720 303.290 89.340 ;
        RECT 303.460 89.120 303.815 89.340 ;
        RECT 303.460 88.530 303.630 89.120 ;
        RECT 303.985 88.920 304.155 89.630 ;
        RECT 305.030 89.560 305.360 90.020 ;
        RECT 305.570 89.660 305.920 89.830 ;
        RECT 304.360 89.090 305.150 89.340 ;
        RECT 305.570 89.270 305.830 89.660 ;
        RECT 306.140 89.570 307.090 89.850 ;
        RECT 307.260 89.580 307.450 90.020 ;
        RECT 307.620 89.640 308.690 89.810 ;
        RECT 305.320 88.920 305.490 89.100 ;
        RECT 302.600 88.100 302.995 88.270 ;
        RECT 303.165 88.140 303.630 88.530 ;
        RECT 303.800 88.750 305.490 88.920 ;
        RECT 302.825 87.970 302.995 88.100 ;
        RECT 303.800 87.970 303.970 88.750 ;
        RECT 305.660 88.580 305.830 89.270 ;
        RECT 304.330 88.410 305.830 88.580 ;
        RECT 306.020 88.610 306.230 89.400 ;
        RECT 306.400 88.780 306.750 89.400 ;
        RECT 306.920 88.790 307.090 89.570 ;
        RECT 307.620 89.410 307.790 89.640 ;
        RECT 307.260 89.240 307.790 89.410 ;
        RECT 307.260 88.960 307.480 89.240 ;
        RECT 307.960 89.070 308.200 89.470 ;
        RECT 306.920 88.620 307.325 88.790 ;
        RECT 307.660 88.700 308.200 89.070 ;
        RECT 308.370 89.285 308.690 89.640 ;
        RECT 308.935 89.560 309.240 90.020 ;
        RECT 309.410 89.310 309.665 89.840 ;
        RECT 308.370 89.110 308.695 89.285 ;
        RECT 308.370 88.810 309.285 89.110 ;
        RECT 308.545 88.780 309.285 88.810 ;
        RECT 306.020 88.450 306.695 88.610 ;
        RECT 307.155 88.530 307.325 88.620 ;
        RECT 306.020 88.440 306.985 88.450 ;
        RECT 305.660 88.270 305.830 88.410 ;
        RECT 302.405 87.470 302.655 87.930 ;
        RECT 302.825 87.640 303.075 87.970 ;
        RECT 303.290 87.640 303.970 87.970 ;
        RECT 304.140 88.070 305.215 88.240 ;
        RECT 305.660 88.100 306.220 88.270 ;
        RECT 306.525 88.150 306.985 88.440 ;
        RECT 307.155 88.360 308.375 88.530 ;
        RECT 304.140 87.730 304.310 88.070 ;
        RECT 304.545 87.470 304.875 87.900 ;
        RECT 305.045 87.730 305.215 88.070 ;
        RECT 305.510 87.470 305.880 87.930 ;
        RECT 306.050 87.640 306.220 88.100 ;
        RECT 307.155 87.980 307.325 88.360 ;
        RECT 308.545 88.190 308.715 88.780 ;
        RECT 309.455 88.660 309.665 89.310 ;
        RECT 309.840 89.270 311.050 90.020 ;
        RECT 306.455 87.640 307.325 87.980 ;
        RECT 307.915 88.020 308.715 88.190 ;
        RECT 307.495 87.470 307.745 87.930 ;
        RECT 307.915 87.730 308.085 88.020 ;
        RECT 308.265 87.470 308.595 87.850 ;
        RECT 308.935 87.470 309.240 88.610 ;
        RECT 309.410 87.780 309.665 88.660 ;
        RECT 309.840 88.560 310.360 89.100 ;
        RECT 310.530 88.730 311.050 89.270 ;
        RECT 309.840 87.470 311.050 88.560 ;
        RECT 162.095 87.300 311.135 87.470 ;
        RECT 162.180 86.210 163.390 87.300 ;
        RECT 163.560 86.865 168.905 87.300 ;
        RECT 162.180 85.500 162.700 86.040 ;
        RECT 162.870 85.670 163.390 86.210 ;
        RECT 162.180 84.750 163.390 85.500 ;
        RECT 165.145 85.295 165.485 86.125 ;
        RECT 166.965 85.615 167.315 86.865 ;
        RECT 169.630 86.370 169.800 87.130 ;
        RECT 169.980 86.540 170.310 87.300 ;
        RECT 169.630 86.200 170.295 86.370 ;
        RECT 170.480 86.225 170.750 87.130 ;
        RECT 170.125 86.055 170.295 86.200 ;
        RECT 169.560 85.650 169.890 86.020 ;
        RECT 170.125 85.725 170.410 86.055 ;
        RECT 170.125 85.470 170.295 85.725 ;
        RECT 169.630 85.300 170.295 85.470 ;
        RECT 170.580 85.425 170.750 86.225 ;
        RECT 163.560 84.750 168.905 85.295 ;
        RECT 169.630 84.920 169.800 85.300 ;
        RECT 169.980 84.750 170.310 85.130 ;
        RECT 170.490 84.920 170.750 85.425 ;
        RECT 170.925 86.160 171.260 87.130 ;
        RECT 171.430 86.160 171.600 87.300 ;
        RECT 171.770 86.960 173.800 87.130 ;
        RECT 170.925 85.490 171.095 86.160 ;
        RECT 171.770 85.990 171.940 86.960 ;
        RECT 171.265 85.660 171.520 85.990 ;
        RECT 171.745 85.660 171.940 85.990 ;
        RECT 172.110 86.620 173.235 86.790 ;
        RECT 171.350 85.490 171.520 85.660 ;
        RECT 172.110 85.490 172.280 86.620 ;
        RECT 170.925 84.920 171.180 85.490 ;
        RECT 171.350 85.320 172.280 85.490 ;
        RECT 172.450 86.280 173.460 86.450 ;
        RECT 172.450 85.480 172.620 86.280 ;
        RECT 172.825 85.940 173.100 86.080 ;
        RECT 172.820 85.770 173.100 85.940 ;
        RECT 172.105 85.285 172.280 85.320 ;
        RECT 171.350 84.750 171.680 85.150 ;
        RECT 172.105 84.920 172.635 85.285 ;
        RECT 172.825 84.920 173.100 85.770 ;
        RECT 173.270 84.920 173.460 86.280 ;
        RECT 173.630 86.295 173.800 86.960 ;
        RECT 173.970 86.540 174.140 87.300 ;
        RECT 174.375 86.540 174.890 86.950 ;
        RECT 173.630 86.105 174.380 86.295 ;
        RECT 174.550 85.730 174.890 86.540 ;
        RECT 175.060 86.135 175.350 87.300 ;
        RECT 175.525 86.160 175.860 87.130 ;
        RECT 176.030 86.160 176.200 87.300 ;
        RECT 176.370 86.960 178.400 87.130 ;
        RECT 173.660 85.560 174.890 85.730 ;
        RECT 173.640 84.750 174.150 85.285 ;
        RECT 174.370 84.955 174.615 85.560 ;
        RECT 175.525 85.490 175.695 86.160 ;
        RECT 176.370 85.990 176.540 86.960 ;
        RECT 175.865 85.660 176.120 85.990 ;
        RECT 176.345 85.660 176.540 85.990 ;
        RECT 176.710 86.620 177.835 86.790 ;
        RECT 175.950 85.490 176.120 85.660 ;
        RECT 176.710 85.490 176.880 86.620 ;
        RECT 175.060 84.750 175.350 85.475 ;
        RECT 175.525 84.920 175.780 85.490 ;
        RECT 175.950 85.320 176.880 85.490 ;
        RECT 177.050 86.280 178.060 86.450 ;
        RECT 177.050 85.480 177.220 86.280 ;
        RECT 177.425 85.940 177.700 86.080 ;
        RECT 177.420 85.770 177.700 85.940 ;
        RECT 176.705 85.285 176.880 85.320 ;
        RECT 175.950 84.750 176.280 85.150 ;
        RECT 176.705 84.920 177.235 85.285 ;
        RECT 177.425 84.920 177.700 85.770 ;
        RECT 177.870 84.920 178.060 86.280 ;
        RECT 178.230 86.295 178.400 86.960 ;
        RECT 178.570 86.540 178.740 87.300 ;
        RECT 178.975 86.540 179.490 86.950 ;
        RECT 178.230 86.105 178.980 86.295 ;
        RECT 179.150 85.730 179.490 86.540 ;
        RECT 179.660 86.210 183.170 87.300 ;
        RECT 184.265 86.630 184.520 87.130 ;
        RECT 184.690 86.800 185.020 87.300 ;
        RECT 184.265 86.460 185.015 86.630 ;
        RECT 178.260 85.560 179.490 85.730 ;
        RECT 178.240 84.750 178.750 85.285 ;
        RECT 178.970 84.955 179.215 85.560 ;
        RECT 179.660 85.520 181.310 86.040 ;
        RECT 181.480 85.690 183.170 86.210 ;
        RECT 184.265 85.640 184.615 86.290 ;
        RECT 179.660 84.750 183.170 85.520 ;
        RECT 184.785 85.470 185.015 86.460 ;
        RECT 184.265 85.300 185.015 85.470 ;
        RECT 184.265 85.010 184.520 85.300 ;
        RECT 184.690 84.750 185.020 85.130 ;
        RECT 185.190 85.010 185.360 87.130 ;
        RECT 185.530 86.330 185.855 87.115 ;
        RECT 186.025 86.840 186.275 87.300 ;
        RECT 186.445 86.800 186.695 87.130 ;
        RECT 186.910 86.800 187.590 87.130 ;
        RECT 186.445 86.670 186.615 86.800 ;
        RECT 186.220 86.500 186.615 86.670 ;
        RECT 185.590 85.280 186.050 86.330 ;
        RECT 186.220 85.140 186.390 86.500 ;
        RECT 186.785 86.240 187.250 86.630 ;
        RECT 186.560 85.430 186.910 86.050 ;
        RECT 187.080 85.650 187.250 86.240 ;
        RECT 187.420 86.020 187.590 86.800 ;
        RECT 187.760 86.700 187.930 87.040 ;
        RECT 188.165 86.870 188.495 87.300 ;
        RECT 188.665 86.700 188.835 87.040 ;
        RECT 189.130 86.840 189.500 87.300 ;
        RECT 187.760 86.530 188.835 86.700 ;
        RECT 189.670 86.670 189.840 87.130 ;
        RECT 190.075 86.790 190.945 87.130 ;
        RECT 191.115 86.840 191.365 87.300 ;
        RECT 189.280 86.500 189.840 86.670 ;
        RECT 189.280 86.360 189.450 86.500 ;
        RECT 187.950 86.190 189.450 86.360 ;
        RECT 190.145 86.330 190.605 86.620 ;
        RECT 187.420 85.850 189.110 86.020 ;
        RECT 187.080 85.430 187.435 85.650 ;
        RECT 187.605 85.140 187.775 85.850 ;
        RECT 187.980 85.430 188.770 85.680 ;
        RECT 188.940 85.670 189.110 85.850 ;
        RECT 189.280 85.500 189.450 86.190 ;
        RECT 185.720 84.750 186.050 85.110 ;
        RECT 186.220 84.970 186.715 85.140 ;
        RECT 186.920 84.970 187.775 85.140 ;
        RECT 188.650 84.750 188.980 85.210 ;
        RECT 189.190 85.110 189.450 85.500 ;
        RECT 189.640 86.320 190.605 86.330 ;
        RECT 190.775 86.410 190.945 86.790 ;
        RECT 191.535 86.750 191.705 87.040 ;
        RECT 191.885 86.920 192.215 87.300 ;
        RECT 191.535 86.580 192.335 86.750 ;
        RECT 189.640 86.160 190.315 86.320 ;
        RECT 190.775 86.240 191.995 86.410 ;
        RECT 189.640 85.370 189.850 86.160 ;
        RECT 190.775 86.150 190.945 86.240 ;
        RECT 190.020 85.370 190.370 85.990 ;
        RECT 190.540 85.980 190.945 86.150 ;
        RECT 190.540 85.200 190.710 85.980 ;
        RECT 190.880 85.530 191.100 85.810 ;
        RECT 191.280 85.700 191.820 86.070 ;
        RECT 192.165 85.990 192.335 86.580 ;
        RECT 192.555 86.160 192.860 87.300 ;
        RECT 193.030 86.110 193.280 86.990 ;
        RECT 193.450 86.160 193.700 87.300 ;
        RECT 193.920 86.865 199.265 87.300 ;
        RECT 192.165 85.960 192.905 85.990 ;
        RECT 190.880 85.360 191.410 85.530 ;
        RECT 189.190 84.940 189.540 85.110 ;
        RECT 189.760 84.920 190.710 85.200 ;
        RECT 190.880 84.750 191.070 85.190 ;
        RECT 191.240 85.130 191.410 85.360 ;
        RECT 191.580 85.300 191.820 85.700 ;
        RECT 191.990 85.660 192.905 85.960 ;
        RECT 191.990 85.485 192.315 85.660 ;
        RECT 191.990 85.130 192.310 85.485 ;
        RECT 193.075 85.460 193.280 86.110 ;
        RECT 191.240 84.960 192.310 85.130 ;
        RECT 192.555 84.750 192.860 85.210 ;
        RECT 193.030 84.930 193.280 85.460 ;
        RECT 193.450 84.750 193.700 85.505 ;
        RECT 195.505 85.295 195.845 86.125 ;
        RECT 197.325 85.615 197.675 86.865 ;
        RECT 199.440 86.210 200.650 87.300 ;
        RECT 199.440 85.500 199.960 86.040 ;
        RECT 200.130 85.670 200.650 86.210 ;
        RECT 200.820 86.135 201.110 87.300 ;
        RECT 201.280 85.695 201.560 87.130 ;
        RECT 201.730 86.525 202.440 87.300 ;
        RECT 202.610 86.355 202.940 87.130 ;
        RECT 201.790 86.140 202.940 86.355 ;
        RECT 193.920 84.750 199.265 85.295 ;
        RECT 199.440 84.750 200.650 85.500 ;
        RECT 200.820 84.750 201.110 85.475 ;
        RECT 201.280 84.920 201.620 85.695 ;
        RECT 201.790 85.570 202.075 86.140 ;
        RECT 202.260 85.740 202.730 85.970 ;
        RECT 203.135 85.940 203.350 87.055 ;
        RECT 203.530 86.580 203.860 87.300 ;
        RECT 204.500 86.330 204.770 87.100 ;
        RECT 204.940 86.520 205.270 87.300 ;
        RECT 205.475 86.695 205.660 87.100 ;
        RECT 205.830 86.875 206.165 87.300 ;
        RECT 206.345 86.945 207.425 87.115 ;
        RECT 205.475 86.520 206.140 86.695 ;
        RECT 203.640 85.940 203.870 86.280 ;
        RECT 202.900 85.760 203.350 85.940 ;
        RECT 202.900 85.740 203.230 85.760 ;
        RECT 203.540 85.740 203.870 85.940 ;
        RECT 204.500 86.160 205.630 86.330 ;
        RECT 201.790 85.380 202.500 85.570 ;
        RECT 202.200 85.240 202.500 85.380 ;
        RECT 202.690 85.380 203.870 85.570 ;
        RECT 202.690 85.300 203.020 85.380 ;
        RECT 202.200 85.230 202.515 85.240 ;
        RECT 202.200 85.220 202.525 85.230 ;
        RECT 202.200 85.215 202.535 85.220 ;
        RECT 201.790 84.750 201.960 85.210 ;
        RECT 202.200 85.205 202.540 85.215 ;
        RECT 202.200 85.200 202.545 85.205 ;
        RECT 202.200 85.190 202.550 85.200 ;
        RECT 202.200 85.185 202.555 85.190 ;
        RECT 202.200 84.920 202.560 85.185 ;
        RECT 203.190 84.750 203.360 85.210 ;
        RECT 203.530 84.920 203.870 85.380 ;
        RECT 204.500 85.250 204.670 86.160 ;
        RECT 204.840 85.410 205.200 85.990 ;
        RECT 205.380 85.660 205.630 86.160 ;
        RECT 205.800 85.490 206.140 86.520 ;
        RECT 206.345 86.160 206.680 86.945 ;
        RECT 206.850 85.990 207.085 86.670 ;
        RECT 207.255 86.330 207.425 86.945 ;
        RECT 207.690 86.500 208.005 87.300 ;
        RECT 207.255 86.160 207.570 86.330 ;
        RECT 206.345 85.660 206.680 85.990 ;
        RECT 206.850 85.660 207.230 85.990 ;
        RECT 207.400 85.490 207.570 86.160 ;
        RECT 205.455 85.320 206.140 85.490 ;
        RECT 206.345 85.320 207.570 85.490 ;
        RECT 207.740 85.320 208.010 86.330 ;
        RECT 208.180 86.160 208.470 87.300 ;
        RECT 208.640 86.580 209.090 87.130 ;
        RECT 209.280 86.580 209.610 87.300 ;
        RECT 204.500 84.920 204.760 85.250 ;
        RECT 204.970 84.750 205.245 85.230 ;
        RECT 205.455 84.920 205.660 85.320 ;
        RECT 205.830 84.750 206.165 85.150 ;
        RECT 206.345 85.050 206.600 85.320 ;
        RECT 206.770 84.750 207.100 85.150 ;
        RECT 207.270 85.050 207.440 85.320 ;
        RECT 207.610 84.750 207.940 85.150 ;
        RECT 208.180 84.750 208.470 85.550 ;
        RECT 208.640 85.210 208.890 86.580 ;
        RECT 209.820 86.410 210.120 86.960 ;
        RECT 210.290 86.630 210.570 87.300 ;
        RECT 209.180 86.240 210.120 86.410 ;
        RECT 209.180 85.990 209.350 86.240 ;
        RECT 210.455 85.990 210.770 86.430 ;
        RECT 209.060 85.660 209.350 85.990 ;
        RECT 209.520 85.740 209.850 85.990 ;
        RECT 210.080 85.740 210.770 85.990 ;
        RECT 210.940 86.330 211.210 87.100 ;
        RECT 211.380 86.520 211.710 87.300 ;
        RECT 211.915 86.695 212.100 87.100 ;
        RECT 212.270 86.875 212.605 87.300 ;
        RECT 212.780 86.865 218.125 87.300 ;
        RECT 211.915 86.520 212.580 86.695 ;
        RECT 210.940 86.160 212.070 86.330 ;
        RECT 209.180 85.570 209.350 85.660 ;
        RECT 209.180 85.380 210.570 85.570 ;
        RECT 208.640 84.920 209.190 85.210 ;
        RECT 209.360 84.750 209.610 85.210 ;
        RECT 210.240 85.020 210.570 85.380 ;
        RECT 210.940 85.250 211.110 86.160 ;
        RECT 211.280 85.410 211.640 85.990 ;
        RECT 211.820 85.660 212.070 86.160 ;
        RECT 212.240 85.490 212.580 86.520 ;
        RECT 211.895 85.320 212.580 85.490 ;
        RECT 210.940 84.920 211.200 85.250 ;
        RECT 211.410 84.750 211.685 85.230 ;
        RECT 211.895 84.920 212.100 85.320 ;
        RECT 214.365 85.295 214.705 86.125 ;
        RECT 216.185 85.615 216.535 86.865 ;
        RECT 218.300 86.210 219.970 87.300 ;
        RECT 218.300 85.520 219.050 86.040 ;
        RECT 219.220 85.690 219.970 86.210 ;
        RECT 220.665 86.290 220.920 87.130 ;
        RECT 221.090 86.460 221.340 87.300 ;
        RECT 221.510 86.290 221.760 87.130 ;
        RECT 221.930 86.460 222.180 87.300 ;
        RECT 222.350 86.750 223.440 87.130 ;
        RECT 222.350 86.290 222.600 86.750 ;
        RECT 220.665 86.120 222.600 86.290 ;
        RECT 222.770 86.290 223.020 86.580 ;
        RECT 223.190 86.460 223.440 86.750 ;
        RECT 223.610 86.960 225.540 87.130 ;
        RECT 223.610 86.290 223.860 86.960 ;
        RECT 224.450 86.800 224.700 86.960 ;
        RECT 225.290 86.800 225.540 86.960 ;
        RECT 225.710 86.790 225.960 87.130 ;
        RECT 224.030 86.630 224.280 86.790 ;
        RECT 224.870 86.630 225.120 86.790 ;
        RECT 224.030 86.620 225.120 86.630 ;
        RECT 226.130 86.620 226.410 87.130 ;
        RECT 224.030 86.450 226.410 86.620 ;
        RECT 222.770 86.120 223.860 86.290 ;
        RECT 224.030 86.110 225.680 86.280 ;
        RECT 224.030 85.950 224.200 86.110 ;
        RECT 220.605 85.740 222.340 85.950 ;
        RECT 222.610 85.740 224.200 85.950 ;
        RECT 225.510 85.950 225.680 86.110 ;
        RECT 224.370 85.740 225.280 85.940 ;
        RECT 225.510 85.740 225.930 85.950 ;
        RECT 226.120 85.570 226.410 86.450 ;
        RECT 226.580 86.135 226.870 87.300 ;
        RECT 227.040 86.865 232.385 87.300 ;
        RECT 212.270 84.750 212.605 85.150 ;
        RECT 212.780 84.750 218.125 85.295 ;
        RECT 218.300 84.750 219.970 85.520 ;
        RECT 220.605 84.750 220.880 85.570 ;
        RECT 221.050 85.390 226.410 85.570 ;
        RECT 221.050 84.920 221.380 85.390 ;
        RECT 221.550 84.750 221.720 85.220 ;
        RECT 221.890 84.920 222.220 85.390 ;
        RECT 222.390 84.750 222.560 85.220 ;
        RECT 222.730 84.920 223.060 85.390 ;
        RECT 223.230 84.750 223.400 85.220 ;
        RECT 223.570 84.920 223.900 85.390 ;
        RECT 224.070 84.750 224.240 85.220 ;
        RECT 224.410 84.920 224.740 85.390 ;
        RECT 224.910 84.750 225.080 85.220 ;
        RECT 225.250 84.920 225.580 85.390 ;
        RECT 225.750 84.750 225.920 85.220 ;
        RECT 226.120 84.920 226.410 85.390 ;
        RECT 226.580 84.750 226.870 85.475 ;
        RECT 228.625 85.295 228.965 86.125 ;
        RECT 230.445 85.615 230.795 86.865 ;
        RECT 233.025 86.330 233.300 87.130 ;
        RECT 233.470 86.500 233.800 87.300 ;
        RECT 233.970 86.330 234.140 87.130 ;
        RECT 234.310 86.500 234.560 87.300 ;
        RECT 234.730 86.960 236.825 87.130 ;
        RECT 234.730 86.330 235.060 86.960 ;
        RECT 233.025 86.120 235.060 86.330 ;
        RECT 235.230 86.410 235.400 86.790 ;
        RECT 235.570 86.600 235.900 86.960 ;
        RECT 236.070 86.410 236.240 86.790 ;
        RECT 236.410 86.580 236.825 86.960 ;
        RECT 235.230 86.110 236.990 86.410 ;
        RECT 237.160 86.210 238.370 87.300 ;
        RECT 233.075 85.740 234.735 85.940 ;
        RECT 235.055 85.740 236.420 85.940 ;
        RECT 236.590 85.570 236.990 86.110 ;
        RECT 227.040 84.750 232.385 85.295 ;
        RECT 233.025 84.750 233.300 85.570 ;
        RECT 233.470 85.390 236.990 85.570 ;
        RECT 237.160 85.500 237.680 86.040 ;
        RECT 237.850 85.670 238.370 86.210 ;
        RECT 238.545 86.580 238.880 87.090 ;
        RECT 233.470 84.920 233.800 85.390 ;
        RECT 233.970 84.750 234.140 85.220 ;
        RECT 234.310 84.920 234.640 85.390 ;
        RECT 234.810 84.750 234.980 85.220 ;
        RECT 235.150 84.920 235.480 85.390 ;
        RECT 235.650 84.750 235.820 85.220 ;
        RECT 235.990 84.920 236.320 85.390 ;
        RECT 236.490 84.750 236.775 85.220 ;
        RECT 237.160 84.750 238.370 85.500 ;
        RECT 238.545 85.225 238.800 86.580 ;
        RECT 239.130 86.500 239.460 87.300 ;
        RECT 239.705 86.710 239.990 87.130 ;
        RECT 240.245 86.880 240.575 87.300 ;
        RECT 240.800 86.960 241.960 87.130 ;
        RECT 240.800 86.710 241.130 86.960 ;
        RECT 239.705 86.540 241.130 86.710 ;
        RECT 241.360 86.330 241.530 86.790 ;
        RECT 241.790 86.460 241.960 86.960 ;
        RECT 239.160 86.160 241.530 86.330 ;
        RECT 242.405 86.330 242.795 86.505 ;
        RECT 243.280 86.500 243.610 87.300 ;
        RECT 243.780 86.510 244.315 87.130 ;
        RECT 244.520 86.865 249.865 87.300 ;
        RECT 239.160 85.990 239.330 86.160 ;
        RECT 241.780 86.110 241.990 86.280 ;
        RECT 242.405 86.160 243.830 86.330 ;
        RECT 241.780 85.990 241.985 86.110 ;
        RECT 239.025 85.660 239.330 85.990 ;
        RECT 239.525 85.660 239.775 85.990 ;
        RECT 239.160 85.490 239.330 85.660 ;
        RECT 239.985 85.600 240.255 85.990 ;
        RECT 240.445 85.600 240.735 85.990 ;
        RECT 239.160 85.320 239.720 85.490 ;
        RECT 239.980 85.430 240.255 85.600 ;
        RECT 240.440 85.430 240.735 85.600 ;
        RECT 239.985 85.330 240.255 85.430 ;
        RECT 240.445 85.330 240.735 85.430 ;
        RECT 240.905 85.325 241.325 85.990 ;
        RECT 241.635 85.660 241.985 85.990 ;
        RECT 238.545 84.965 238.880 85.225 ;
        RECT 239.550 85.150 239.720 85.320 ;
        RECT 239.050 84.750 239.380 85.150 ;
        RECT 239.550 84.980 241.165 85.150 ;
        RECT 241.710 84.750 242.040 85.470 ;
        RECT 242.280 85.430 242.635 85.990 ;
        RECT 242.805 85.260 242.975 86.160 ;
        RECT 243.145 85.430 243.410 85.990 ;
        RECT 243.660 85.660 243.830 86.160 ;
        RECT 244.000 85.490 244.315 86.510 ;
        RECT 242.385 84.750 242.625 85.260 ;
        RECT 242.805 84.930 243.085 85.260 ;
        RECT 243.315 84.750 243.530 85.260 ;
        RECT 243.700 84.920 244.315 85.490 ;
        RECT 246.105 85.295 246.445 86.125 ;
        RECT 247.925 85.615 248.275 86.865 ;
        RECT 250.040 86.210 251.710 87.300 ;
        RECT 250.040 85.520 250.790 86.040 ;
        RECT 250.960 85.690 251.710 86.210 ;
        RECT 252.340 86.135 252.630 87.300 ;
        RECT 252.800 86.210 255.390 87.300 ;
        RECT 252.800 85.520 254.010 86.040 ;
        RECT 254.180 85.690 255.390 86.210 ;
        RECT 256.060 86.350 256.350 87.120 ;
        RECT 256.920 86.760 257.180 87.120 ;
        RECT 257.350 86.930 257.680 87.300 ;
        RECT 257.850 86.760 258.110 87.120 ;
        RECT 256.920 86.530 258.110 86.760 ;
        RECT 258.300 86.580 258.630 87.300 ;
        RECT 258.800 86.350 259.065 87.120 ;
        RECT 256.060 86.170 258.555 86.350 ;
        RECT 256.030 85.660 256.300 85.990 ;
        RECT 256.480 85.660 256.915 85.990 ;
        RECT 257.095 85.660 257.670 85.990 ;
        RECT 257.850 85.660 258.130 85.990 ;
        RECT 244.520 84.750 249.865 85.295 ;
        RECT 250.040 84.750 251.710 85.520 ;
        RECT 252.340 84.750 252.630 85.475 ;
        RECT 252.800 84.750 255.390 85.520 ;
        RECT 258.330 85.480 258.555 86.170 ;
        RECT 256.070 85.290 258.555 85.480 ;
        RECT 256.070 84.930 256.295 85.290 ;
        RECT 256.475 84.750 256.805 85.120 ;
        RECT 256.985 84.930 257.240 85.290 ;
        RECT 257.805 84.750 258.550 85.120 ;
        RECT 258.730 84.930 259.065 86.350 ;
        RECT 259.855 86.290 260.155 87.130 ;
        RECT 260.350 86.460 260.600 87.300 ;
        RECT 261.190 86.710 261.995 87.130 ;
        RECT 260.770 86.540 262.335 86.710 ;
        RECT 260.770 86.290 260.940 86.540 ;
        RECT 259.855 86.120 260.940 86.290 ;
        RECT 259.700 85.660 260.030 85.950 ;
        RECT 260.200 85.490 260.370 86.120 ;
        RECT 261.110 85.990 261.430 86.370 ;
        RECT 261.620 86.280 261.995 86.370 ;
        RECT 261.600 86.110 261.995 86.280 ;
        RECT 262.165 86.290 262.335 86.540 ;
        RECT 262.505 86.460 262.835 87.300 ;
        RECT 263.005 86.540 263.670 87.130 ;
        RECT 262.165 86.120 263.085 86.290 ;
        RECT 260.540 85.740 260.870 85.950 ;
        RECT 261.050 85.740 261.430 85.990 ;
        RECT 261.620 85.950 261.995 86.110 ;
        RECT 262.915 85.950 263.085 86.120 ;
        RECT 261.620 85.740 262.105 85.950 ;
        RECT 262.295 85.740 262.745 85.950 ;
        RECT 262.915 85.740 263.250 85.950 ;
        RECT 263.420 85.570 263.670 86.540 ;
        RECT 263.995 86.290 264.295 87.130 ;
        RECT 264.490 86.460 264.740 87.300 ;
        RECT 265.330 86.710 266.135 87.130 ;
        RECT 264.910 86.540 266.475 86.710 ;
        RECT 264.910 86.290 265.080 86.540 ;
        RECT 263.995 86.120 265.080 86.290 ;
        RECT 263.840 85.660 264.170 85.950 ;
        RECT 259.860 85.310 260.370 85.490 ;
        RECT 260.775 85.400 262.475 85.570 ;
        RECT 260.775 85.310 261.160 85.400 ;
        RECT 259.860 84.920 260.190 85.310 ;
        RECT 260.360 84.970 261.545 85.140 ;
        RECT 261.805 84.750 261.975 85.220 ;
        RECT 262.145 84.935 262.475 85.400 ;
        RECT 262.645 84.750 262.815 85.570 ;
        RECT 262.985 84.930 263.670 85.570 ;
        RECT 264.340 85.490 264.510 86.120 ;
        RECT 265.250 85.990 265.570 86.370 ;
        RECT 265.760 86.280 266.135 86.370 ;
        RECT 265.740 86.110 266.135 86.280 ;
        RECT 266.305 86.290 266.475 86.540 ;
        RECT 266.645 86.460 266.975 87.300 ;
        RECT 267.145 86.540 267.810 87.130 ;
        RECT 266.305 86.120 267.225 86.290 ;
        RECT 264.680 85.740 265.010 85.950 ;
        RECT 265.190 85.740 265.570 85.990 ;
        RECT 265.760 85.950 266.135 86.110 ;
        RECT 267.055 85.950 267.225 86.120 ;
        RECT 265.760 85.740 266.245 85.950 ;
        RECT 266.435 85.740 266.885 85.950 ;
        RECT 267.055 85.740 267.390 85.950 ;
        RECT 267.560 85.570 267.810 86.540 ;
        RECT 268.185 86.330 268.515 87.130 ;
        RECT 268.685 86.500 269.015 87.300 ;
        RECT 269.315 86.330 269.645 87.130 ;
        RECT 270.290 86.500 270.540 87.300 ;
        RECT 268.185 86.160 270.620 86.330 ;
        RECT 270.810 86.160 270.980 87.300 ;
        RECT 271.150 86.160 271.490 87.130 ;
        RECT 271.660 86.865 277.005 87.300 ;
        RECT 267.980 85.740 268.330 85.990 ;
        RECT 264.000 85.310 264.510 85.490 ;
        RECT 264.915 85.400 266.615 85.570 ;
        RECT 264.915 85.310 265.300 85.400 ;
        RECT 264.000 84.920 264.330 85.310 ;
        RECT 264.500 84.970 265.685 85.140 ;
        RECT 265.945 84.750 266.115 85.220 ;
        RECT 266.285 84.935 266.615 85.400 ;
        RECT 266.785 84.750 266.955 85.570 ;
        RECT 267.125 84.930 267.810 85.570 ;
        RECT 268.515 85.530 268.685 86.160 ;
        RECT 268.855 85.740 269.185 85.940 ;
        RECT 269.355 85.740 269.685 85.940 ;
        RECT 269.855 85.740 270.275 85.940 ;
        RECT 270.450 85.910 270.620 86.160 ;
        RECT 270.450 85.740 271.145 85.910 ;
        RECT 268.185 84.920 268.685 85.530 ;
        RECT 269.315 85.400 270.540 85.570 ;
        RECT 271.315 85.550 271.490 86.160 ;
        RECT 269.315 84.920 269.645 85.400 ;
        RECT 269.815 84.750 270.040 85.210 ;
        RECT 270.210 84.920 270.540 85.400 ;
        RECT 270.730 84.750 270.980 85.550 ;
        RECT 271.150 84.920 271.490 85.550 ;
        RECT 273.245 85.295 273.585 86.125 ;
        RECT 275.065 85.615 275.415 86.865 ;
        RECT 278.100 86.135 278.390 87.300 ;
        RECT 278.570 86.580 278.900 87.300 ;
        RECT 278.560 85.940 278.790 86.280 ;
        RECT 279.080 85.940 279.295 87.055 ;
        RECT 279.490 86.355 279.820 87.130 ;
        RECT 279.990 86.525 280.700 87.300 ;
        RECT 279.490 86.140 280.640 86.355 ;
        RECT 278.560 85.740 278.890 85.940 ;
        RECT 279.080 85.760 279.530 85.940 ;
        RECT 279.200 85.740 279.530 85.760 ;
        RECT 279.700 85.740 280.170 85.970 ;
        RECT 280.355 85.570 280.640 86.140 ;
        RECT 280.870 85.695 281.150 87.130 ;
        RECT 281.320 86.210 282.990 87.300 ;
        RECT 283.165 86.630 283.420 87.130 ;
        RECT 283.590 86.800 283.920 87.300 ;
        RECT 283.165 86.460 283.915 86.630 ;
        RECT 271.660 84.750 277.005 85.295 ;
        RECT 278.100 84.750 278.390 85.475 ;
        RECT 278.560 85.380 279.740 85.570 ;
        RECT 278.560 84.920 278.900 85.380 ;
        RECT 279.410 85.300 279.740 85.380 ;
        RECT 279.930 85.380 280.640 85.570 ;
        RECT 279.930 85.240 280.230 85.380 ;
        RECT 279.915 85.230 280.230 85.240 ;
        RECT 279.905 85.220 280.230 85.230 ;
        RECT 279.895 85.215 280.230 85.220 ;
        RECT 279.070 84.750 279.240 85.210 ;
        RECT 279.890 85.205 280.230 85.215 ;
        RECT 279.885 85.200 280.230 85.205 ;
        RECT 279.880 85.190 280.230 85.200 ;
        RECT 279.875 85.185 280.230 85.190 ;
        RECT 279.870 84.920 280.230 85.185 ;
        RECT 280.470 84.750 280.640 85.210 ;
        RECT 280.810 84.920 281.150 85.695 ;
        RECT 281.320 85.520 282.070 86.040 ;
        RECT 282.240 85.690 282.990 86.210 ;
        RECT 283.165 85.640 283.515 86.290 ;
        RECT 281.320 84.750 282.990 85.520 ;
        RECT 283.685 85.470 283.915 86.460 ;
        RECT 283.165 85.300 283.915 85.470 ;
        RECT 283.165 85.010 283.420 85.300 ;
        RECT 283.590 84.750 283.920 85.130 ;
        RECT 284.090 85.010 284.260 87.130 ;
        RECT 284.430 86.330 284.755 87.115 ;
        RECT 284.925 86.840 285.175 87.300 ;
        RECT 285.345 86.800 285.595 87.130 ;
        RECT 285.810 86.800 286.490 87.130 ;
        RECT 285.345 86.670 285.515 86.800 ;
        RECT 285.120 86.500 285.515 86.670 ;
        RECT 284.490 85.280 284.950 86.330 ;
        RECT 285.120 85.140 285.290 86.500 ;
        RECT 285.685 86.240 286.150 86.630 ;
        RECT 285.460 85.430 285.810 86.050 ;
        RECT 285.980 85.650 286.150 86.240 ;
        RECT 286.320 86.020 286.490 86.800 ;
        RECT 286.660 86.700 286.830 87.040 ;
        RECT 287.065 86.870 287.395 87.300 ;
        RECT 287.565 86.700 287.735 87.040 ;
        RECT 288.030 86.840 288.400 87.300 ;
        RECT 286.660 86.530 287.735 86.700 ;
        RECT 288.570 86.670 288.740 87.130 ;
        RECT 288.975 86.790 289.845 87.130 ;
        RECT 290.015 86.840 290.265 87.300 ;
        RECT 288.180 86.500 288.740 86.670 ;
        RECT 288.180 86.360 288.350 86.500 ;
        RECT 286.850 86.190 288.350 86.360 ;
        RECT 289.045 86.330 289.505 86.620 ;
        RECT 286.320 85.850 288.010 86.020 ;
        RECT 285.980 85.430 286.335 85.650 ;
        RECT 286.505 85.140 286.675 85.850 ;
        RECT 286.880 85.430 287.670 85.680 ;
        RECT 287.840 85.670 288.010 85.850 ;
        RECT 288.180 85.500 288.350 86.190 ;
        RECT 284.620 84.750 284.950 85.110 ;
        RECT 285.120 84.970 285.615 85.140 ;
        RECT 285.820 84.970 286.675 85.140 ;
        RECT 287.550 84.750 287.880 85.210 ;
        RECT 288.090 85.110 288.350 85.500 ;
        RECT 288.540 86.320 289.505 86.330 ;
        RECT 289.675 86.410 289.845 86.790 ;
        RECT 290.435 86.750 290.605 87.040 ;
        RECT 290.785 86.920 291.115 87.300 ;
        RECT 290.435 86.580 291.235 86.750 ;
        RECT 288.540 86.160 289.215 86.320 ;
        RECT 289.675 86.240 290.895 86.410 ;
        RECT 288.540 85.370 288.750 86.160 ;
        RECT 289.675 86.150 289.845 86.240 ;
        RECT 288.920 85.370 289.270 85.990 ;
        RECT 289.440 85.980 289.845 86.150 ;
        RECT 289.440 85.200 289.610 85.980 ;
        RECT 289.780 85.530 290.000 85.810 ;
        RECT 290.180 85.700 290.720 86.070 ;
        RECT 291.065 85.990 291.235 86.580 ;
        RECT 291.455 86.160 291.760 87.300 ;
        RECT 291.930 86.110 292.180 86.990 ;
        RECT 292.350 86.160 292.600 87.300 ;
        RECT 293.370 86.370 293.540 87.130 ;
        RECT 293.720 86.540 294.050 87.300 ;
        RECT 293.370 86.200 294.035 86.370 ;
        RECT 294.220 86.225 294.490 87.130 ;
        RECT 291.065 85.960 291.805 85.990 ;
        RECT 289.780 85.360 290.310 85.530 ;
        RECT 288.090 84.940 288.440 85.110 ;
        RECT 288.660 84.920 289.610 85.200 ;
        RECT 289.780 84.750 289.970 85.190 ;
        RECT 290.140 85.130 290.310 85.360 ;
        RECT 290.480 85.300 290.720 85.700 ;
        RECT 290.890 85.660 291.805 85.960 ;
        RECT 290.890 85.485 291.215 85.660 ;
        RECT 290.890 85.130 291.210 85.485 ;
        RECT 291.975 85.460 292.180 86.110 ;
        RECT 293.865 86.055 294.035 86.200 ;
        RECT 293.300 85.650 293.630 86.020 ;
        RECT 293.865 85.725 294.150 86.055 ;
        RECT 290.140 84.960 291.210 85.130 ;
        RECT 291.455 84.750 291.760 85.210 ;
        RECT 291.930 84.930 292.180 85.460 ;
        RECT 292.350 84.750 292.600 85.505 ;
        RECT 293.865 85.470 294.035 85.725 ;
        RECT 293.370 85.300 294.035 85.470 ;
        RECT 294.320 85.425 294.490 86.225 ;
        RECT 295.120 86.540 295.635 86.950 ;
        RECT 295.870 86.540 296.040 87.300 ;
        RECT 296.210 86.960 298.240 87.130 ;
        RECT 295.120 85.730 295.460 86.540 ;
        RECT 296.210 86.295 296.380 86.960 ;
        RECT 296.775 86.620 297.900 86.790 ;
        RECT 295.630 86.105 296.380 86.295 ;
        RECT 296.550 86.280 297.560 86.450 ;
        RECT 295.120 85.560 296.350 85.730 ;
        RECT 293.370 84.920 293.540 85.300 ;
        RECT 293.720 84.750 294.050 85.130 ;
        RECT 294.230 84.920 294.490 85.425 ;
        RECT 295.395 84.955 295.640 85.560 ;
        RECT 295.860 84.750 296.370 85.285 ;
        RECT 296.550 84.920 296.740 86.280 ;
        RECT 296.910 85.940 297.185 86.080 ;
        RECT 296.910 85.770 297.190 85.940 ;
        RECT 296.910 84.920 297.185 85.770 ;
        RECT 297.390 85.480 297.560 86.280 ;
        RECT 297.730 85.490 297.900 86.620 ;
        RECT 298.070 85.990 298.240 86.960 ;
        RECT 298.410 86.160 298.580 87.300 ;
        RECT 298.750 86.160 299.085 87.130 ;
        RECT 299.350 86.370 299.520 87.130 ;
        RECT 299.700 86.540 300.030 87.300 ;
        RECT 299.350 86.200 300.015 86.370 ;
        RECT 300.200 86.225 300.470 87.130 ;
        RECT 298.070 85.660 298.265 85.990 ;
        RECT 298.490 85.660 298.745 85.990 ;
        RECT 298.490 85.490 298.660 85.660 ;
        RECT 298.915 85.490 299.085 86.160 ;
        RECT 299.845 86.055 300.015 86.200 ;
        RECT 299.280 85.650 299.610 86.020 ;
        RECT 299.845 85.725 300.130 86.055 ;
        RECT 297.730 85.320 298.660 85.490 ;
        RECT 297.730 85.285 297.905 85.320 ;
        RECT 297.375 84.920 297.905 85.285 ;
        RECT 298.330 84.750 298.660 85.150 ;
        RECT 298.830 84.920 299.085 85.490 ;
        RECT 299.845 85.470 300.015 85.725 ;
        RECT 299.350 85.300 300.015 85.470 ;
        RECT 300.300 85.425 300.470 86.225 ;
        RECT 300.640 86.210 303.230 87.300 ;
        RECT 299.350 84.920 299.520 85.300 ;
        RECT 299.700 84.750 300.030 85.130 ;
        RECT 300.210 84.920 300.470 85.425 ;
        RECT 300.640 85.520 301.850 86.040 ;
        RECT 302.020 85.690 303.230 86.210 ;
        RECT 303.860 86.135 304.150 87.300 ;
        RECT 304.320 86.210 307.830 87.300 ;
        RECT 304.320 85.520 305.970 86.040 ;
        RECT 306.140 85.690 307.830 86.210 ;
        RECT 308.460 86.225 308.730 87.130 ;
        RECT 308.900 86.540 309.230 87.300 ;
        RECT 309.410 86.370 309.580 87.130 ;
        RECT 300.640 84.750 303.230 85.520 ;
        RECT 303.860 84.750 304.150 85.475 ;
        RECT 304.320 84.750 307.830 85.520 ;
        RECT 308.460 85.425 308.630 86.225 ;
        RECT 308.915 86.200 309.580 86.370 ;
        RECT 309.840 86.210 311.050 87.300 ;
        RECT 308.915 86.055 309.085 86.200 ;
        RECT 308.800 85.725 309.085 86.055 ;
        RECT 308.915 85.470 309.085 85.725 ;
        RECT 309.320 85.650 309.650 86.020 ;
        RECT 309.840 85.670 310.360 86.210 ;
        RECT 310.530 85.500 311.050 86.040 ;
        RECT 308.460 84.920 308.720 85.425 ;
        RECT 308.915 85.300 309.580 85.470 ;
        RECT 308.900 84.750 309.230 85.130 ;
        RECT 309.410 84.920 309.580 85.300 ;
        RECT 309.840 84.750 311.050 85.500 ;
        RECT 162.095 84.580 311.135 84.750 ;
        RECT 162.180 83.830 163.390 84.580 ;
        RECT 163.560 84.035 168.905 84.580 ;
        RECT 169.080 84.035 174.425 84.580 ;
        RECT 162.180 83.290 162.700 83.830 ;
        RECT 162.870 83.120 163.390 83.660 ;
        RECT 165.145 83.205 165.485 84.035 ;
        RECT 162.180 82.030 163.390 83.120 ;
        RECT 166.965 82.465 167.315 83.715 ;
        RECT 170.665 83.205 171.005 84.035 ;
        RECT 174.600 83.810 178.110 84.580 ;
        RECT 178.330 83.825 178.580 84.580 ;
        RECT 178.750 83.870 179.000 84.400 ;
        RECT 179.170 84.120 179.475 84.580 ;
        RECT 179.720 84.200 180.790 84.370 ;
        RECT 172.485 82.465 172.835 83.715 ;
        RECT 174.600 83.290 176.250 83.810 ;
        RECT 176.420 83.120 178.110 83.640 ;
        RECT 178.750 83.220 178.955 83.870 ;
        RECT 179.720 83.845 180.040 84.200 ;
        RECT 179.715 83.670 180.040 83.845 ;
        RECT 179.125 83.370 180.040 83.670 ;
        RECT 180.210 83.630 180.450 84.030 ;
        RECT 180.620 83.970 180.790 84.200 ;
        RECT 180.960 84.140 181.150 84.580 ;
        RECT 181.320 84.130 182.270 84.410 ;
        RECT 182.490 84.220 182.840 84.390 ;
        RECT 180.620 83.800 181.150 83.970 ;
        RECT 179.125 83.340 179.865 83.370 ;
        RECT 163.560 82.030 168.905 82.465 ;
        RECT 169.080 82.030 174.425 82.465 ;
        RECT 174.600 82.030 178.110 83.120 ;
        RECT 178.330 82.030 178.580 83.170 ;
        RECT 178.750 82.340 179.000 83.220 ;
        RECT 179.170 82.030 179.475 83.170 ;
        RECT 179.695 82.750 179.865 83.340 ;
        RECT 180.210 83.260 180.750 83.630 ;
        RECT 180.930 83.520 181.150 83.800 ;
        RECT 181.320 83.350 181.490 84.130 ;
        RECT 181.085 83.180 181.490 83.350 ;
        RECT 181.660 83.340 182.010 83.960 ;
        RECT 181.085 83.090 181.255 83.180 ;
        RECT 182.180 83.170 182.390 83.960 ;
        RECT 180.035 82.920 181.255 83.090 ;
        RECT 181.715 83.010 182.390 83.170 ;
        RECT 179.695 82.580 180.495 82.750 ;
        RECT 179.815 82.030 180.145 82.410 ;
        RECT 180.325 82.290 180.495 82.580 ;
        RECT 181.085 82.540 181.255 82.920 ;
        RECT 181.425 83.000 182.390 83.010 ;
        RECT 182.580 83.830 182.840 84.220 ;
        RECT 183.050 84.120 183.380 84.580 ;
        RECT 184.255 84.190 185.110 84.360 ;
        RECT 185.315 84.190 185.810 84.360 ;
        RECT 185.980 84.220 186.310 84.580 ;
        RECT 182.580 83.140 182.750 83.830 ;
        RECT 182.920 83.480 183.090 83.660 ;
        RECT 183.260 83.650 184.050 83.900 ;
        RECT 184.255 83.480 184.425 84.190 ;
        RECT 184.595 83.680 184.950 83.900 ;
        RECT 182.920 83.310 184.610 83.480 ;
        RECT 181.425 82.710 181.885 83.000 ;
        RECT 182.580 82.970 184.080 83.140 ;
        RECT 182.580 82.830 182.750 82.970 ;
        RECT 182.190 82.660 182.750 82.830 ;
        RECT 180.665 82.030 180.915 82.490 ;
        RECT 181.085 82.200 181.955 82.540 ;
        RECT 182.190 82.200 182.360 82.660 ;
        RECT 183.195 82.630 184.270 82.800 ;
        RECT 182.530 82.030 182.900 82.490 ;
        RECT 183.195 82.290 183.365 82.630 ;
        RECT 183.535 82.030 183.865 82.460 ;
        RECT 184.100 82.290 184.270 82.630 ;
        RECT 184.440 82.530 184.610 83.310 ;
        RECT 184.780 83.090 184.950 83.680 ;
        RECT 185.120 83.280 185.470 83.900 ;
        RECT 184.780 82.700 185.245 83.090 ;
        RECT 185.640 82.830 185.810 84.190 ;
        RECT 185.980 83.000 186.440 84.050 ;
        RECT 185.415 82.660 185.810 82.830 ;
        RECT 185.415 82.530 185.585 82.660 ;
        RECT 184.440 82.200 185.120 82.530 ;
        RECT 185.335 82.200 185.585 82.530 ;
        RECT 185.755 82.030 186.005 82.490 ;
        RECT 186.175 82.215 186.500 83.000 ;
        RECT 186.670 82.200 186.840 84.320 ;
        RECT 187.010 84.200 187.340 84.580 ;
        RECT 187.510 84.030 187.765 84.320 ;
        RECT 187.015 83.860 187.765 84.030 ;
        RECT 187.015 82.870 187.245 83.860 ;
        RECT 187.940 83.855 188.230 84.580 ;
        RECT 189.320 83.905 189.580 84.410 ;
        RECT 189.760 84.200 190.090 84.580 ;
        RECT 190.270 84.030 190.440 84.410 ;
        RECT 191.865 84.100 192.165 84.580 ;
        RECT 187.415 83.040 187.765 83.690 ;
        RECT 187.015 82.700 187.765 82.870 ;
        RECT 187.010 82.030 187.340 82.530 ;
        RECT 187.510 82.200 187.765 82.700 ;
        RECT 187.940 82.030 188.230 83.195 ;
        RECT 189.320 83.105 189.490 83.905 ;
        RECT 189.775 83.860 190.440 84.030 ;
        RECT 192.335 83.930 192.595 84.385 ;
        RECT 192.765 84.100 193.025 84.580 ;
        RECT 193.195 83.930 193.455 84.385 ;
        RECT 193.625 84.100 193.885 84.580 ;
        RECT 194.055 83.930 194.315 84.385 ;
        RECT 194.485 84.100 194.745 84.580 ;
        RECT 194.915 83.930 195.175 84.385 ;
        RECT 195.345 84.055 195.605 84.580 ;
        RECT 189.775 83.605 189.945 83.860 ;
        RECT 191.865 83.760 195.175 83.930 ;
        RECT 189.660 83.275 189.945 83.605 ;
        RECT 190.180 83.310 190.510 83.680 ;
        RECT 189.775 83.130 189.945 83.275 ;
        RECT 191.865 83.170 192.835 83.760 ;
        RECT 195.775 83.590 196.025 84.400 ;
        RECT 196.205 84.120 196.450 84.580 ;
        RECT 193.005 83.340 196.025 83.590 ;
        RECT 196.195 83.340 196.510 83.950 ;
        RECT 196.680 83.810 200.190 84.580 ;
        RECT 200.360 83.830 201.570 84.580 ;
        RECT 201.800 84.120 202.045 84.580 ;
        RECT 189.320 82.200 189.590 83.105 ;
        RECT 189.775 82.960 190.440 83.130 ;
        RECT 189.760 82.030 190.090 82.790 ;
        RECT 190.270 82.200 190.440 82.960 ;
        RECT 191.865 82.930 195.175 83.170 ;
        RECT 191.870 82.030 192.165 82.760 ;
        RECT 192.335 82.205 192.595 82.930 ;
        RECT 192.765 82.030 193.025 82.760 ;
        RECT 193.195 82.205 193.455 82.930 ;
        RECT 193.625 82.030 193.885 82.760 ;
        RECT 194.055 82.205 194.315 82.930 ;
        RECT 194.485 82.030 194.745 82.760 ;
        RECT 194.915 82.205 195.175 82.930 ;
        RECT 195.345 82.030 195.605 83.140 ;
        RECT 195.775 82.205 196.025 83.340 ;
        RECT 196.680 83.290 198.330 83.810 ;
        RECT 196.205 82.030 196.500 83.140 ;
        RECT 198.500 83.120 200.190 83.640 ;
        RECT 200.360 83.290 200.880 83.830 ;
        RECT 201.050 83.120 201.570 83.660 ;
        RECT 201.740 83.340 202.055 83.950 ;
        RECT 202.225 83.590 202.475 84.400 ;
        RECT 202.645 84.055 202.905 84.580 ;
        RECT 203.075 83.930 203.335 84.385 ;
        RECT 203.505 84.100 203.765 84.580 ;
        RECT 203.935 83.930 204.195 84.385 ;
        RECT 204.365 84.100 204.625 84.580 ;
        RECT 204.795 83.930 205.055 84.385 ;
        RECT 205.225 84.100 205.485 84.580 ;
        RECT 205.655 83.930 205.915 84.385 ;
        RECT 206.085 84.100 206.385 84.580 ;
        RECT 203.075 83.760 206.385 83.930 ;
        RECT 207.260 83.780 207.550 84.580 ;
        RECT 207.720 84.120 208.270 84.410 ;
        RECT 208.440 84.120 208.690 84.580 ;
        RECT 202.225 83.340 205.245 83.590 ;
        RECT 196.680 82.030 200.190 83.120 ;
        RECT 200.360 82.030 201.570 83.120 ;
        RECT 201.750 82.030 202.045 83.140 ;
        RECT 202.225 82.205 202.475 83.340 ;
        RECT 205.415 83.170 206.385 83.760 ;
        RECT 202.645 82.030 202.905 83.140 ;
        RECT 203.075 82.930 206.385 83.170 ;
        RECT 203.075 82.205 203.335 82.930 ;
        RECT 203.505 82.030 203.765 82.760 ;
        RECT 203.935 82.205 204.195 82.930 ;
        RECT 204.365 82.030 204.625 82.760 ;
        RECT 204.795 82.205 205.055 82.930 ;
        RECT 205.225 82.030 205.485 82.760 ;
        RECT 205.655 82.205 205.915 82.930 ;
        RECT 206.085 82.030 206.380 82.760 ;
        RECT 207.260 82.030 207.550 83.170 ;
        RECT 207.720 82.750 207.970 84.120 ;
        RECT 209.320 83.950 209.650 84.310 ;
        RECT 208.260 83.760 209.650 83.950 ;
        RECT 210.480 83.780 210.770 84.580 ;
        RECT 210.940 84.120 211.490 84.410 ;
        RECT 211.660 84.120 211.910 84.580 ;
        RECT 208.260 83.670 208.430 83.760 ;
        RECT 208.140 83.340 208.430 83.670 ;
        RECT 208.600 83.340 208.930 83.590 ;
        RECT 209.160 83.340 209.850 83.590 ;
        RECT 208.260 83.090 208.430 83.340 ;
        RECT 208.260 82.920 209.200 83.090 ;
        RECT 207.720 82.200 208.170 82.750 ;
        RECT 208.360 82.030 208.690 82.750 ;
        RECT 208.900 82.370 209.200 82.920 ;
        RECT 209.535 82.900 209.850 83.340 ;
        RECT 209.370 82.030 209.650 82.700 ;
        RECT 210.480 82.030 210.770 83.170 ;
        RECT 210.940 82.750 211.190 84.120 ;
        RECT 212.540 83.950 212.870 84.310 ;
        RECT 211.480 83.760 212.870 83.950 ;
        RECT 213.700 83.855 213.990 84.580 ;
        RECT 214.160 84.035 219.505 84.580 ;
        RECT 211.480 83.670 211.650 83.760 ;
        RECT 211.360 83.340 211.650 83.670 ;
        RECT 211.820 83.340 212.150 83.590 ;
        RECT 212.380 83.340 213.070 83.590 ;
        RECT 211.480 83.090 211.650 83.340 ;
        RECT 211.480 82.920 212.420 83.090 ;
        RECT 210.940 82.200 211.390 82.750 ;
        RECT 211.580 82.030 211.910 82.750 ;
        RECT 212.120 82.370 212.420 82.920 ;
        RECT 212.755 82.900 213.070 83.340 ;
        RECT 215.745 83.205 216.085 84.035 ;
        RECT 220.165 83.930 220.500 84.410 ;
        RECT 220.670 84.110 220.840 84.580 ;
        RECT 221.010 83.940 221.340 84.410 ;
        RECT 221.510 84.110 221.680 84.580 ;
        RECT 221.850 83.940 222.180 84.410 ;
        RECT 222.350 84.110 223.040 84.580 ;
        RECT 223.210 83.940 223.540 84.410 ;
        RECT 223.710 84.110 223.880 84.580 ;
        RECT 224.050 83.940 224.380 84.410 ;
        RECT 224.550 84.110 224.720 84.580 ;
        RECT 224.890 83.940 225.220 84.410 ;
        RECT 225.390 84.110 225.560 84.580 ;
        RECT 225.730 83.940 226.060 84.410 ;
        RECT 226.230 84.110 226.400 84.580 ;
        RECT 226.570 83.940 226.815 84.350 ;
        RECT 227.060 84.095 227.850 84.360 ;
        RECT 220.165 83.760 220.840 83.930 ;
        RECT 221.010 83.760 226.815 83.940 ;
        RECT 212.590 82.030 212.870 82.700 ;
        RECT 213.700 82.030 213.990 83.195 ;
        RECT 217.565 82.465 217.915 83.715 ;
        RECT 220.165 83.380 220.500 83.590 ;
        RECT 220.670 83.210 220.840 83.760 ;
        RECT 221.090 83.380 222.745 83.590 ;
        RECT 223.090 83.380 224.355 83.590 ;
        RECT 224.590 83.380 226.180 83.590 ;
        RECT 224.590 83.210 224.760 83.380 ;
        RECT 226.475 83.210 226.815 83.760 ;
        RECT 227.040 83.420 227.425 83.900 ;
        RECT 227.595 83.240 227.850 84.095 ;
        RECT 228.020 83.915 228.250 84.360 ;
        RECT 228.430 84.085 228.760 84.580 ;
        RECT 228.935 83.950 229.185 84.410 ;
        RECT 228.020 83.420 228.430 83.915 ;
        RECT 229.015 83.740 229.185 83.950 ;
        RECT 229.355 83.920 229.630 84.580 ;
        RECT 229.800 84.080 230.100 84.410 ;
        RECT 230.270 84.100 230.545 84.580 ;
        RECT 228.615 83.240 228.845 83.670 ;
        RECT 220.165 83.040 224.760 83.210 ;
        RECT 224.930 83.040 226.815 83.210 ;
        RECT 214.160 82.030 219.505 82.465 ;
        RECT 220.165 82.200 220.460 83.040 ;
        RECT 220.630 82.030 220.880 82.870 ;
        RECT 221.050 82.700 224.340 82.870 ;
        RECT 221.050 82.200 221.300 82.700 ;
        RECT 221.470 82.030 221.720 82.530 ;
        RECT 221.890 82.200 222.140 82.700 ;
        RECT 223.250 82.540 223.500 82.700 ;
        RECT 224.090 82.540 224.340 82.700 ;
        RECT 222.310 82.030 222.560 82.530 ;
        RECT 222.830 82.370 223.080 82.530 ;
        RECT 223.670 82.370 223.920 82.530 ;
        RECT 224.510 82.370 224.760 82.870 ;
        RECT 224.930 82.540 225.180 83.040 ;
        RECT 225.350 82.370 225.600 82.870 ;
        RECT 225.770 82.540 226.020 83.040 ;
        RECT 226.190 82.370 226.440 82.870 ;
        RECT 222.830 82.200 226.440 82.370 ;
        RECT 226.610 82.250 226.815 83.040 ;
        RECT 227.055 83.070 228.845 83.240 ;
        RECT 229.015 83.220 229.630 83.740 ;
        RECT 227.055 82.705 227.310 83.070 ;
        RECT 227.480 82.710 227.810 82.900 ;
        RECT 228.035 82.775 228.285 83.070 ;
        RECT 229.030 82.880 229.200 83.220 ;
        RECT 229.800 83.170 229.970 84.080 ;
        RECT 230.725 83.930 231.020 84.320 ;
        RECT 231.190 84.100 231.445 84.580 ;
        RECT 231.620 83.930 231.880 84.320 ;
        RECT 232.050 84.100 232.330 84.580 ;
        RECT 232.560 84.035 237.905 84.580 ;
        RECT 230.140 83.340 230.490 83.910 ;
        RECT 230.725 83.760 232.375 83.930 ;
        RECT 230.660 83.420 231.800 83.590 ;
        RECT 230.660 83.170 230.830 83.420 ;
        RECT 231.970 83.250 232.375 83.760 ;
        RECT 227.480 82.535 227.670 82.710 ;
        RECT 227.040 82.030 227.670 82.535 ;
        RECT 227.850 82.200 228.325 82.540 ;
        RECT 228.510 82.030 228.725 82.875 ;
        RECT 228.940 82.870 229.200 82.880 ;
        RECT 228.925 82.200 229.200 82.870 ;
        RECT 229.370 82.030 229.630 83.040 ;
        RECT 229.800 83.000 230.830 83.170 ;
        RECT 231.620 83.080 232.375 83.250 ;
        RECT 234.145 83.205 234.485 84.035 ;
        RECT 238.080 83.830 239.290 84.580 ;
        RECT 239.460 83.855 239.750 84.580 ;
        RECT 229.800 82.200 230.110 83.000 ;
        RECT 231.620 82.830 231.880 83.080 ;
        RECT 230.280 82.030 230.590 82.830 ;
        RECT 230.760 82.660 231.880 82.830 ;
        RECT 230.760 82.200 231.020 82.660 ;
        RECT 231.190 82.030 231.445 82.490 ;
        RECT 231.620 82.200 231.880 82.660 ;
        RECT 232.050 82.030 232.335 82.900 ;
        RECT 235.965 82.465 236.315 83.715 ;
        RECT 238.080 83.290 238.600 83.830 ;
        RECT 239.920 83.810 241.590 84.580 ;
        RECT 242.310 83.930 242.480 84.410 ;
        RECT 242.650 84.100 242.980 84.580 ;
        RECT 243.205 84.160 244.740 84.410 ;
        RECT 243.205 83.930 243.375 84.160 ;
        RECT 238.770 83.120 239.290 83.660 ;
        RECT 239.920 83.290 240.670 83.810 ;
        RECT 242.310 83.760 243.375 83.930 ;
        RECT 232.560 82.030 237.905 82.465 ;
        RECT 238.080 82.030 239.290 83.120 ;
        RECT 239.460 82.030 239.750 83.195 ;
        RECT 240.840 83.120 241.590 83.640 ;
        RECT 243.555 83.590 243.835 83.990 ;
        RECT 242.225 83.380 242.575 83.590 ;
        RECT 242.745 83.390 243.190 83.590 ;
        RECT 243.360 83.390 243.835 83.590 ;
        RECT 244.105 83.590 244.390 83.990 ;
        RECT 244.570 83.930 244.740 84.160 ;
        RECT 244.910 84.100 245.240 84.580 ;
        RECT 245.455 84.080 245.710 84.410 ;
        RECT 245.500 84.070 245.710 84.080 ;
        RECT 245.525 84.000 245.710 84.070 ;
        RECT 244.570 83.760 245.370 83.930 ;
        RECT 244.105 83.390 244.435 83.590 ;
        RECT 244.605 83.390 244.970 83.590 ;
        RECT 245.200 83.210 245.370 83.760 ;
        RECT 239.920 82.030 241.590 83.120 ;
        RECT 242.310 83.040 245.370 83.210 ;
        RECT 242.310 82.200 242.480 83.040 ;
        RECT 245.540 82.870 245.710 84.000 ;
        RECT 242.650 82.370 242.980 82.870 ;
        RECT 243.150 82.630 244.785 82.870 ;
        RECT 243.150 82.540 243.380 82.630 ;
        RECT 243.490 82.370 243.820 82.410 ;
        RECT 242.650 82.200 243.820 82.370 ;
        RECT 244.010 82.030 244.365 82.450 ;
        RECT 244.535 82.200 244.785 82.630 ;
        RECT 244.955 82.030 245.285 82.790 ;
        RECT 245.455 82.200 245.710 82.870 ;
        RECT 245.910 83.855 246.240 84.365 ;
        RECT 246.410 84.180 246.740 84.580 ;
        RECT 247.790 84.010 248.120 84.350 ;
        RECT 248.290 84.180 248.620 84.580 ;
        RECT 249.120 84.035 254.465 84.580 ;
        RECT 254.640 84.035 259.985 84.580 ;
        RECT 245.910 83.090 246.100 83.855 ;
        RECT 246.410 83.840 248.775 84.010 ;
        RECT 246.410 83.670 246.580 83.840 ;
        RECT 246.270 83.340 246.580 83.670 ;
        RECT 246.750 83.340 247.055 83.670 ;
        RECT 245.910 82.240 246.240 83.090 ;
        RECT 246.410 82.030 246.660 83.170 ;
        RECT 246.840 83.010 247.055 83.340 ;
        RECT 247.230 83.010 247.515 83.670 ;
        RECT 247.710 83.010 247.975 83.670 ;
        RECT 248.190 83.010 248.435 83.670 ;
        RECT 248.605 82.840 248.775 83.840 ;
        RECT 250.705 83.205 251.045 84.035 ;
        RECT 246.850 82.670 248.140 82.840 ;
        RECT 246.850 82.250 247.100 82.670 ;
        RECT 247.330 82.030 247.660 82.500 ;
        RECT 247.890 82.250 248.140 82.670 ;
        RECT 248.320 82.670 248.775 82.840 ;
        RECT 248.320 82.240 248.650 82.670 ;
        RECT 252.525 82.465 252.875 83.715 ;
        RECT 256.225 83.205 256.565 84.035 ;
        RECT 260.160 83.810 261.830 84.580 ;
        RECT 262.330 84.180 262.660 84.580 ;
        RECT 262.830 84.010 263.160 84.350 ;
        RECT 264.210 84.180 264.540 84.580 ;
        RECT 262.175 83.840 264.540 84.010 ;
        RECT 264.710 83.855 265.040 84.365 ;
        RECT 265.220 83.855 265.510 84.580 ;
        RECT 265.845 84.070 266.085 84.580 ;
        RECT 266.265 84.070 266.545 84.400 ;
        RECT 266.775 84.070 266.990 84.580 ;
        RECT 258.045 82.465 258.395 83.715 ;
        RECT 260.160 83.290 260.910 83.810 ;
        RECT 261.080 83.120 261.830 83.640 ;
        RECT 249.120 82.030 254.465 82.465 ;
        RECT 254.640 82.030 259.985 82.465 ;
        RECT 260.160 82.030 261.830 83.120 ;
        RECT 262.175 82.840 262.345 83.840 ;
        RECT 264.370 83.670 264.540 83.840 ;
        RECT 262.515 83.010 262.760 83.670 ;
        RECT 262.975 83.010 263.240 83.670 ;
        RECT 263.435 83.010 263.720 83.670 ;
        RECT 263.895 83.340 264.200 83.670 ;
        RECT 264.370 83.340 264.680 83.670 ;
        RECT 263.895 83.010 264.110 83.340 ;
        RECT 262.175 82.670 262.630 82.840 ;
        RECT 262.300 82.240 262.630 82.670 ;
        RECT 262.810 82.670 264.100 82.840 ;
        RECT 262.810 82.250 263.060 82.670 ;
        RECT 263.290 82.030 263.620 82.500 ;
        RECT 263.850 82.250 264.100 82.670 ;
        RECT 264.290 82.030 264.540 83.170 ;
        RECT 264.850 83.090 265.040 83.855 ;
        RECT 265.740 83.340 266.095 83.900 ;
        RECT 264.710 82.240 265.040 83.090 ;
        RECT 265.220 82.030 265.510 83.195 ;
        RECT 266.265 83.170 266.435 84.070 ;
        RECT 266.605 83.340 266.870 83.900 ;
        RECT 267.160 83.840 267.775 84.410 ;
        RECT 267.120 83.170 267.290 83.670 ;
        RECT 265.865 83.000 267.290 83.170 ;
        RECT 265.865 82.825 266.255 83.000 ;
        RECT 266.740 82.030 267.070 82.830 ;
        RECT 267.460 82.820 267.775 83.840 ;
        RECT 267.980 83.810 271.490 84.580 ;
        RECT 271.660 83.830 272.870 84.580 ;
        RECT 273.045 84.030 273.300 84.320 ;
        RECT 273.470 84.200 273.800 84.580 ;
        RECT 273.045 83.860 273.795 84.030 ;
        RECT 267.980 83.290 269.630 83.810 ;
        RECT 269.800 83.120 271.490 83.640 ;
        RECT 271.660 83.290 272.180 83.830 ;
        RECT 272.350 83.120 272.870 83.660 ;
        RECT 267.240 82.200 267.775 82.820 ;
        RECT 267.980 82.030 271.490 83.120 ;
        RECT 271.660 82.030 272.870 83.120 ;
        RECT 273.045 83.040 273.395 83.690 ;
        RECT 273.565 82.870 273.795 83.860 ;
        RECT 273.045 82.700 273.795 82.870 ;
        RECT 273.045 82.200 273.300 82.700 ;
        RECT 273.470 82.030 273.800 82.530 ;
        RECT 273.970 82.200 274.140 84.320 ;
        RECT 274.500 84.220 274.830 84.580 ;
        RECT 275.000 84.190 275.495 84.360 ;
        RECT 275.700 84.190 276.555 84.360 ;
        RECT 274.370 83.000 274.830 84.050 ;
        RECT 274.310 82.215 274.635 83.000 ;
        RECT 275.000 82.830 275.170 84.190 ;
        RECT 275.340 83.280 275.690 83.900 ;
        RECT 275.860 83.680 276.215 83.900 ;
        RECT 275.860 83.090 276.030 83.680 ;
        RECT 276.385 83.480 276.555 84.190 ;
        RECT 277.430 84.120 277.760 84.580 ;
        RECT 277.970 84.220 278.320 84.390 ;
        RECT 276.760 83.650 277.550 83.900 ;
        RECT 277.970 83.830 278.230 84.220 ;
        RECT 278.540 84.130 279.490 84.410 ;
        RECT 279.660 84.140 279.850 84.580 ;
        RECT 280.020 84.200 281.090 84.370 ;
        RECT 277.720 83.480 277.890 83.660 ;
        RECT 275.000 82.660 275.395 82.830 ;
        RECT 275.565 82.700 276.030 83.090 ;
        RECT 276.200 83.310 277.890 83.480 ;
        RECT 275.225 82.530 275.395 82.660 ;
        RECT 276.200 82.530 276.370 83.310 ;
        RECT 278.060 83.140 278.230 83.830 ;
        RECT 276.730 82.970 278.230 83.140 ;
        RECT 278.420 83.170 278.630 83.960 ;
        RECT 278.800 83.340 279.150 83.960 ;
        RECT 279.320 83.350 279.490 84.130 ;
        RECT 280.020 83.970 280.190 84.200 ;
        RECT 279.660 83.800 280.190 83.970 ;
        RECT 279.660 83.520 279.880 83.800 ;
        RECT 280.360 83.630 280.600 84.030 ;
        RECT 279.320 83.180 279.725 83.350 ;
        RECT 280.060 83.260 280.600 83.630 ;
        RECT 280.770 83.845 281.090 84.200 ;
        RECT 281.335 84.120 281.640 84.580 ;
        RECT 281.810 83.870 282.065 84.400 ;
        RECT 282.300 84.120 282.545 84.580 ;
        RECT 280.770 83.670 281.095 83.845 ;
        RECT 280.770 83.370 281.685 83.670 ;
        RECT 280.945 83.340 281.685 83.370 ;
        RECT 278.420 83.010 279.095 83.170 ;
        RECT 279.555 83.090 279.725 83.180 ;
        RECT 278.420 83.000 279.385 83.010 ;
        RECT 278.060 82.830 278.230 82.970 ;
        RECT 274.805 82.030 275.055 82.490 ;
        RECT 275.225 82.200 275.475 82.530 ;
        RECT 275.690 82.200 276.370 82.530 ;
        RECT 276.540 82.630 277.615 82.800 ;
        RECT 278.060 82.660 278.620 82.830 ;
        RECT 278.925 82.710 279.385 83.000 ;
        RECT 279.555 82.920 280.775 83.090 ;
        RECT 276.540 82.290 276.710 82.630 ;
        RECT 276.945 82.030 277.275 82.460 ;
        RECT 277.445 82.290 277.615 82.630 ;
        RECT 277.910 82.030 278.280 82.490 ;
        RECT 278.450 82.200 278.620 82.660 ;
        RECT 279.555 82.540 279.725 82.920 ;
        RECT 280.945 82.750 281.115 83.340 ;
        RECT 281.855 83.220 282.065 83.870 ;
        RECT 282.240 83.340 282.555 83.950 ;
        RECT 282.725 83.590 282.975 84.400 ;
        RECT 283.145 84.055 283.405 84.580 ;
        RECT 283.575 83.930 283.835 84.385 ;
        RECT 284.005 84.100 284.265 84.580 ;
        RECT 284.435 83.930 284.695 84.385 ;
        RECT 284.865 84.100 285.125 84.580 ;
        RECT 285.295 83.930 285.555 84.385 ;
        RECT 285.725 84.100 285.985 84.580 ;
        RECT 286.155 83.930 286.415 84.385 ;
        RECT 286.585 84.100 286.885 84.580 ;
        RECT 283.575 83.760 286.885 83.930 ;
        RECT 282.725 83.340 285.745 83.590 ;
        RECT 278.855 82.200 279.725 82.540 ;
        RECT 280.315 82.580 281.115 82.750 ;
        RECT 279.895 82.030 280.145 82.490 ;
        RECT 280.315 82.290 280.485 82.580 ;
        RECT 280.665 82.030 280.995 82.410 ;
        RECT 281.335 82.030 281.640 83.170 ;
        RECT 281.810 82.340 282.065 83.220 ;
        RECT 282.250 82.030 282.545 83.140 ;
        RECT 282.725 82.205 282.975 83.340 ;
        RECT 285.915 83.170 286.885 83.760 ;
        RECT 283.145 82.030 283.405 83.140 ;
        RECT 283.575 82.930 286.885 83.170 ;
        RECT 287.300 83.905 287.560 84.410 ;
        RECT 287.740 84.200 288.070 84.580 ;
        RECT 288.250 84.030 288.420 84.410 ;
        RECT 287.300 83.105 287.470 83.905 ;
        RECT 287.755 83.860 288.420 84.030 ;
        RECT 287.755 83.605 287.925 83.860 ;
        RECT 288.680 83.810 290.350 84.580 ;
        RECT 290.980 83.855 291.270 84.580 ;
        RECT 292.420 84.100 292.700 84.580 ;
        RECT 292.870 83.930 293.130 84.320 ;
        RECT 293.305 84.100 293.560 84.580 ;
        RECT 293.730 83.930 294.025 84.320 ;
        RECT 294.205 84.100 294.480 84.580 ;
        RECT 294.650 84.080 294.950 84.410 ;
        RECT 287.640 83.275 287.925 83.605 ;
        RECT 288.160 83.310 288.490 83.680 ;
        RECT 288.680 83.290 289.430 83.810 ;
        RECT 292.375 83.760 294.025 83.930 ;
        RECT 287.755 83.130 287.925 83.275 ;
        RECT 283.575 82.205 283.835 82.930 ;
        RECT 284.005 82.030 284.265 82.760 ;
        RECT 284.435 82.205 284.695 82.930 ;
        RECT 284.865 82.030 285.125 82.760 ;
        RECT 285.295 82.205 285.555 82.930 ;
        RECT 285.725 82.030 285.985 82.760 ;
        RECT 286.155 82.205 286.415 82.930 ;
        RECT 286.585 82.030 286.880 82.760 ;
        RECT 287.300 82.200 287.570 83.105 ;
        RECT 287.755 82.960 288.420 83.130 ;
        RECT 289.600 83.120 290.350 83.640 ;
        RECT 292.375 83.250 292.780 83.760 ;
        RECT 292.950 83.420 294.090 83.590 ;
        RECT 287.740 82.030 288.070 82.790 ;
        RECT 288.250 82.200 288.420 82.960 ;
        RECT 288.680 82.030 290.350 83.120 ;
        RECT 290.980 82.030 291.270 83.195 ;
        RECT 292.375 83.080 293.130 83.250 ;
        RECT 292.415 82.030 292.700 82.900 ;
        RECT 292.870 82.830 293.130 83.080 ;
        RECT 293.920 83.170 294.090 83.420 ;
        RECT 294.260 83.340 294.610 83.910 ;
        RECT 294.780 83.170 294.950 84.080 ;
        RECT 293.920 83.000 294.950 83.170 ;
        RECT 292.870 82.660 293.990 82.830 ;
        RECT 292.870 82.200 293.130 82.660 ;
        RECT 293.305 82.030 293.560 82.490 ;
        RECT 293.730 82.200 293.990 82.660 ;
        RECT 294.160 82.030 294.470 82.830 ;
        RECT 294.640 82.200 294.950 83.000 ;
        RECT 295.585 83.840 295.840 84.410 ;
        RECT 296.010 84.180 296.340 84.580 ;
        RECT 296.765 84.045 297.295 84.410 ;
        RECT 296.765 84.010 296.940 84.045 ;
        RECT 296.010 83.840 296.940 84.010 ;
        RECT 297.485 83.900 297.760 84.410 ;
        RECT 295.585 83.170 295.755 83.840 ;
        RECT 296.010 83.670 296.180 83.840 ;
        RECT 295.925 83.340 296.180 83.670 ;
        RECT 296.405 83.340 296.600 83.670 ;
        RECT 295.585 82.200 295.920 83.170 ;
        RECT 296.090 82.030 296.260 83.170 ;
        RECT 296.430 82.370 296.600 83.340 ;
        RECT 296.770 82.710 296.940 83.840 ;
        RECT 297.110 83.050 297.280 83.850 ;
        RECT 297.480 83.730 297.760 83.900 ;
        RECT 297.485 83.250 297.760 83.730 ;
        RECT 297.930 83.050 298.120 84.410 ;
        RECT 298.300 84.045 298.810 84.580 ;
        RECT 299.030 83.770 299.275 84.375 ;
        RECT 299.725 84.030 299.980 84.320 ;
        RECT 300.150 84.200 300.480 84.580 ;
        RECT 299.725 83.860 300.475 84.030 ;
        RECT 298.320 83.600 299.550 83.770 ;
        RECT 297.110 82.880 298.120 83.050 ;
        RECT 298.290 83.035 299.040 83.225 ;
        RECT 296.770 82.540 297.895 82.710 ;
        RECT 298.290 82.370 298.460 83.035 ;
        RECT 299.210 82.790 299.550 83.600 ;
        RECT 299.725 83.040 300.075 83.690 ;
        RECT 300.245 82.870 300.475 83.860 ;
        RECT 296.430 82.200 298.460 82.370 ;
        RECT 298.630 82.030 298.800 82.790 ;
        RECT 299.035 82.380 299.550 82.790 ;
        RECT 299.725 82.700 300.475 82.870 ;
        RECT 299.725 82.200 299.980 82.700 ;
        RECT 300.150 82.030 300.480 82.530 ;
        RECT 300.650 82.200 300.820 84.320 ;
        RECT 301.180 84.220 301.510 84.580 ;
        RECT 301.680 84.190 302.175 84.360 ;
        RECT 302.380 84.190 303.235 84.360 ;
        RECT 301.050 83.000 301.510 84.050 ;
        RECT 300.990 82.215 301.315 83.000 ;
        RECT 301.680 82.830 301.850 84.190 ;
        RECT 302.020 83.280 302.370 83.900 ;
        RECT 302.540 83.680 302.895 83.900 ;
        RECT 302.540 83.090 302.710 83.680 ;
        RECT 303.065 83.480 303.235 84.190 ;
        RECT 304.110 84.120 304.440 84.580 ;
        RECT 304.650 84.220 305.000 84.390 ;
        RECT 303.440 83.650 304.230 83.900 ;
        RECT 304.650 83.830 304.910 84.220 ;
        RECT 305.220 84.130 306.170 84.410 ;
        RECT 306.340 84.140 306.530 84.580 ;
        RECT 306.700 84.200 307.770 84.370 ;
        RECT 304.400 83.480 304.570 83.660 ;
        RECT 301.680 82.660 302.075 82.830 ;
        RECT 302.245 82.700 302.710 83.090 ;
        RECT 302.880 83.310 304.570 83.480 ;
        RECT 301.905 82.530 302.075 82.660 ;
        RECT 302.880 82.530 303.050 83.310 ;
        RECT 304.740 83.140 304.910 83.830 ;
        RECT 303.410 82.970 304.910 83.140 ;
        RECT 305.100 83.170 305.310 83.960 ;
        RECT 305.480 83.340 305.830 83.960 ;
        RECT 306.000 83.350 306.170 84.130 ;
        RECT 306.700 83.970 306.870 84.200 ;
        RECT 306.340 83.800 306.870 83.970 ;
        RECT 306.340 83.520 306.560 83.800 ;
        RECT 307.040 83.630 307.280 84.030 ;
        RECT 306.000 83.180 306.405 83.350 ;
        RECT 306.740 83.260 307.280 83.630 ;
        RECT 307.450 83.845 307.770 84.200 ;
        RECT 308.015 84.120 308.320 84.580 ;
        RECT 308.490 83.870 308.740 84.400 ;
        RECT 307.450 83.670 307.775 83.845 ;
        RECT 307.450 83.370 308.365 83.670 ;
        RECT 307.625 83.340 308.365 83.370 ;
        RECT 305.100 83.010 305.775 83.170 ;
        RECT 306.235 83.090 306.405 83.180 ;
        RECT 305.100 83.000 306.065 83.010 ;
        RECT 304.740 82.830 304.910 82.970 ;
        RECT 301.485 82.030 301.735 82.490 ;
        RECT 301.905 82.200 302.155 82.530 ;
        RECT 302.370 82.200 303.050 82.530 ;
        RECT 303.220 82.630 304.295 82.800 ;
        RECT 304.740 82.660 305.300 82.830 ;
        RECT 305.605 82.710 306.065 83.000 ;
        RECT 306.235 82.920 307.455 83.090 ;
        RECT 303.220 82.290 303.390 82.630 ;
        RECT 303.625 82.030 303.955 82.460 ;
        RECT 304.125 82.290 304.295 82.630 ;
        RECT 304.590 82.030 304.960 82.490 ;
        RECT 305.130 82.200 305.300 82.660 ;
        RECT 306.235 82.540 306.405 82.920 ;
        RECT 307.625 82.750 307.795 83.340 ;
        RECT 308.535 83.220 308.740 83.870 ;
        RECT 308.910 83.825 309.160 84.580 ;
        RECT 309.840 83.830 311.050 84.580 ;
        RECT 305.535 82.200 306.405 82.540 ;
        RECT 306.995 82.580 307.795 82.750 ;
        RECT 306.575 82.030 306.825 82.490 ;
        RECT 306.995 82.290 307.165 82.580 ;
        RECT 307.345 82.030 307.675 82.410 ;
        RECT 308.015 82.030 308.320 83.170 ;
        RECT 308.490 82.340 308.740 83.220 ;
        RECT 308.910 82.030 309.160 83.170 ;
        RECT 309.840 83.120 310.360 83.660 ;
        RECT 310.530 83.290 311.050 83.830 ;
        RECT 309.840 82.030 311.050 83.120 ;
        RECT 162.095 81.860 311.135 82.030 ;
        RECT 162.180 80.770 163.390 81.860 ;
        RECT 163.560 81.425 168.905 81.860 ;
        RECT 162.180 80.060 162.700 80.600 ;
        RECT 162.870 80.230 163.390 80.770 ;
        RECT 162.180 79.310 163.390 80.060 ;
        RECT 165.145 79.855 165.485 80.685 ;
        RECT 166.965 80.175 167.315 81.425 ;
        RECT 169.540 80.785 169.810 81.690 ;
        RECT 169.980 81.100 170.310 81.860 ;
        RECT 170.490 80.930 170.660 81.690 ;
        RECT 169.540 79.985 169.710 80.785 ;
        RECT 169.995 80.760 170.660 80.930 ;
        RECT 170.920 80.785 171.190 81.690 ;
        RECT 171.360 81.100 171.690 81.860 ;
        RECT 171.870 80.930 172.040 81.690 ;
        RECT 169.995 80.615 170.165 80.760 ;
        RECT 169.880 80.285 170.165 80.615 ;
        RECT 169.995 80.030 170.165 80.285 ;
        RECT 170.400 80.210 170.730 80.580 ;
        RECT 163.560 79.310 168.905 79.855 ;
        RECT 169.540 79.480 169.800 79.985 ;
        RECT 169.995 79.860 170.660 80.030 ;
        RECT 169.980 79.310 170.310 79.690 ;
        RECT 170.490 79.480 170.660 79.860 ;
        RECT 170.920 79.985 171.090 80.785 ;
        RECT 171.375 80.760 172.040 80.930 ;
        RECT 173.310 80.930 173.480 81.690 ;
        RECT 173.660 81.100 173.990 81.860 ;
        RECT 173.310 80.760 173.975 80.930 ;
        RECT 174.160 80.785 174.430 81.690 ;
        RECT 171.375 80.615 171.545 80.760 ;
        RECT 171.260 80.285 171.545 80.615 ;
        RECT 173.805 80.615 173.975 80.760 ;
        RECT 171.375 80.030 171.545 80.285 ;
        RECT 171.780 80.210 172.110 80.580 ;
        RECT 173.240 80.210 173.570 80.580 ;
        RECT 173.805 80.285 174.090 80.615 ;
        RECT 173.805 80.030 173.975 80.285 ;
        RECT 170.920 79.480 171.180 79.985 ;
        RECT 171.375 79.860 172.040 80.030 ;
        RECT 171.360 79.310 171.690 79.690 ;
        RECT 171.870 79.480 172.040 79.860 ;
        RECT 173.310 79.860 173.975 80.030 ;
        RECT 174.260 79.985 174.430 80.785 ;
        RECT 175.060 80.695 175.350 81.860 ;
        RECT 175.525 80.720 175.860 81.690 ;
        RECT 176.030 80.720 176.200 81.860 ;
        RECT 176.370 81.520 178.400 81.690 ;
        RECT 175.525 80.050 175.695 80.720 ;
        RECT 176.370 80.550 176.540 81.520 ;
        RECT 175.865 80.220 176.120 80.550 ;
        RECT 176.345 80.220 176.540 80.550 ;
        RECT 176.710 81.180 177.835 81.350 ;
        RECT 175.950 80.050 176.120 80.220 ;
        RECT 176.710 80.050 176.880 81.180 ;
        RECT 173.310 79.480 173.480 79.860 ;
        RECT 173.660 79.310 173.990 79.690 ;
        RECT 174.170 79.480 174.430 79.985 ;
        RECT 175.060 79.310 175.350 80.035 ;
        RECT 175.525 79.480 175.780 80.050 ;
        RECT 175.950 79.880 176.880 80.050 ;
        RECT 177.050 80.840 178.060 81.010 ;
        RECT 177.050 80.040 177.220 80.840 ;
        RECT 177.425 80.500 177.700 80.640 ;
        RECT 177.420 80.330 177.700 80.500 ;
        RECT 176.705 79.845 176.880 79.880 ;
        RECT 175.950 79.310 176.280 79.710 ;
        RECT 176.705 79.480 177.235 79.845 ;
        RECT 177.425 79.480 177.700 80.330 ;
        RECT 177.870 79.480 178.060 80.840 ;
        RECT 178.230 80.855 178.400 81.520 ;
        RECT 178.570 81.100 178.740 81.860 ;
        RECT 178.975 81.100 179.490 81.510 ;
        RECT 179.660 81.425 185.005 81.860 ;
        RECT 178.230 80.665 178.980 80.855 ;
        RECT 179.150 80.290 179.490 81.100 ;
        RECT 178.260 80.120 179.490 80.290 ;
        RECT 178.240 79.310 178.750 79.845 ;
        RECT 178.970 79.515 179.215 80.120 ;
        RECT 181.245 79.855 181.585 80.685 ;
        RECT 183.065 80.175 183.415 81.425 ;
        RECT 185.730 80.930 185.900 81.690 ;
        RECT 186.080 81.100 186.410 81.860 ;
        RECT 185.730 80.760 186.395 80.930 ;
        RECT 186.580 80.785 186.850 81.690 ;
        RECT 187.025 81.190 187.280 81.690 ;
        RECT 187.450 81.360 187.780 81.860 ;
        RECT 187.025 81.020 187.775 81.190 ;
        RECT 186.225 80.615 186.395 80.760 ;
        RECT 185.660 80.210 185.990 80.580 ;
        RECT 186.225 80.285 186.510 80.615 ;
        RECT 186.225 80.030 186.395 80.285 ;
        RECT 185.730 79.860 186.395 80.030 ;
        RECT 186.680 79.985 186.850 80.785 ;
        RECT 187.025 80.200 187.375 80.850 ;
        RECT 187.545 80.030 187.775 81.020 ;
        RECT 179.660 79.310 185.005 79.855 ;
        RECT 185.730 79.480 185.900 79.860 ;
        RECT 186.080 79.310 186.410 79.690 ;
        RECT 186.590 79.480 186.850 79.985 ;
        RECT 187.025 79.860 187.775 80.030 ;
        RECT 187.025 79.570 187.280 79.860 ;
        RECT 187.450 79.310 187.780 79.690 ;
        RECT 187.950 79.570 188.120 81.690 ;
        RECT 188.290 80.890 188.615 81.675 ;
        RECT 188.785 81.400 189.035 81.860 ;
        RECT 189.205 81.360 189.455 81.690 ;
        RECT 189.670 81.360 190.350 81.690 ;
        RECT 189.205 81.230 189.375 81.360 ;
        RECT 188.980 81.060 189.375 81.230 ;
        RECT 188.350 79.840 188.810 80.890 ;
        RECT 188.980 79.700 189.150 81.060 ;
        RECT 189.545 80.800 190.010 81.190 ;
        RECT 189.320 79.990 189.670 80.610 ;
        RECT 189.840 80.210 190.010 80.800 ;
        RECT 190.180 80.580 190.350 81.360 ;
        RECT 190.520 81.260 190.690 81.600 ;
        RECT 190.925 81.430 191.255 81.860 ;
        RECT 191.425 81.260 191.595 81.600 ;
        RECT 191.890 81.400 192.260 81.860 ;
        RECT 190.520 81.090 191.595 81.260 ;
        RECT 192.430 81.230 192.600 81.690 ;
        RECT 192.835 81.350 193.705 81.690 ;
        RECT 193.875 81.400 194.125 81.860 ;
        RECT 192.040 81.060 192.600 81.230 ;
        RECT 192.040 80.920 192.210 81.060 ;
        RECT 190.710 80.750 192.210 80.920 ;
        RECT 192.905 80.890 193.365 81.180 ;
        RECT 190.180 80.410 191.870 80.580 ;
        RECT 189.840 79.990 190.195 80.210 ;
        RECT 190.365 79.700 190.535 80.410 ;
        RECT 190.740 79.990 191.530 80.240 ;
        RECT 191.700 80.230 191.870 80.410 ;
        RECT 192.040 80.060 192.210 80.750 ;
        RECT 188.480 79.310 188.810 79.670 ;
        RECT 188.980 79.530 189.475 79.700 ;
        RECT 189.680 79.530 190.535 79.700 ;
        RECT 191.410 79.310 191.740 79.770 ;
        RECT 191.950 79.670 192.210 80.060 ;
        RECT 192.400 80.880 193.365 80.890 ;
        RECT 193.535 80.970 193.705 81.350 ;
        RECT 194.295 81.310 194.465 81.600 ;
        RECT 194.645 81.480 194.975 81.860 ;
        RECT 194.295 81.140 195.095 81.310 ;
        RECT 192.400 80.720 193.075 80.880 ;
        RECT 193.535 80.800 194.755 80.970 ;
        RECT 192.400 79.930 192.610 80.720 ;
        RECT 193.535 80.710 193.705 80.800 ;
        RECT 192.780 79.930 193.130 80.550 ;
        RECT 193.300 80.540 193.705 80.710 ;
        RECT 193.300 79.760 193.470 80.540 ;
        RECT 193.640 80.090 193.860 80.370 ;
        RECT 194.040 80.260 194.580 80.630 ;
        RECT 194.925 80.550 195.095 81.140 ;
        RECT 195.315 80.720 195.620 81.860 ;
        RECT 195.790 80.670 196.045 81.550 ;
        RECT 196.220 80.770 199.730 81.860 ;
        RECT 194.925 80.520 195.665 80.550 ;
        RECT 193.640 79.920 194.170 80.090 ;
        RECT 191.950 79.500 192.300 79.670 ;
        RECT 192.520 79.480 193.470 79.760 ;
        RECT 193.640 79.310 193.830 79.750 ;
        RECT 194.000 79.690 194.170 79.920 ;
        RECT 194.340 79.860 194.580 80.260 ;
        RECT 194.750 80.220 195.665 80.520 ;
        RECT 194.750 80.045 195.075 80.220 ;
        RECT 194.750 79.690 195.070 80.045 ;
        RECT 195.835 80.020 196.045 80.670 ;
        RECT 194.000 79.520 195.070 79.690 ;
        RECT 195.315 79.310 195.620 79.770 ;
        RECT 195.790 79.490 196.045 80.020 ;
        RECT 196.220 80.080 197.870 80.600 ;
        RECT 198.040 80.250 199.730 80.770 ;
        RECT 200.820 80.695 201.110 81.860 ;
        RECT 201.280 81.425 206.625 81.860 ;
        RECT 196.220 79.310 199.730 80.080 ;
        RECT 200.820 79.310 201.110 80.035 ;
        RECT 202.865 79.855 203.205 80.685 ;
        RECT 204.685 80.175 205.035 81.425 ;
        RECT 207.720 80.720 208.010 81.860 ;
        RECT 208.180 81.140 208.630 81.690 ;
        RECT 208.820 81.140 209.150 81.860 ;
        RECT 201.280 79.310 206.625 79.855 ;
        RECT 207.720 79.310 208.010 80.110 ;
        RECT 208.180 79.770 208.430 81.140 ;
        RECT 209.360 80.970 209.660 81.520 ;
        RECT 209.830 81.190 210.110 81.860 ;
        RECT 210.480 81.425 215.825 81.860 ;
        RECT 208.720 80.800 209.660 80.970 ;
        RECT 208.720 80.550 208.890 80.800 ;
        RECT 209.995 80.550 210.310 80.990 ;
        RECT 208.600 80.220 208.890 80.550 ;
        RECT 209.060 80.300 209.390 80.550 ;
        RECT 209.620 80.300 210.310 80.550 ;
        RECT 208.720 80.130 208.890 80.220 ;
        RECT 208.720 79.940 210.110 80.130 ;
        RECT 208.180 79.480 208.730 79.770 ;
        RECT 208.900 79.310 209.150 79.770 ;
        RECT 209.780 79.580 210.110 79.940 ;
        RECT 212.065 79.855 212.405 80.685 ;
        RECT 213.885 80.175 214.235 81.425 ;
        RECT 216.000 80.770 218.590 81.860 ;
        RECT 219.900 81.500 220.230 81.860 ;
        RECT 220.755 81.500 221.090 81.860 ;
        RECT 221.660 81.500 221.990 81.860 ;
        RECT 222.555 81.500 223.005 81.860 ;
        RECT 216.000 80.080 217.210 80.600 ;
        RECT 217.380 80.250 218.590 80.770 ;
        RECT 219.290 81.100 223.055 81.330 ;
        RECT 210.480 79.310 215.825 79.855 ;
        RECT 216.000 79.310 218.590 80.080 ;
        RECT 219.290 79.650 219.570 81.100 ;
        RECT 219.740 79.840 220.020 80.930 ;
        RECT 220.200 80.760 221.510 80.930 ;
        RECT 220.200 80.070 220.465 80.760 ;
        RECT 221.680 80.750 222.455 80.920 ;
        RECT 221.680 80.580 221.850 80.750 ;
        RECT 220.635 80.245 221.850 80.580 ;
        RECT 220.200 79.840 221.450 80.070 ;
        RECT 221.620 80.030 221.850 80.245 ;
        RECT 222.020 80.220 222.210 80.565 ;
        RECT 221.620 79.840 222.315 80.030 ;
        RECT 222.500 79.950 222.715 80.565 ;
        RECT 222.885 80.550 223.055 81.100 ;
        RECT 223.225 80.720 223.585 81.390 ;
        RECT 223.820 80.770 226.410 81.860 ;
        RECT 222.885 80.220 223.195 80.550 ;
        RECT 223.365 80.030 223.585 80.720 ;
        RECT 219.900 79.310 220.230 79.670 ;
        RECT 220.400 79.480 220.590 79.840 ;
        RECT 221.260 79.740 221.450 79.840 ;
        RECT 222.135 79.770 222.315 79.840 ;
        RECT 223.100 79.770 223.585 80.030 ;
        RECT 220.760 79.310 221.090 79.670 ;
        RECT 221.625 79.310 221.955 79.670 ;
        RECT 222.135 79.580 223.585 79.770 ;
        RECT 223.100 79.480 223.585 79.580 ;
        RECT 223.820 80.080 225.030 80.600 ;
        RECT 225.200 80.250 226.410 80.770 ;
        RECT 226.580 80.695 226.870 81.860 ;
        RECT 227.040 81.010 227.300 81.690 ;
        RECT 227.470 81.080 227.720 81.860 ;
        RECT 227.970 81.310 228.220 81.690 ;
        RECT 228.390 81.480 228.745 81.860 ;
        RECT 229.750 81.470 230.085 81.690 ;
        RECT 229.350 81.310 229.580 81.350 ;
        RECT 227.970 81.110 229.580 81.310 ;
        RECT 227.970 81.100 228.805 81.110 ;
        RECT 229.395 81.020 229.580 81.110 ;
        RECT 223.820 79.310 226.410 80.080 ;
        RECT 226.580 79.310 226.870 80.035 ;
        RECT 227.040 79.820 227.210 81.010 ;
        RECT 228.910 80.910 229.240 80.940 ;
        RECT 227.440 80.850 229.240 80.910 ;
        RECT 229.830 80.850 230.085 81.470 ;
        RECT 230.260 81.425 235.605 81.860 ;
        RECT 236.705 81.470 237.040 81.690 ;
        RECT 238.045 81.480 238.400 81.860 ;
        RECT 227.380 80.740 230.085 80.850 ;
        RECT 227.380 80.705 227.580 80.740 ;
        RECT 227.380 80.130 227.550 80.705 ;
        RECT 228.910 80.680 230.085 80.740 ;
        RECT 227.780 80.265 228.190 80.570 ;
        RECT 228.360 80.300 228.690 80.510 ;
        RECT 227.380 80.010 227.650 80.130 ;
        RECT 227.380 79.965 228.225 80.010 ;
        RECT 227.470 79.840 228.225 79.965 ;
        RECT 228.480 79.900 228.690 80.300 ;
        RECT 228.935 80.300 229.410 80.510 ;
        RECT 229.600 80.300 230.090 80.500 ;
        RECT 228.935 79.900 229.155 80.300 ;
        RECT 227.040 79.810 227.270 79.820 ;
        RECT 227.040 79.480 227.300 79.810 ;
        RECT 228.055 79.690 228.225 79.840 ;
        RECT 227.470 79.310 227.800 79.670 ;
        RECT 228.055 79.480 229.355 79.690 ;
        RECT 229.630 79.310 230.085 80.075 ;
        RECT 231.845 79.855 232.185 80.685 ;
        RECT 233.665 80.175 234.015 81.425 ;
        RECT 236.705 80.850 236.960 81.470 ;
        RECT 237.210 81.310 237.440 81.350 ;
        RECT 238.570 81.310 238.820 81.690 ;
        RECT 237.210 81.110 238.820 81.310 ;
        RECT 237.210 81.020 237.395 81.110 ;
        RECT 237.985 81.100 238.820 81.110 ;
        RECT 239.070 81.080 239.320 81.860 ;
        RECT 239.490 81.010 239.750 81.690 ;
        RECT 237.550 80.910 237.880 80.940 ;
        RECT 237.550 80.850 239.350 80.910 ;
        RECT 236.705 80.740 239.410 80.850 ;
        RECT 236.705 80.680 237.880 80.740 ;
        RECT 239.210 80.705 239.410 80.740 ;
        RECT 236.700 80.300 237.190 80.500 ;
        RECT 237.380 80.300 237.855 80.510 ;
        RECT 230.260 79.310 235.605 79.855 ;
        RECT 236.705 79.310 237.160 80.075 ;
        RECT 237.635 79.900 237.855 80.300 ;
        RECT 238.100 80.300 238.430 80.510 ;
        RECT 238.100 79.900 238.310 80.300 ;
        RECT 238.600 80.265 239.010 80.570 ;
        RECT 239.240 80.130 239.410 80.705 ;
        RECT 239.140 80.010 239.410 80.130 ;
        RECT 238.565 79.965 239.410 80.010 ;
        RECT 238.565 79.840 239.320 79.965 ;
        RECT 238.565 79.690 238.735 79.840 ;
        RECT 239.580 79.820 239.750 81.010 ;
        RECT 240.010 80.850 240.180 81.690 ;
        RECT 240.350 81.520 241.520 81.690 ;
        RECT 240.350 81.020 240.680 81.520 ;
        RECT 241.190 81.480 241.520 81.520 ;
        RECT 241.710 81.440 242.065 81.860 ;
        RECT 240.850 81.260 241.080 81.350 ;
        RECT 242.235 81.260 242.485 81.690 ;
        RECT 240.850 81.020 242.485 81.260 ;
        RECT 242.655 81.100 242.985 81.860 ;
        RECT 243.155 81.020 243.410 81.690 ;
        RECT 240.010 80.680 243.070 80.850 ;
        RECT 239.925 80.300 240.275 80.510 ;
        RECT 240.445 80.300 240.890 80.500 ;
        RECT 241.060 80.300 241.535 80.500 ;
        RECT 239.520 79.810 239.750 79.820 ;
        RECT 237.435 79.480 238.735 79.690 ;
        RECT 238.990 79.310 239.320 79.670 ;
        RECT 239.490 79.480 239.750 79.810 ;
        RECT 240.010 79.960 241.075 80.130 ;
        RECT 240.010 79.480 240.180 79.960 ;
        RECT 240.350 79.310 240.680 79.790 ;
        RECT 240.905 79.730 241.075 79.960 ;
        RECT 241.255 79.900 241.535 80.300 ;
        RECT 241.805 80.300 242.135 80.500 ;
        RECT 242.305 80.330 242.680 80.500 ;
        RECT 242.305 80.300 242.670 80.330 ;
        RECT 241.805 79.900 242.090 80.300 ;
        RECT 242.900 80.130 243.070 80.680 ;
        RECT 242.270 79.960 243.070 80.130 ;
        RECT 242.270 79.730 242.440 79.960 ;
        RECT 243.240 79.890 243.410 81.020 ;
        RECT 243.690 80.850 243.860 81.690 ;
        RECT 244.030 81.520 245.200 81.690 ;
        RECT 244.030 81.020 244.360 81.520 ;
        RECT 244.870 81.480 245.200 81.520 ;
        RECT 245.390 81.440 245.745 81.860 ;
        RECT 244.530 81.260 244.760 81.350 ;
        RECT 245.915 81.260 246.165 81.690 ;
        RECT 244.530 81.020 246.165 81.260 ;
        RECT 246.335 81.100 246.665 81.860 ;
        RECT 246.835 81.020 247.090 81.690 ;
        RECT 243.690 80.680 246.750 80.850 ;
        RECT 243.605 80.300 243.955 80.510 ;
        RECT 244.125 80.300 244.570 80.500 ;
        RECT 244.740 80.300 245.215 80.500 ;
        RECT 243.225 79.820 243.410 79.890 ;
        RECT 243.200 79.810 243.410 79.820 ;
        RECT 240.905 79.480 242.440 79.730 ;
        RECT 242.610 79.310 242.940 79.790 ;
        RECT 243.155 79.480 243.410 79.810 ;
        RECT 243.690 79.960 244.755 80.130 ;
        RECT 243.690 79.480 243.860 79.960 ;
        RECT 244.030 79.310 244.360 79.790 ;
        RECT 244.585 79.730 244.755 79.960 ;
        RECT 244.935 79.900 245.215 80.300 ;
        RECT 245.485 80.300 245.815 80.500 ;
        RECT 245.985 80.330 246.360 80.500 ;
        RECT 245.985 80.300 246.350 80.330 ;
        RECT 245.485 79.900 245.770 80.300 ;
        RECT 246.580 80.130 246.750 80.680 ;
        RECT 245.950 79.960 246.750 80.130 ;
        RECT 245.950 79.730 246.120 79.960 ;
        RECT 246.920 79.890 247.090 81.020 ;
        RECT 247.280 80.770 250.790 81.860 ;
        RECT 250.960 80.770 252.170 81.860 ;
        RECT 246.905 79.820 247.090 79.890 ;
        RECT 246.880 79.810 247.090 79.820 ;
        RECT 244.585 79.480 246.120 79.730 ;
        RECT 246.290 79.310 246.620 79.790 ;
        RECT 246.835 79.480 247.090 79.810 ;
        RECT 247.280 80.080 248.930 80.600 ;
        RECT 249.100 80.250 250.790 80.770 ;
        RECT 247.280 79.310 250.790 80.080 ;
        RECT 250.960 80.060 251.480 80.600 ;
        RECT 251.650 80.230 252.170 80.770 ;
        RECT 252.340 80.695 252.630 81.860 ;
        RECT 252.800 81.425 258.145 81.860 ;
        RECT 250.960 79.310 252.170 80.060 ;
        RECT 252.340 79.310 252.630 80.035 ;
        RECT 254.385 79.855 254.725 80.685 ;
        RECT 256.205 80.175 256.555 81.425 ;
        RECT 258.320 81.010 258.580 81.690 ;
        RECT 258.750 81.080 259.000 81.860 ;
        RECT 259.250 81.310 259.500 81.690 ;
        RECT 259.670 81.480 260.025 81.860 ;
        RECT 261.030 81.470 261.365 81.690 ;
        RECT 260.630 81.310 260.860 81.350 ;
        RECT 259.250 81.110 260.860 81.310 ;
        RECT 259.250 81.100 260.085 81.110 ;
        RECT 260.675 81.020 260.860 81.110 ;
        RECT 252.800 79.310 258.145 79.855 ;
        RECT 258.320 79.820 258.490 81.010 ;
        RECT 260.190 80.910 260.520 80.940 ;
        RECT 258.720 80.850 260.520 80.910 ;
        RECT 261.110 80.850 261.365 81.470 ;
        RECT 261.540 81.425 266.885 81.860 ;
        RECT 267.060 81.425 272.405 81.860 ;
        RECT 258.660 80.740 261.365 80.850 ;
        RECT 258.660 80.705 258.860 80.740 ;
        RECT 258.660 80.130 258.830 80.705 ;
        RECT 260.190 80.680 261.365 80.740 ;
        RECT 259.060 80.265 259.470 80.570 ;
        RECT 259.640 80.300 259.970 80.510 ;
        RECT 258.660 80.010 258.930 80.130 ;
        RECT 258.660 79.965 259.505 80.010 ;
        RECT 258.750 79.840 259.505 79.965 ;
        RECT 259.760 79.900 259.970 80.300 ;
        RECT 260.215 80.300 260.690 80.510 ;
        RECT 260.880 80.300 261.370 80.500 ;
        RECT 260.215 79.900 260.435 80.300 ;
        RECT 258.320 79.810 258.550 79.820 ;
        RECT 258.320 79.480 258.580 79.810 ;
        RECT 259.335 79.690 259.505 79.840 ;
        RECT 258.750 79.310 259.080 79.670 ;
        RECT 259.335 79.480 260.635 79.690 ;
        RECT 260.910 79.310 261.365 80.075 ;
        RECT 263.125 79.855 263.465 80.685 ;
        RECT 264.945 80.175 265.295 81.425 ;
        RECT 268.645 79.855 268.985 80.685 ;
        RECT 270.465 80.175 270.815 81.425 ;
        RECT 272.580 80.770 273.790 81.860 ;
        RECT 272.580 80.060 273.100 80.600 ;
        RECT 273.270 80.230 273.790 80.770 ;
        RECT 273.960 80.785 274.230 81.690 ;
        RECT 274.400 81.100 274.730 81.860 ;
        RECT 274.910 80.930 275.080 81.690 ;
        RECT 261.540 79.310 266.885 79.855 ;
        RECT 267.060 79.310 272.405 79.855 ;
        RECT 272.580 79.310 273.790 80.060 ;
        RECT 273.960 79.985 274.130 80.785 ;
        RECT 274.415 80.760 275.080 80.930 ;
        RECT 275.340 80.785 275.610 81.690 ;
        RECT 275.780 81.100 276.110 81.860 ;
        RECT 276.290 80.930 276.460 81.690 ;
        RECT 274.415 80.615 274.585 80.760 ;
        RECT 274.300 80.285 274.585 80.615 ;
        RECT 274.415 80.030 274.585 80.285 ;
        RECT 274.820 80.210 275.150 80.580 ;
        RECT 273.960 79.480 274.220 79.985 ;
        RECT 274.415 79.860 275.080 80.030 ;
        RECT 274.400 79.310 274.730 79.690 ;
        RECT 274.910 79.480 275.080 79.860 ;
        RECT 275.340 79.985 275.510 80.785 ;
        RECT 275.795 80.760 276.460 80.930 ;
        RECT 276.720 80.770 277.930 81.860 ;
        RECT 275.795 80.615 275.965 80.760 ;
        RECT 275.680 80.285 275.965 80.615 ;
        RECT 275.795 80.030 275.965 80.285 ;
        RECT 276.200 80.210 276.530 80.580 ;
        RECT 276.720 80.060 277.240 80.600 ;
        RECT 277.410 80.230 277.930 80.770 ;
        RECT 278.100 80.695 278.390 81.860 ;
        RECT 278.560 81.425 283.905 81.860 ;
        RECT 275.340 79.480 275.600 79.985 ;
        RECT 275.795 79.860 276.460 80.030 ;
        RECT 275.780 79.310 276.110 79.690 ;
        RECT 276.290 79.480 276.460 79.860 ;
        RECT 276.720 79.310 277.930 80.060 ;
        RECT 278.100 79.310 278.390 80.035 ;
        RECT 280.145 79.855 280.485 80.685 ;
        RECT 281.965 80.175 282.315 81.425 ;
        RECT 285.005 81.190 285.260 81.690 ;
        RECT 285.430 81.360 285.760 81.860 ;
        RECT 285.005 81.020 285.755 81.190 ;
        RECT 285.005 80.200 285.355 80.850 ;
        RECT 285.525 80.030 285.755 81.020 ;
        RECT 285.005 79.860 285.755 80.030 ;
        RECT 278.560 79.310 283.905 79.855 ;
        RECT 285.005 79.570 285.260 79.860 ;
        RECT 285.430 79.310 285.760 79.690 ;
        RECT 285.930 79.570 286.100 81.690 ;
        RECT 286.270 80.890 286.595 81.675 ;
        RECT 286.765 81.400 287.015 81.860 ;
        RECT 287.185 81.360 287.435 81.690 ;
        RECT 287.650 81.360 288.330 81.690 ;
        RECT 287.185 81.230 287.355 81.360 ;
        RECT 286.960 81.060 287.355 81.230 ;
        RECT 286.330 79.840 286.790 80.890 ;
        RECT 286.960 79.700 287.130 81.060 ;
        RECT 287.525 80.800 287.990 81.190 ;
        RECT 287.300 79.990 287.650 80.610 ;
        RECT 287.820 80.210 287.990 80.800 ;
        RECT 288.160 80.580 288.330 81.360 ;
        RECT 288.500 81.260 288.670 81.600 ;
        RECT 288.905 81.430 289.235 81.860 ;
        RECT 289.405 81.260 289.575 81.600 ;
        RECT 289.870 81.400 290.240 81.860 ;
        RECT 288.500 81.090 289.575 81.260 ;
        RECT 290.410 81.230 290.580 81.690 ;
        RECT 290.815 81.350 291.685 81.690 ;
        RECT 291.855 81.400 292.105 81.860 ;
        RECT 290.020 81.060 290.580 81.230 ;
        RECT 290.020 80.920 290.190 81.060 ;
        RECT 288.690 80.750 290.190 80.920 ;
        RECT 290.885 80.890 291.345 81.180 ;
        RECT 288.160 80.410 289.850 80.580 ;
        RECT 287.820 79.990 288.175 80.210 ;
        RECT 288.345 79.700 288.515 80.410 ;
        RECT 288.720 79.990 289.510 80.240 ;
        RECT 289.680 80.230 289.850 80.410 ;
        RECT 290.020 80.060 290.190 80.750 ;
        RECT 286.460 79.310 286.790 79.670 ;
        RECT 286.960 79.530 287.455 79.700 ;
        RECT 287.660 79.530 288.515 79.700 ;
        RECT 289.390 79.310 289.720 79.770 ;
        RECT 289.930 79.670 290.190 80.060 ;
        RECT 290.380 80.880 291.345 80.890 ;
        RECT 291.515 80.970 291.685 81.350 ;
        RECT 292.275 81.310 292.445 81.600 ;
        RECT 292.625 81.480 292.955 81.860 ;
        RECT 292.275 81.140 293.075 81.310 ;
        RECT 290.380 80.720 291.055 80.880 ;
        RECT 291.515 80.800 292.735 80.970 ;
        RECT 290.380 79.930 290.590 80.720 ;
        RECT 291.515 80.710 291.685 80.800 ;
        RECT 290.760 79.930 291.110 80.550 ;
        RECT 291.280 80.540 291.685 80.710 ;
        RECT 291.280 79.760 291.450 80.540 ;
        RECT 291.620 80.090 291.840 80.370 ;
        RECT 292.020 80.260 292.560 80.630 ;
        RECT 292.905 80.550 293.075 81.140 ;
        RECT 293.295 80.720 293.600 81.860 ;
        RECT 293.770 80.670 294.020 81.550 ;
        RECT 294.190 80.720 294.440 81.860 ;
        RECT 294.665 80.720 295.000 81.690 ;
        RECT 295.170 80.720 295.340 81.860 ;
        RECT 295.510 81.520 297.540 81.690 ;
        RECT 292.905 80.520 293.645 80.550 ;
        RECT 291.620 79.920 292.150 80.090 ;
        RECT 289.930 79.500 290.280 79.670 ;
        RECT 290.500 79.480 291.450 79.760 ;
        RECT 291.620 79.310 291.810 79.750 ;
        RECT 291.980 79.690 292.150 79.920 ;
        RECT 292.320 79.860 292.560 80.260 ;
        RECT 292.730 80.220 293.645 80.520 ;
        RECT 292.730 80.045 293.055 80.220 ;
        RECT 292.730 79.690 293.050 80.045 ;
        RECT 293.815 80.020 294.020 80.670 ;
        RECT 291.980 79.520 293.050 79.690 ;
        RECT 293.295 79.310 293.600 79.770 ;
        RECT 293.770 79.490 294.020 80.020 ;
        RECT 294.190 79.310 294.440 80.065 ;
        RECT 294.665 80.050 294.835 80.720 ;
        RECT 295.510 80.550 295.680 81.520 ;
        RECT 295.005 80.220 295.260 80.550 ;
        RECT 295.485 80.220 295.680 80.550 ;
        RECT 295.850 81.180 296.975 81.350 ;
        RECT 295.090 80.050 295.260 80.220 ;
        RECT 295.850 80.050 296.020 81.180 ;
        RECT 294.665 79.480 294.920 80.050 ;
        RECT 295.090 79.880 296.020 80.050 ;
        RECT 296.190 80.840 297.200 81.010 ;
        RECT 296.190 80.040 296.360 80.840 ;
        RECT 295.845 79.845 296.020 79.880 ;
        RECT 295.090 79.310 295.420 79.710 ;
        RECT 295.845 79.480 296.375 79.845 ;
        RECT 296.565 79.820 296.840 80.640 ;
        RECT 296.560 79.650 296.840 79.820 ;
        RECT 296.565 79.480 296.840 79.650 ;
        RECT 297.010 79.480 297.200 80.840 ;
        RECT 297.370 80.855 297.540 81.520 ;
        RECT 297.710 81.100 297.880 81.860 ;
        RECT 298.115 81.100 298.630 81.510 ;
        RECT 297.370 80.665 298.120 80.855 ;
        RECT 298.290 80.290 298.630 81.100 ;
        RECT 297.400 80.120 298.630 80.290 ;
        RECT 298.805 80.720 299.140 81.690 ;
        RECT 299.310 80.720 299.480 81.860 ;
        RECT 299.650 81.520 301.680 81.690 ;
        RECT 297.380 79.310 297.890 79.845 ;
        RECT 298.110 79.515 298.355 80.120 ;
        RECT 298.805 80.050 298.975 80.720 ;
        RECT 299.650 80.550 299.820 81.520 ;
        RECT 299.145 80.220 299.400 80.550 ;
        RECT 299.625 80.220 299.820 80.550 ;
        RECT 299.990 81.180 301.115 81.350 ;
        RECT 299.230 80.050 299.400 80.220 ;
        RECT 299.990 80.050 300.160 81.180 ;
        RECT 298.805 79.480 299.060 80.050 ;
        RECT 299.230 79.880 300.160 80.050 ;
        RECT 300.330 80.840 301.340 81.010 ;
        RECT 300.330 80.040 300.500 80.840 ;
        RECT 300.705 80.500 300.980 80.640 ;
        RECT 300.700 80.330 300.980 80.500 ;
        RECT 299.985 79.845 300.160 79.880 ;
        RECT 299.230 79.310 299.560 79.710 ;
        RECT 299.985 79.480 300.515 79.845 ;
        RECT 300.705 79.480 300.980 80.330 ;
        RECT 301.150 79.480 301.340 80.840 ;
        RECT 301.510 80.855 301.680 81.520 ;
        RECT 301.850 81.100 302.020 81.860 ;
        RECT 302.255 81.100 302.770 81.510 ;
        RECT 301.510 80.665 302.260 80.855 ;
        RECT 302.430 80.290 302.770 81.100 ;
        RECT 303.860 80.695 304.150 81.860 ;
        RECT 304.320 80.785 304.590 81.690 ;
        RECT 304.760 81.100 305.090 81.860 ;
        RECT 305.270 80.930 305.440 81.690 ;
        RECT 301.540 80.120 302.770 80.290 ;
        RECT 301.520 79.310 302.030 79.845 ;
        RECT 302.250 79.515 302.495 80.120 ;
        RECT 303.860 79.310 304.150 80.035 ;
        RECT 304.320 79.985 304.490 80.785 ;
        RECT 304.775 80.760 305.440 80.930 ;
        RECT 305.700 80.770 309.210 81.860 ;
        RECT 304.775 80.615 304.945 80.760 ;
        RECT 304.660 80.285 304.945 80.615 ;
        RECT 304.775 80.030 304.945 80.285 ;
        RECT 305.180 80.210 305.510 80.580 ;
        RECT 305.700 80.080 307.350 80.600 ;
        RECT 307.520 80.250 309.210 80.770 ;
        RECT 309.840 80.770 311.050 81.860 ;
        RECT 309.840 80.230 310.360 80.770 ;
        RECT 304.320 79.480 304.580 79.985 ;
        RECT 304.775 79.860 305.440 80.030 ;
        RECT 304.760 79.310 305.090 79.690 ;
        RECT 305.270 79.480 305.440 79.860 ;
        RECT 305.700 79.310 309.210 80.080 ;
        RECT 310.530 80.060 311.050 80.600 ;
        RECT 309.840 79.310 311.050 80.060 ;
        RECT 162.095 79.140 311.135 79.310 ;
        RECT 162.180 78.390 163.390 79.140 ;
        RECT 162.180 77.850 162.700 78.390 ;
        RECT 163.560 78.370 167.070 79.140 ;
        RECT 168.165 78.590 168.420 78.880 ;
        RECT 168.590 78.760 168.920 79.140 ;
        RECT 168.165 78.420 168.915 78.590 ;
        RECT 162.870 77.680 163.390 78.220 ;
        RECT 163.560 77.850 165.210 78.370 ;
        RECT 165.380 77.680 167.070 78.200 ;
        RECT 162.180 76.590 163.390 77.680 ;
        RECT 163.560 76.590 167.070 77.680 ;
        RECT 168.165 77.600 168.515 78.250 ;
        RECT 168.685 77.430 168.915 78.420 ;
        RECT 168.165 77.260 168.915 77.430 ;
        RECT 168.165 76.760 168.420 77.260 ;
        RECT 168.590 76.590 168.920 77.090 ;
        RECT 169.090 76.760 169.260 78.880 ;
        RECT 169.620 78.780 169.950 79.140 ;
        RECT 170.120 78.750 170.615 78.920 ;
        RECT 170.820 78.750 171.675 78.920 ;
        RECT 169.490 77.560 169.950 78.610 ;
        RECT 169.430 76.775 169.755 77.560 ;
        RECT 170.120 77.390 170.290 78.750 ;
        RECT 170.460 77.840 170.810 78.460 ;
        RECT 170.980 78.240 171.335 78.460 ;
        RECT 170.980 77.650 171.150 78.240 ;
        RECT 171.505 78.040 171.675 78.750 ;
        RECT 172.550 78.680 172.880 79.140 ;
        RECT 173.090 78.780 173.440 78.950 ;
        RECT 171.880 78.210 172.670 78.460 ;
        RECT 173.090 78.390 173.350 78.780 ;
        RECT 173.660 78.690 174.610 78.970 ;
        RECT 174.780 78.700 174.970 79.140 ;
        RECT 175.140 78.760 176.210 78.930 ;
        RECT 172.840 78.040 173.010 78.220 ;
        RECT 170.120 77.220 170.515 77.390 ;
        RECT 170.685 77.260 171.150 77.650 ;
        RECT 171.320 77.870 173.010 78.040 ;
        RECT 170.345 77.090 170.515 77.220 ;
        RECT 171.320 77.090 171.490 77.870 ;
        RECT 173.180 77.700 173.350 78.390 ;
        RECT 171.850 77.530 173.350 77.700 ;
        RECT 173.540 77.730 173.750 78.520 ;
        RECT 173.920 77.900 174.270 78.520 ;
        RECT 174.440 77.910 174.610 78.690 ;
        RECT 175.140 78.530 175.310 78.760 ;
        RECT 174.780 78.360 175.310 78.530 ;
        RECT 174.780 78.080 175.000 78.360 ;
        RECT 175.480 78.190 175.720 78.590 ;
        RECT 174.440 77.740 174.845 77.910 ;
        RECT 175.180 77.820 175.720 78.190 ;
        RECT 175.890 78.405 176.210 78.760 ;
        RECT 176.455 78.680 176.760 79.140 ;
        RECT 176.930 78.430 177.180 78.960 ;
        RECT 175.890 78.230 176.215 78.405 ;
        RECT 175.890 77.930 176.805 78.230 ;
        RECT 176.065 77.900 176.805 77.930 ;
        RECT 173.540 77.570 174.215 77.730 ;
        RECT 174.675 77.650 174.845 77.740 ;
        RECT 173.540 77.560 174.505 77.570 ;
        RECT 173.180 77.390 173.350 77.530 ;
        RECT 169.925 76.590 170.175 77.050 ;
        RECT 170.345 76.760 170.595 77.090 ;
        RECT 170.810 76.760 171.490 77.090 ;
        RECT 171.660 77.190 172.735 77.360 ;
        RECT 173.180 77.220 173.740 77.390 ;
        RECT 174.045 77.270 174.505 77.560 ;
        RECT 174.675 77.480 175.895 77.650 ;
        RECT 171.660 76.850 171.830 77.190 ;
        RECT 172.065 76.590 172.395 77.020 ;
        RECT 172.565 76.850 172.735 77.190 ;
        RECT 173.030 76.590 173.400 77.050 ;
        RECT 173.570 76.760 173.740 77.220 ;
        RECT 174.675 77.100 174.845 77.480 ;
        RECT 176.065 77.310 176.235 77.900 ;
        RECT 176.975 77.780 177.180 78.430 ;
        RECT 177.350 78.385 177.600 79.140 ;
        RECT 177.825 78.590 178.080 78.880 ;
        RECT 178.250 78.760 178.580 79.140 ;
        RECT 177.825 78.420 178.575 78.590 ;
        RECT 173.975 76.760 174.845 77.100 ;
        RECT 175.435 77.140 176.235 77.310 ;
        RECT 175.015 76.590 175.265 77.050 ;
        RECT 175.435 76.850 175.605 77.140 ;
        RECT 175.785 76.590 176.115 76.970 ;
        RECT 176.455 76.590 176.760 77.730 ;
        RECT 176.930 76.900 177.180 77.780 ;
        RECT 177.350 76.590 177.600 77.730 ;
        RECT 177.825 77.600 178.175 78.250 ;
        RECT 178.345 77.430 178.575 78.420 ;
        RECT 177.825 77.260 178.575 77.430 ;
        RECT 177.825 76.760 178.080 77.260 ;
        RECT 178.250 76.590 178.580 77.090 ;
        RECT 178.750 76.760 178.920 78.880 ;
        RECT 179.280 78.780 179.610 79.140 ;
        RECT 179.780 78.750 180.275 78.920 ;
        RECT 180.480 78.750 181.335 78.920 ;
        RECT 179.150 77.560 179.610 78.610 ;
        RECT 179.090 76.775 179.415 77.560 ;
        RECT 179.780 77.390 179.950 78.750 ;
        RECT 180.120 77.840 180.470 78.460 ;
        RECT 180.640 78.240 180.995 78.460 ;
        RECT 180.640 77.650 180.810 78.240 ;
        RECT 181.165 78.040 181.335 78.750 ;
        RECT 182.210 78.680 182.540 79.140 ;
        RECT 182.750 78.780 183.100 78.950 ;
        RECT 181.540 78.210 182.330 78.460 ;
        RECT 182.750 78.390 183.010 78.780 ;
        RECT 183.320 78.690 184.270 78.970 ;
        RECT 184.440 78.700 184.630 79.140 ;
        RECT 184.800 78.760 185.870 78.930 ;
        RECT 182.500 78.040 182.670 78.220 ;
        RECT 179.780 77.220 180.175 77.390 ;
        RECT 180.345 77.260 180.810 77.650 ;
        RECT 180.980 77.870 182.670 78.040 ;
        RECT 180.005 77.090 180.175 77.220 ;
        RECT 180.980 77.090 181.150 77.870 ;
        RECT 182.840 77.700 183.010 78.390 ;
        RECT 181.510 77.530 183.010 77.700 ;
        RECT 183.200 77.730 183.410 78.520 ;
        RECT 183.580 77.900 183.930 78.520 ;
        RECT 184.100 77.910 184.270 78.690 ;
        RECT 184.800 78.530 184.970 78.760 ;
        RECT 184.440 78.360 184.970 78.530 ;
        RECT 184.440 78.080 184.660 78.360 ;
        RECT 185.140 78.190 185.380 78.590 ;
        RECT 184.100 77.740 184.505 77.910 ;
        RECT 184.840 77.820 185.380 78.190 ;
        RECT 185.550 78.405 185.870 78.760 ;
        RECT 186.115 78.680 186.420 79.140 ;
        RECT 186.590 78.430 186.840 78.960 ;
        RECT 185.550 78.230 185.875 78.405 ;
        RECT 185.550 77.930 186.465 78.230 ;
        RECT 185.725 77.900 186.465 77.930 ;
        RECT 183.200 77.570 183.875 77.730 ;
        RECT 184.335 77.650 184.505 77.740 ;
        RECT 183.200 77.560 184.165 77.570 ;
        RECT 182.840 77.390 183.010 77.530 ;
        RECT 179.585 76.590 179.835 77.050 ;
        RECT 180.005 76.760 180.255 77.090 ;
        RECT 180.470 76.760 181.150 77.090 ;
        RECT 181.320 77.190 182.395 77.360 ;
        RECT 182.840 77.220 183.400 77.390 ;
        RECT 183.705 77.270 184.165 77.560 ;
        RECT 184.335 77.480 185.555 77.650 ;
        RECT 181.320 76.850 181.490 77.190 ;
        RECT 181.725 76.590 182.055 77.020 ;
        RECT 182.225 76.850 182.395 77.190 ;
        RECT 182.690 76.590 183.060 77.050 ;
        RECT 183.230 76.760 183.400 77.220 ;
        RECT 184.335 77.100 184.505 77.480 ;
        RECT 185.725 77.310 185.895 77.900 ;
        RECT 186.635 77.780 186.840 78.430 ;
        RECT 187.010 78.385 187.260 79.140 ;
        RECT 187.940 78.415 188.230 79.140 ;
        RECT 188.405 78.590 188.660 78.880 ;
        RECT 188.830 78.760 189.160 79.140 ;
        RECT 188.405 78.420 189.155 78.590 ;
        RECT 183.635 76.760 184.505 77.100 ;
        RECT 185.095 77.140 185.895 77.310 ;
        RECT 184.675 76.590 184.925 77.050 ;
        RECT 185.095 76.850 185.265 77.140 ;
        RECT 185.445 76.590 185.775 76.970 ;
        RECT 186.115 76.590 186.420 77.730 ;
        RECT 186.590 76.900 186.840 77.780 ;
        RECT 187.010 76.590 187.260 77.730 ;
        RECT 187.940 76.590 188.230 77.755 ;
        RECT 188.405 77.600 188.755 78.250 ;
        RECT 188.925 77.430 189.155 78.420 ;
        RECT 188.405 77.260 189.155 77.430 ;
        RECT 188.405 76.760 188.660 77.260 ;
        RECT 188.830 76.590 189.160 77.090 ;
        RECT 189.330 76.760 189.500 78.880 ;
        RECT 189.860 78.780 190.190 79.140 ;
        RECT 190.360 78.750 190.855 78.920 ;
        RECT 191.060 78.750 191.915 78.920 ;
        RECT 189.730 77.560 190.190 78.610 ;
        RECT 189.670 76.775 189.995 77.560 ;
        RECT 190.360 77.390 190.530 78.750 ;
        RECT 190.700 77.840 191.050 78.460 ;
        RECT 191.220 78.240 191.575 78.460 ;
        RECT 191.220 77.650 191.390 78.240 ;
        RECT 191.745 78.040 191.915 78.750 ;
        RECT 192.790 78.680 193.120 79.140 ;
        RECT 193.330 78.780 193.680 78.950 ;
        RECT 192.120 78.210 192.910 78.460 ;
        RECT 193.330 78.390 193.590 78.780 ;
        RECT 193.900 78.690 194.850 78.970 ;
        RECT 195.020 78.700 195.210 79.140 ;
        RECT 195.380 78.760 196.450 78.930 ;
        RECT 193.080 78.040 193.250 78.220 ;
        RECT 190.360 77.220 190.755 77.390 ;
        RECT 190.925 77.260 191.390 77.650 ;
        RECT 191.560 77.870 193.250 78.040 ;
        RECT 190.585 77.090 190.755 77.220 ;
        RECT 191.560 77.090 191.730 77.870 ;
        RECT 193.420 77.700 193.590 78.390 ;
        RECT 192.090 77.530 193.590 77.700 ;
        RECT 193.780 77.730 193.990 78.520 ;
        RECT 194.160 77.900 194.510 78.520 ;
        RECT 194.680 77.910 194.850 78.690 ;
        RECT 195.380 78.530 195.550 78.760 ;
        RECT 195.020 78.360 195.550 78.530 ;
        RECT 195.020 78.080 195.240 78.360 ;
        RECT 195.720 78.190 195.960 78.590 ;
        RECT 194.680 77.740 195.085 77.910 ;
        RECT 195.420 77.820 195.960 78.190 ;
        RECT 196.130 78.405 196.450 78.760 ;
        RECT 196.695 78.680 197.000 79.140 ;
        RECT 197.170 78.430 197.420 78.960 ;
        RECT 196.130 78.230 196.455 78.405 ;
        RECT 196.130 77.930 197.045 78.230 ;
        RECT 196.305 77.900 197.045 77.930 ;
        RECT 193.780 77.570 194.455 77.730 ;
        RECT 194.915 77.650 195.085 77.740 ;
        RECT 193.780 77.560 194.745 77.570 ;
        RECT 193.420 77.390 193.590 77.530 ;
        RECT 190.165 76.590 190.415 77.050 ;
        RECT 190.585 76.760 190.835 77.090 ;
        RECT 191.050 76.760 191.730 77.090 ;
        RECT 191.900 77.190 192.975 77.360 ;
        RECT 193.420 77.220 193.980 77.390 ;
        RECT 194.285 77.270 194.745 77.560 ;
        RECT 194.915 77.480 196.135 77.650 ;
        RECT 191.900 76.850 192.070 77.190 ;
        RECT 192.305 76.590 192.635 77.020 ;
        RECT 192.805 76.850 192.975 77.190 ;
        RECT 193.270 76.590 193.640 77.050 ;
        RECT 193.810 76.760 193.980 77.220 ;
        RECT 194.915 77.100 195.085 77.480 ;
        RECT 196.305 77.310 196.475 77.900 ;
        RECT 197.215 77.780 197.420 78.430 ;
        RECT 197.590 78.385 197.840 79.140 ;
        RECT 198.065 78.400 198.320 78.970 ;
        RECT 198.490 78.740 198.820 79.140 ;
        RECT 199.245 78.605 199.775 78.970 ;
        RECT 199.965 78.800 200.240 78.970 ;
        RECT 199.960 78.630 200.240 78.800 ;
        RECT 199.245 78.570 199.420 78.605 ;
        RECT 198.490 78.400 199.420 78.570 ;
        RECT 194.215 76.760 195.085 77.100 ;
        RECT 195.675 77.140 196.475 77.310 ;
        RECT 195.255 76.590 195.505 77.050 ;
        RECT 195.675 76.850 195.845 77.140 ;
        RECT 196.025 76.590 196.355 76.970 ;
        RECT 196.695 76.590 197.000 77.730 ;
        RECT 197.170 76.900 197.420 77.780 ;
        RECT 198.065 77.730 198.235 78.400 ;
        RECT 198.490 78.230 198.660 78.400 ;
        RECT 198.405 77.900 198.660 78.230 ;
        RECT 198.885 77.900 199.080 78.230 ;
        RECT 197.590 76.590 197.840 77.730 ;
        RECT 198.065 76.760 198.400 77.730 ;
        RECT 198.570 76.590 198.740 77.730 ;
        RECT 198.910 76.930 199.080 77.900 ;
        RECT 199.250 77.270 199.420 78.400 ;
        RECT 199.590 77.610 199.760 78.410 ;
        RECT 199.965 77.810 200.240 78.630 ;
        RECT 200.410 77.610 200.600 78.970 ;
        RECT 200.780 78.605 201.290 79.140 ;
        RECT 201.510 78.330 201.755 78.935 ;
        RECT 202.200 78.370 205.710 79.140 ;
        RECT 205.965 78.640 206.460 78.970 ;
        RECT 200.800 78.160 202.030 78.330 ;
        RECT 199.590 77.440 200.600 77.610 ;
        RECT 200.770 77.595 201.520 77.785 ;
        RECT 199.250 77.100 200.375 77.270 ;
        RECT 200.770 76.930 200.940 77.595 ;
        RECT 201.690 77.350 202.030 78.160 ;
        RECT 202.200 77.850 203.850 78.370 ;
        RECT 204.020 77.680 205.710 78.200 ;
        RECT 198.910 76.760 200.940 76.930 ;
        RECT 201.110 76.590 201.280 77.350 ;
        RECT 201.515 76.940 202.030 77.350 ;
        RECT 202.200 76.590 205.710 77.680 ;
        RECT 205.880 77.150 206.120 78.460 ;
        RECT 206.290 77.730 206.460 78.640 ;
        RECT 206.680 77.900 207.030 78.865 ;
        RECT 207.210 77.900 207.510 78.870 ;
        RECT 207.690 77.900 207.970 78.870 ;
        RECT 208.150 78.340 208.420 79.140 ;
        RECT 208.590 78.420 208.930 78.930 ;
        RECT 208.165 77.900 208.495 78.150 ;
        RECT 208.165 77.730 208.480 77.900 ;
        RECT 206.290 77.560 208.480 77.730 ;
        RECT 205.885 76.590 206.220 76.970 ;
        RECT 206.390 76.760 206.640 77.560 ;
        RECT 206.860 76.590 207.190 77.310 ;
        RECT 207.375 76.760 207.625 77.560 ;
        RECT 208.090 76.590 208.420 77.390 ;
        RECT 208.670 77.020 208.930 78.420 ;
        RECT 208.590 76.760 208.930 77.020 ;
        RECT 209.100 78.640 209.360 78.970 ;
        RECT 209.570 78.660 209.845 79.140 ;
        RECT 209.100 77.730 209.270 78.640 ;
        RECT 210.055 78.570 210.260 78.970 ;
        RECT 210.430 78.740 210.765 79.140 ;
        RECT 209.440 77.900 209.800 78.480 ;
        RECT 210.055 78.400 210.740 78.570 ;
        RECT 209.980 77.730 210.230 78.230 ;
        RECT 209.100 77.560 210.230 77.730 ;
        RECT 209.100 76.790 209.370 77.560 ;
        RECT 210.400 77.370 210.740 78.400 ;
        RECT 210.940 78.370 213.530 79.140 ;
        RECT 213.700 78.415 213.990 79.140 ;
        RECT 214.160 78.370 217.670 79.140 ;
        RECT 218.850 78.490 219.020 78.970 ;
        RECT 219.190 78.660 219.520 79.140 ;
        RECT 219.745 78.720 221.280 78.970 ;
        RECT 219.745 78.490 219.915 78.720 ;
        RECT 210.940 77.850 212.150 78.370 ;
        RECT 212.320 77.680 213.530 78.200 ;
        RECT 214.160 77.850 215.810 78.370 ;
        RECT 218.850 78.320 219.915 78.490 ;
        RECT 209.540 76.590 209.870 77.370 ;
        RECT 210.075 77.195 210.740 77.370 ;
        RECT 210.075 76.790 210.260 77.195 ;
        RECT 210.430 76.590 210.765 77.015 ;
        RECT 210.940 76.590 213.530 77.680 ;
        RECT 213.700 76.590 213.990 77.755 ;
        RECT 215.980 77.680 217.670 78.200 ;
        RECT 220.095 78.150 220.375 78.550 ;
        RECT 218.765 77.940 219.115 78.150 ;
        RECT 219.285 77.950 219.730 78.150 ;
        RECT 219.900 77.950 220.375 78.150 ;
        RECT 220.645 78.150 220.930 78.550 ;
        RECT 221.110 78.490 221.280 78.720 ;
        RECT 221.450 78.660 221.780 79.140 ;
        RECT 221.995 78.640 222.250 78.970 ;
        RECT 222.065 78.560 222.250 78.640 ;
        RECT 221.110 78.320 221.910 78.490 ;
        RECT 220.645 77.950 220.975 78.150 ;
        RECT 221.145 77.950 221.510 78.150 ;
        RECT 221.740 77.770 221.910 78.320 ;
        RECT 214.160 76.590 217.670 77.680 ;
        RECT 218.850 77.600 221.910 77.770 ;
        RECT 218.850 76.760 219.020 77.600 ;
        RECT 222.080 77.440 222.250 78.560 ;
        RECT 222.440 78.390 223.650 79.140 ;
        RECT 223.910 78.490 224.080 78.970 ;
        RECT 224.250 78.660 224.580 79.140 ;
        RECT 224.805 78.720 226.340 78.970 ;
        RECT 224.805 78.490 224.975 78.720 ;
        RECT 222.440 77.850 222.960 78.390 ;
        RECT 223.910 78.320 224.975 78.490 ;
        RECT 223.130 77.680 223.650 78.220 ;
        RECT 225.155 78.150 225.435 78.550 ;
        RECT 223.825 77.940 224.175 78.150 ;
        RECT 224.345 77.950 224.790 78.150 ;
        RECT 224.960 77.950 225.435 78.150 ;
        RECT 225.705 78.150 225.990 78.550 ;
        RECT 226.170 78.490 226.340 78.720 ;
        RECT 226.510 78.660 226.840 79.140 ;
        RECT 227.055 78.640 227.310 78.970 ;
        RECT 227.100 78.630 227.310 78.640 ;
        RECT 227.125 78.560 227.310 78.630 ;
        RECT 226.170 78.320 226.970 78.490 ;
        RECT 225.705 77.950 226.035 78.150 ;
        RECT 226.205 78.120 226.570 78.150 ;
        RECT 226.205 77.950 226.580 78.120 ;
        RECT 226.800 77.770 226.970 78.320 ;
        RECT 222.040 77.430 222.250 77.440 ;
        RECT 219.190 76.930 219.520 77.430 ;
        RECT 219.690 77.190 221.325 77.430 ;
        RECT 219.690 77.100 219.920 77.190 ;
        RECT 220.030 76.930 220.360 76.970 ;
        RECT 219.190 76.760 220.360 76.930 ;
        RECT 220.550 76.590 220.905 77.010 ;
        RECT 221.075 76.760 221.325 77.190 ;
        RECT 221.495 76.590 221.825 77.350 ;
        RECT 221.995 76.760 222.250 77.430 ;
        RECT 222.440 76.590 223.650 77.680 ;
        RECT 223.910 77.600 226.970 77.770 ;
        RECT 223.910 76.760 224.080 77.600 ;
        RECT 227.140 77.430 227.310 78.560 ;
        RECT 227.505 78.320 227.780 79.140 ;
        RECT 227.950 78.500 228.280 78.970 ;
        RECT 228.450 78.670 228.620 79.140 ;
        RECT 228.790 78.500 229.120 78.970 ;
        RECT 229.290 78.670 229.580 79.140 ;
        RECT 229.800 78.595 235.145 79.140 ;
        RECT 227.950 78.490 229.120 78.500 ;
        RECT 227.950 78.320 229.550 78.490 ;
        RECT 227.505 77.950 228.225 78.150 ;
        RECT 228.395 77.950 229.165 78.150 ;
        RECT 229.335 77.780 229.550 78.320 ;
        RECT 224.250 76.930 224.580 77.430 ;
        RECT 224.750 77.190 226.385 77.430 ;
        RECT 224.750 77.100 224.980 77.190 ;
        RECT 225.090 76.930 225.420 76.970 ;
        RECT 224.250 76.760 225.420 76.930 ;
        RECT 225.610 76.590 225.965 77.010 ;
        RECT 226.135 76.760 226.385 77.190 ;
        RECT 226.555 76.590 226.885 77.350 ;
        RECT 227.055 76.760 227.310 77.430 ;
        RECT 227.505 77.560 228.620 77.770 ;
        RECT 227.505 76.760 227.780 77.560 ;
        RECT 227.950 76.590 228.280 77.390 ;
        RECT 228.450 76.930 228.620 77.560 ;
        RECT 228.790 77.560 229.550 77.780 ;
        RECT 231.385 77.765 231.725 78.595 ;
        RECT 235.865 78.570 236.040 78.970 ;
        RECT 236.210 78.760 236.540 79.140 ;
        RECT 236.785 78.640 237.015 78.970 ;
        RECT 235.865 78.400 236.495 78.570 ;
        RECT 228.790 77.100 229.120 77.560 ;
        RECT 229.290 76.930 229.590 77.390 ;
        RECT 233.205 77.025 233.555 78.275 ;
        RECT 236.325 78.230 236.495 78.400 ;
        RECT 235.780 77.550 236.145 78.230 ;
        RECT 236.325 77.900 236.675 78.230 ;
        RECT 236.325 77.380 236.495 77.900 ;
        RECT 235.865 77.210 236.495 77.380 ;
        RECT 236.845 77.350 237.015 78.640 ;
        RECT 237.215 77.530 237.495 78.805 ;
        RECT 237.720 78.120 237.990 78.805 ;
        RECT 238.450 78.760 238.780 79.140 ;
        RECT 238.950 78.885 239.285 78.930 ;
        RECT 237.680 77.950 237.990 78.120 ;
        RECT 237.720 77.530 237.990 77.950 ;
        RECT 238.180 77.530 238.520 78.560 ;
        RECT 238.950 78.420 239.290 78.885 ;
        RECT 238.690 77.900 238.950 78.230 ;
        RECT 238.690 77.350 238.860 77.900 ;
        RECT 239.120 77.730 239.290 78.420 ;
        RECT 239.460 78.415 239.750 79.140 ;
        RECT 240.010 78.490 240.180 78.970 ;
        RECT 240.350 78.660 240.680 79.140 ;
        RECT 240.905 78.720 242.440 78.970 ;
        RECT 240.905 78.490 241.075 78.720 ;
        RECT 240.010 78.320 241.075 78.490 ;
        RECT 241.255 78.150 241.535 78.550 ;
        RECT 239.925 77.940 240.275 78.150 ;
        RECT 240.445 77.950 240.890 78.150 ;
        RECT 241.060 77.950 241.535 78.150 ;
        RECT 241.805 78.150 242.090 78.550 ;
        RECT 242.270 78.490 242.440 78.720 ;
        RECT 242.610 78.660 242.940 79.140 ;
        RECT 243.155 78.640 243.410 78.970 ;
        RECT 243.200 78.630 243.410 78.640 ;
        RECT 243.225 78.560 243.410 78.630 ;
        RECT 242.270 78.320 243.070 78.490 ;
        RECT 241.805 77.950 242.135 78.150 ;
        RECT 242.305 77.950 242.670 78.150 ;
        RECT 242.900 77.770 243.070 78.320 ;
        RECT 228.450 76.760 229.590 76.930 ;
        RECT 229.800 76.590 235.145 77.025 ;
        RECT 235.865 76.760 236.040 77.210 ;
        RECT 236.845 77.180 238.860 77.350 ;
        RECT 236.210 76.590 236.540 77.030 ;
        RECT 236.845 76.760 237.015 77.180 ;
        RECT 237.250 76.590 237.920 77.000 ;
        RECT 238.135 76.760 238.305 77.180 ;
        RECT 238.505 76.590 238.835 77.000 ;
        RECT 239.030 76.760 239.290 77.730 ;
        RECT 239.460 76.590 239.750 77.755 ;
        RECT 240.010 77.600 243.070 77.770 ;
        RECT 240.010 76.760 240.180 77.600 ;
        RECT 243.240 77.430 243.410 78.560 ;
        RECT 243.605 78.375 244.060 79.140 ;
        RECT 244.335 78.760 245.635 78.970 ;
        RECT 245.890 78.780 246.220 79.140 ;
        RECT 245.465 78.610 245.635 78.760 ;
        RECT 246.390 78.640 246.650 78.970 ;
        RECT 244.535 78.150 244.755 78.550 ;
        RECT 243.600 77.950 244.090 78.150 ;
        RECT 244.280 77.940 244.755 78.150 ;
        RECT 245.000 78.150 245.210 78.550 ;
        RECT 245.465 78.485 246.220 78.610 ;
        RECT 245.465 78.440 246.310 78.485 ;
        RECT 246.040 78.320 246.310 78.440 ;
        RECT 245.000 77.940 245.330 78.150 ;
        RECT 245.500 77.880 245.910 78.185 ;
        RECT 240.350 76.930 240.680 77.430 ;
        RECT 240.850 77.190 242.485 77.430 ;
        RECT 240.850 77.100 241.080 77.190 ;
        RECT 241.190 76.930 241.520 76.970 ;
        RECT 240.350 76.760 241.520 76.930 ;
        RECT 241.710 76.590 242.065 77.010 ;
        RECT 242.235 76.760 242.485 77.190 ;
        RECT 242.655 76.590 242.985 77.350 ;
        RECT 243.155 76.760 243.410 77.430 ;
        RECT 243.605 77.710 244.780 77.770 ;
        RECT 246.140 77.745 246.310 78.320 ;
        RECT 246.110 77.710 246.310 77.745 ;
        RECT 243.605 77.600 246.310 77.710 ;
        RECT 243.605 76.980 243.860 77.600 ;
        RECT 244.450 77.540 246.250 77.600 ;
        RECT 244.450 77.510 244.780 77.540 ;
        RECT 246.480 77.440 246.650 78.640 ;
        RECT 246.835 78.570 247.090 78.920 ;
        RECT 247.260 78.740 247.590 79.140 ;
        RECT 247.760 78.570 247.930 78.920 ;
        RECT 248.100 78.740 248.480 79.140 ;
        RECT 246.835 78.400 248.500 78.570 ;
        RECT 248.670 78.465 248.945 78.810 ;
        RECT 249.120 78.595 254.465 79.140 ;
        RECT 248.330 78.230 248.500 78.400 ;
        RECT 246.820 77.900 247.165 78.230 ;
        RECT 247.335 77.900 248.160 78.230 ;
        RECT 248.330 77.900 248.605 78.230 ;
        RECT 244.110 77.340 244.295 77.430 ;
        RECT 244.885 77.340 245.720 77.350 ;
        RECT 244.110 77.140 245.720 77.340 ;
        RECT 244.110 77.100 244.340 77.140 ;
        RECT 243.605 76.760 243.940 76.980 ;
        RECT 244.945 76.590 245.300 76.970 ;
        RECT 245.470 76.760 245.720 77.140 ;
        RECT 245.970 76.590 246.220 77.370 ;
        RECT 246.390 76.760 246.650 77.440 ;
        RECT 246.840 77.440 247.165 77.730 ;
        RECT 247.335 77.610 247.530 77.900 ;
        RECT 248.330 77.730 248.500 77.900 ;
        RECT 248.775 77.730 248.945 78.465 ;
        RECT 250.705 77.765 251.045 78.595 ;
        RECT 254.640 78.370 256.310 79.140 ;
        RECT 256.570 78.490 256.740 78.970 ;
        RECT 256.910 78.660 257.240 79.140 ;
        RECT 257.465 78.720 259.000 78.970 ;
        RECT 257.465 78.490 257.635 78.720 ;
        RECT 247.840 77.560 248.500 77.730 ;
        RECT 247.840 77.440 248.010 77.560 ;
        RECT 246.840 77.270 248.010 77.440 ;
        RECT 246.820 76.810 248.010 77.100 ;
        RECT 248.180 76.590 248.460 77.390 ;
        RECT 248.670 76.760 248.945 77.730 ;
        RECT 252.525 77.025 252.875 78.275 ;
        RECT 254.640 77.850 255.390 78.370 ;
        RECT 256.570 78.320 257.635 78.490 ;
        RECT 255.560 77.680 256.310 78.200 ;
        RECT 257.815 78.150 258.095 78.550 ;
        RECT 256.485 77.940 256.835 78.150 ;
        RECT 257.005 77.950 257.450 78.150 ;
        RECT 257.620 77.950 258.095 78.150 ;
        RECT 258.365 78.150 258.650 78.550 ;
        RECT 258.830 78.490 259.000 78.720 ;
        RECT 259.170 78.660 259.500 79.140 ;
        RECT 259.715 78.640 259.970 78.970 ;
        RECT 259.785 78.560 259.970 78.640 ;
        RECT 258.830 78.320 259.630 78.490 ;
        RECT 258.365 77.950 258.695 78.150 ;
        RECT 258.865 77.950 259.230 78.150 ;
        RECT 259.460 77.770 259.630 78.320 ;
        RECT 249.120 76.590 254.465 77.025 ;
        RECT 254.640 76.590 256.310 77.680 ;
        RECT 256.570 77.600 259.630 77.770 ;
        RECT 256.570 76.760 256.740 77.600 ;
        RECT 259.800 77.440 259.970 78.560 ;
        RECT 260.250 78.490 260.420 78.970 ;
        RECT 260.590 78.660 260.920 79.140 ;
        RECT 261.145 78.720 262.680 78.970 ;
        RECT 261.145 78.490 261.315 78.720 ;
        RECT 260.250 78.320 261.315 78.490 ;
        RECT 261.495 78.150 261.775 78.550 ;
        RECT 260.165 77.940 260.515 78.150 ;
        RECT 260.685 77.950 261.130 78.150 ;
        RECT 261.300 77.950 261.775 78.150 ;
        RECT 262.045 78.150 262.330 78.550 ;
        RECT 262.510 78.490 262.680 78.720 ;
        RECT 262.850 78.660 263.180 79.140 ;
        RECT 263.395 78.640 263.650 78.970 ;
        RECT 263.465 78.560 263.650 78.640 ;
        RECT 262.510 78.320 263.310 78.490 ;
        RECT 262.045 77.950 262.375 78.150 ;
        RECT 262.545 77.950 262.910 78.150 ;
        RECT 263.140 77.770 263.310 78.320 ;
        RECT 259.760 77.430 259.970 77.440 ;
        RECT 256.910 76.930 257.240 77.430 ;
        RECT 257.410 77.190 259.045 77.430 ;
        RECT 257.410 77.100 257.640 77.190 ;
        RECT 257.750 76.930 258.080 76.970 ;
        RECT 256.910 76.760 258.080 76.930 ;
        RECT 258.270 76.590 258.625 77.010 ;
        RECT 258.795 76.760 259.045 77.190 ;
        RECT 259.215 76.590 259.545 77.350 ;
        RECT 259.715 76.760 259.970 77.430 ;
        RECT 260.250 77.600 263.310 77.770 ;
        RECT 260.250 76.760 260.420 77.600 ;
        RECT 263.480 77.430 263.650 78.560 ;
        RECT 263.840 78.390 265.050 79.140 ;
        RECT 265.220 78.415 265.510 79.140 ;
        RECT 265.680 78.595 271.025 79.140 ;
        RECT 263.840 77.850 264.360 78.390 ;
        RECT 264.530 77.680 265.050 78.220 ;
        RECT 267.265 77.765 267.605 78.595 ;
        RECT 271.200 78.390 272.410 79.140 ;
        RECT 272.585 78.590 272.840 78.880 ;
        RECT 273.010 78.760 273.340 79.140 ;
        RECT 272.585 78.420 273.335 78.590 ;
        RECT 260.590 76.930 260.920 77.430 ;
        RECT 261.090 77.190 262.725 77.430 ;
        RECT 261.090 77.100 261.320 77.190 ;
        RECT 261.430 76.930 261.760 76.970 ;
        RECT 260.590 76.760 261.760 76.930 ;
        RECT 261.950 76.590 262.305 77.010 ;
        RECT 262.475 76.760 262.725 77.190 ;
        RECT 262.895 76.590 263.225 77.350 ;
        RECT 263.395 76.760 263.650 77.430 ;
        RECT 263.840 76.590 265.050 77.680 ;
        RECT 265.220 76.590 265.510 77.755 ;
        RECT 269.085 77.025 269.435 78.275 ;
        RECT 271.200 77.850 271.720 78.390 ;
        RECT 271.890 77.680 272.410 78.220 ;
        RECT 265.680 76.590 271.025 77.025 ;
        RECT 271.200 76.590 272.410 77.680 ;
        RECT 272.585 77.600 272.935 78.250 ;
        RECT 273.105 77.430 273.335 78.420 ;
        RECT 272.585 77.260 273.335 77.430 ;
        RECT 272.585 76.760 272.840 77.260 ;
        RECT 273.010 76.590 273.340 77.090 ;
        RECT 273.510 76.760 273.680 78.880 ;
        RECT 274.040 78.780 274.370 79.140 ;
        RECT 274.540 78.750 275.035 78.920 ;
        RECT 275.240 78.750 276.095 78.920 ;
        RECT 273.910 77.560 274.370 78.610 ;
        RECT 273.850 76.775 274.175 77.560 ;
        RECT 274.540 77.390 274.710 78.750 ;
        RECT 274.880 77.840 275.230 78.460 ;
        RECT 275.400 78.240 275.755 78.460 ;
        RECT 275.400 77.650 275.570 78.240 ;
        RECT 275.925 78.040 276.095 78.750 ;
        RECT 276.970 78.680 277.300 79.140 ;
        RECT 277.510 78.780 277.860 78.950 ;
        RECT 276.300 78.210 277.090 78.460 ;
        RECT 277.510 78.390 277.770 78.780 ;
        RECT 278.080 78.690 279.030 78.970 ;
        RECT 279.200 78.700 279.390 79.140 ;
        RECT 279.560 78.760 280.630 78.930 ;
        RECT 277.260 78.040 277.430 78.220 ;
        RECT 274.540 77.220 274.935 77.390 ;
        RECT 275.105 77.260 275.570 77.650 ;
        RECT 275.740 77.870 277.430 78.040 ;
        RECT 274.765 77.090 274.935 77.220 ;
        RECT 275.740 77.090 275.910 77.870 ;
        RECT 277.600 77.700 277.770 78.390 ;
        RECT 276.270 77.530 277.770 77.700 ;
        RECT 277.960 77.730 278.170 78.520 ;
        RECT 278.340 77.900 278.690 78.520 ;
        RECT 278.860 77.910 279.030 78.690 ;
        RECT 279.560 78.530 279.730 78.760 ;
        RECT 279.200 78.360 279.730 78.530 ;
        RECT 279.200 78.080 279.420 78.360 ;
        RECT 279.900 78.190 280.140 78.590 ;
        RECT 278.860 77.740 279.265 77.910 ;
        RECT 279.600 77.820 280.140 78.190 ;
        RECT 280.310 78.405 280.630 78.760 ;
        RECT 280.875 78.680 281.180 79.140 ;
        RECT 281.350 78.430 281.600 78.960 ;
        RECT 280.310 78.230 280.635 78.405 ;
        RECT 280.310 77.930 281.225 78.230 ;
        RECT 280.485 77.900 281.225 77.930 ;
        RECT 277.960 77.570 278.635 77.730 ;
        RECT 279.095 77.650 279.265 77.740 ;
        RECT 277.960 77.560 278.925 77.570 ;
        RECT 277.600 77.390 277.770 77.530 ;
        RECT 274.345 76.590 274.595 77.050 ;
        RECT 274.765 76.760 275.015 77.090 ;
        RECT 275.230 76.760 275.910 77.090 ;
        RECT 276.080 77.190 277.155 77.360 ;
        RECT 277.600 77.220 278.160 77.390 ;
        RECT 278.465 77.270 278.925 77.560 ;
        RECT 279.095 77.480 280.315 77.650 ;
        RECT 276.080 76.850 276.250 77.190 ;
        RECT 276.485 76.590 276.815 77.020 ;
        RECT 276.985 76.850 277.155 77.190 ;
        RECT 277.450 76.590 277.820 77.050 ;
        RECT 277.990 76.760 278.160 77.220 ;
        RECT 279.095 77.100 279.265 77.480 ;
        RECT 280.485 77.310 280.655 77.900 ;
        RECT 281.395 77.780 281.600 78.430 ;
        RECT 281.770 78.385 282.020 79.140 ;
        RECT 282.240 78.370 285.750 79.140 ;
        RECT 285.980 78.680 286.225 79.140 ;
        RECT 282.240 77.850 283.890 78.370 ;
        RECT 278.395 76.760 279.265 77.100 ;
        RECT 279.855 77.140 280.655 77.310 ;
        RECT 279.435 76.590 279.685 77.050 ;
        RECT 279.855 76.850 280.025 77.140 ;
        RECT 280.205 76.590 280.535 76.970 ;
        RECT 280.875 76.590 281.180 77.730 ;
        RECT 281.350 76.900 281.600 77.780 ;
        RECT 281.770 76.590 282.020 77.730 ;
        RECT 284.060 77.680 285.750 78.200 ;
        RECT 285.920 77.900 286.235 78.510 ;
        RECT 286.405 78.150 286.655 78.960 ;
        RECT 286.825 78.615 287.085 79.140 ;
        RECT 287.255 78.490 287.515 78.945 ;
        RECT 287.685 78.660 287.945 79.140 ;
        RECT 288.115 78.490 288.375 78.945 ;
        RECT 288.545 78.660 288.805 79.140 ;
        RECT 288.975 78.490 289.235 78.945 ;
        RECT 289.405 78.660 289.665 79.140 ;
        RECT 289.835 78.490 290.095 78.945 ;
        RECT 290.265 78.660 290.565 79.140 ;
        RECT 287.255 78.320 290.565 78.490 ;
        RECT 290.980 78.415 291.270 79.140 ;
        RECT 286.405 77.900 289.425 78.150 ;
        RECT 282.240 76.590 285.750 77.680 ;
        RECT 285.930 76.590 286.225 77.700 ;
        RECT 286.405 76.765 286.655 77.900 ;
        RECT 289.595 77.730 290.565 78.320 ;
        RECT 291.440 78.370 294.030 79.140 ;
        RECT 294.665 78.590 294.920 78.880 ;
        RECT 295.090 78.760 295.420 79.140 ;
        RECT 294.665 78.420 295.415 78.590 ;
        RECT 291.440 77.850 292.650 78.370 ;
        RECT 286.825 76.590 287.085 77.700 ;
        RECT 287.255 77.490 290.565 77.730 ;
        RECT 287.255 76.765 287.515 77.490 ;
        RECT 287.685 76.590 287.945 77.320 ;
        RECT 288.115 76.765 288.375 77.490 ;
        RECT 288.545 76.590 288.805 77.320 ;
        RECT 288.975 76.765 289.235 77.490 ;
        RECT 289.405 76.590 289.665 77.320 ;
        RECT 289.835 76.765 290.095 77.490 ;
        RECT 290.265 76.590 290.560 77.320 ;
        RECT 290.980 76.590 291.270 77.755 ;
        RECT 292.820 77.680 294.030 78.200 ;
        RECT 291.440 76.590 294.030 77.680 ;
        RECT 294.665 77.600 295.015 78.250 ;
        RECT 295.185 77.430 295.415 78.420 ;
        RECT 294.665 77.260 295.415 77.430 ;
        RECT 294.665 76.760 294.920 77.260 ;
        RECT 295.090 76.590 295.420 77.090 ;
        RECT 295.590 76.760 295.760 78.880 ;
        RECT 296.120 78.780 296.450 79.140 ;
        RECT 296.620 78.750 297.115 78.920 ;
        RECT 297.320 78.750 298.175 78.920 ;
        RECT 295.990 77.560 296.450 78.610 ;
        RECT 295.930 76.775 296.255 77.560 ;
        RECT 296.620 77.390 296.790 78.750 ;
        RECT 296.960 77.840 297.310 78.460 ;
        RECT 297.480 78.240 297.835 78.460 ;
        RECT 297.480 77.650 297.650 78.240 ;
        RECT 298.005 78.040 298.175 78.750 ;
        RECT 299.050 78.680 299.380 79.140 ;
        RECT 299.590 78.780 299.940 78.950 ;
        RECT 298.380 78.210 299.170 78.460 ;
        RECT 299.590 78.390 299.850 78.780 ;
        RECT 300.160 78.690 301.110 78.970 ;
        RECT 301.280 78.700 301.470 79.140 ;
        RECT 301.640 78.760 302.710 78.930 ;
        RECT 299.340 78.040 299.510 78.220 ;
        RECT 296.620 77.220 297.015 77.390 ;
        RECT 297.185 77.260 297.650 77.650 ;
        RECT 297.820 77.870 299.510 78.040 ;
        RECT 296.845 77.090 297.015 77.220 ;
        RECT 297.820 77.090 297.990 77.870 ;
        RECT 299.680 77.700 299.850 78.390 ;
        RECT 298.350 77.530 299.850 77.700 ;
        RECT 300.040 77.730 300.250 78.520 ;
        RECT 300.420 77.900 300.770 78.520 ;
        RECT 300.940 77.910 301.110 78.690 ;
        RECT 301.640 78.530 301.810 78.760 ;
        RECT 301.280 78.360 301.810 78.530 ;
        RECT 301.280 78.080 301.500 78.360 ;
        RECT 301.980 78.190 302.220 78.590 ;
        RECT 300.940 77.740 301.345 77.910 ;
        RECT 301.680 77.820 302.220 78.190 ;
        RECT 302.390 78.405 302.710 78.760 ;
        RECT 302.955 78.680 303.260 79.140 ;
        RECT 303.430 78.430 303.680 78.960 ;
        RECT 302.390 78.230 302.715 78.405 ;
        RECT 302.390 77.930 303.305 78.230 ;
        RECT 302.565 77.900 303.305 77.930 ;
        RECT 300.040 77.570 300.715 77.730 ;
        RECT 301.175 77.650 301.345 77.740 ;
        RECT 300.040 77.560 301.005 77.570 ;
        RECT 299.680 77.390 299.850 77.530 ;
        RECT 296.425 76.590 296.675 77.050 ;
        RECT 296.845 76.760 297.095 77.090 ;
        RECT 297.310 76.760 297.990 77.090 ;
        RECT 298.160 77.190 299.235 77.360 ;
        RECT 299.680 77.220 300.240 77.390 ;
        RECT 300.545 77.270 301.005 77.560 ;
        RECT 301.175 77.480 302.395 77.650 ;
        RECT 298.160 76.850 298.330 77.190 ;
        RECT 298.565 76.590 298.895 77.020 ;
        RECT 299.065 76.850 299.235 77.190 ;
        RECT 299.530 76.590 299.900 77.050 ;
        RECT 300.070 76.760 300.240 77.220 ;
        RECT 301.175 77.100 301.345 77.480 ;
        RECT 302.565 77.310 302.735 77.900 ;
        RECT 303.475 77.780 303.680 78.430 ;
        RECT 303.850 78.385 304.100 79.140 ;
        RECT 304.320 78.595 309.665 79.140 ;
        RECT 300.475 76.760 301.345 77.100 ;
        RECT 301.935 77.140 302.735 77.310 ;
        RECT 301.515 76.590 301.765 77.050 ;
        RECT 301.935 76.850 302.105 77.140 ;
        RECT 302.285 76.590 302.615 76.970 ;
        RECT 302.955 76.590 303.260 77.730 ;
        RECT 303.430 76.900 303.680 77.780 ;
        RECT 305.905 77.765 306.245 78.595 ;
        RECT 309.840 78.390 311.050 79.140 ;
        RECT 303.850 76.590 304.100 77.730 ;
        RECT 307.725 77.025 308.075 78.275 ;
        RECT 309.840 77.680 310.360 78.220 ;
        RECT 310.530 77.850 311.050 78.390 ;
        RECT 304.320 76.590 309.665 77.025 ;
        RECT 309.840 76.590 311.050 77.680 ;
        RECT 162.095 76.420 311.135 76.590 ;
        RECT 162.180 75.330 163.390 76.420 ;
        RECT 163.560 75.330 165.230 76.420 ;
        RECT 165.405 75.750 165.660 76.250 ;
        RECT 165.830 75.920 166.160 76.420 ;
        RECT 165.405 75.580 166.155 75.750 ;
        RECT 162.180 74.620 162.700 75.160 ;
        RECT 162.870 74.790 163.390 75.330 ;
        RECT 163.560 74.640 164.310 75.160 ;
        RECT 164.480 74.810 165.230 75.330 ;
        RECT 165.405 74.760 165.755 75.410 ;
        RECT 162.180 73.870 163.390 74.620 ;
        RECT 163.560 73.870 165.230 74.640 ;
        RECT 165.925 74.590 166.155 75.580 ;
        RECT 165.405 74.420 166.155 74.590 ;
        RECT 165.405 74.130 165.660 74.420 ;
        RECT 165.830 73.870 166.160 74.250 ;
        RECT 166.330 74.130 166.500 76.250 ;
        RECT 166.670 75.450 166.995 76.235 ;
        RECT 167.165 75.960 167.415 76.420 ;
        RECT 167.585 75.920 167.835 76.250 ;
        RECT 168.050 75.920 168.730 76.250 ;
        RECT 167.585 75.790 167.755 75.920 ;
        RECT 167.360 75.620 167.755 75.790 ;
        RECT 166.730 74.400 167.190 75.450 ;
        RECT 167.360 74.260 167.530 75.620 ;
        RECT 167.925 75.360 168.390 75.750 ;
        RECT 167.700 74.550 168.050 75.170 ;
        RECT 168.220 74.770 168.390 75.360 ;
        RECT 168.560 75.140 168.730 75.920 ;
        RECT 168.900 75.820 169.070 76.160 ;
        RECT 169.305 75.990 169.635 76.420 ;
        RECT 169.805 75.820 169.975 76.160 ;
        RECT 170.270 75.960 170.640 76.420 ;
        RECT 168.900 75.650 169.975 75.820 ;
        RECT 170.810 75.790 170.980 76.250 ;
        RECT 171.215 75.910 172.085 76.250 ;
        RECT 172.255 75.960 172.505 76.420 ;
        RECT 170.420 75.620 170.980 75.790 ;
        RECT 170.420 75.480 170.590 75.620 ;
        RECT 169.090 75.310 170.590 75.480 ;
        RECT 171.285 75.450 171.745 75.740 ;
        RECT 168.560 74.970 170.250 75.140 ;
        RECT 168.220 74.550 168.575 74.770 ;
        RECT 168.745 74.260 168.915 74.970 ;
        RECT 169.120 74.550 169.910 74.800 ;
        RECT 170.080 74.790 170.250 74.970 ;
        RECT 170.420 74.620 170.590 75.310 ;
        RECT 166.860 73.870 167.190 74.230 ;
        RECT 167.360 74.090 167.855 74.260 ;
        RECT 168.060 74.090 168.915 74.260 ;
        RECT 169.790 73.870 170.120 74.330 ;
        RECT 170.330 74.230 170.590 74.620 ;
        RECT 170.780 75.440 171.745 75.450 ;
        RECT 171.915 75.530 172.085 75.910 ;
        RECT 172.675 75.870 172.845 76.160 ;
        RECT 173.025 76.040 173.355 76.420 ;
        RECT 172.675 75.700 173.475 75.870 ;
        RECT 170.780 75.280 171.455 75.440 ;
        RECT 171.915 75.360 173.135 75.530 ;
        RECT 170.780 74.490 170.990 75.280 ;
        RECT 171.915 75.270 172.085 75.360 ;
        RECT 171.160 74.490 171.510 75.110 ;
        RECT 171.680 75.100 172.085 75.270 ;
        RECT 171.680 74.320 171.850 75.100 ;
        RECT 172.020 74.650 172.240 74.930 ;
        RECT 172.420 74.820 172.960 75.190 ;
        RECT 173.305 75.110 173.475 75.700 ;
        RECT 173.695 75.280 174.000 76.420 ;
        RECT 174.170 75.230 174.420 76.110 ;
        RECT 174.590 75.280 174.840 76.420 ;
        RECT 175.060 75.255 175.350 76.420 ;
        RECT 175.985 75.280 176.320 76.250 ;
        RECT 176.490 75.280 176.660 76.420 ;
        RECT 176.830 76.080 178.860 76.250 ;
        RECT 173.305 75.080 174.045 75.110 ;
        RECT 172.020 74.480 172.550 74.650 ;
        RECT 170.330 74.060 170.680 74.230 ;
        RECT 170.900 74.040 171.850 74.320 ;
        RECT 172.020 73.870 172.210 74.310 ;
        RECT 172.380 74.250 172.550 74.480 ;
        RECT 172.720 74.420 172.960 74.820 ;
        RECT 173.130 74.780 174.045 75.080 ;
        RECT 173.130 74.605 173.455 74.780 ;
        RECT 173.130 74.250 173.450 74.605 ;
        RECT 174.215 74.580 174.420 75.230 ;
        RECT 172.380 74.080 173.450 74.250 ;
        RECT 173.695 73.870 174.000 74.330 ;
        RECT 174.170 74.050 174.420 74.580 ;
        RECT 174.590 73.870 174.840 74.625 ;
        RECT 175.985 74.610 176.155 75.280 ;
        RECT 176.830 75.110 177.000 76.080 ;
        RECT 176.325 74.780 176.580 75.110 ;
        RECT 176.805 74.780 177.000 75.110 ;
        RECT 177.170 75.740 178.295 75.910 ;
        RECT 176.410 74.610 176.580 74.780 ;
        RECT 177.170 74.610 177.340 75.740 ;
        RECT 175.060 73.870 175.350 74.595 ;
        RECT 175.985 74.040 176.240 74.610 ;
        RECT 176.410 74.440 177.340 74.610 ;
        RECT 177.510 75.400 178.520 75.570 ;
        RECT 177.510 74.600 177.680 75.400 ;
        RECT 177.165 74.405 177.340 74.440 ;
        RECT 176.410 73.870 176.740 74.270 ;
        RECT 177.165 74.040 177.695 74.405 ;
        RECT 177.885 74.380 178.160 75.200 ;
        RECT 177.880 74.210 178.160 74.380 ;
        RECT 177.885 74.040 178.160 74.210 ;
        RECT 178.330 74.040 178.520 75.400 ;
        RECT 178.690 75.415 178.860 76.080 ;
        RECT 179.030 75.660 179.200 76.420 ;
        RECT 179.435 75.660 179.950 76.070 ;
        RECT 180.830 75.690 181.125 76.420 ;
        RECT 178.690 75.225 179.440 75.415 ;
        RECT 179.610 74.850 179.950 75.660 ;
        RECT 181.295 75.520 181.555 76.245 ;
        RECT 181.725 75.690 181.985 76.420 ;
        RECT 182.155 75.520 182.415 76.245 ;
        RECT 182.585 75.690 182.845 76.420 ;
        RECT 183.015 75.520 183.275 76.245 ;
        RECT 183.445 75.690 183.705 76.420 ;
        RECT 183.875 75.520 184.135 76.245 ;
        RECT 178.720 74.680 179.950 74.850 ;
        RECT 180.825 75.280 184.135 75.520 ;
        RECT 184.305 75.310 184.565 76.420 ;
        RECT 180.825 74.690 181.795 75.280 ;
        RECT 184.735 75.110 184.985 76.245 ;
        RECT 185.165 75.310 185.460 76.420 ;
        RECT 185.645 75.750 185.900 76.250 ;
        RECT 186.070 75.920 186.400 76.420 ;
        RECT 185.645 75.580 186.395 75.750 ;
        RECT 181.965 74.860 184.985 75.110 ;
        RECT 178.700 73.870 179.210 74.405 ;
        RECT 179.430 74.075 179.675 74.680 ;
        RECT 180.825 74.520 184.135 74.690 ;
        RECT 180.825 73.870 181.125 74.350 ;
        RECT 181.295 74.065 181.555 74.520 ;
        RECT 181.725 73.870 181.985 74.350 ;
        RECT 182.155 74.065 182.415 74.520 ;
        RECT 182.585 73.870 182.845 74.350 ;
        RECT 183.015 74.065 183.275 74.520 ;
        RECT 183.445 73.870 183.705 74.350 ;
        RECT 183.875 74.065 184.135 74.520 ;
        RECT 184.305 73.870 184.565 74.395 ;
        RECT 184.735 74.050 184.985 74.860 ;
        RECT 185.155 74.500 185.470 75.110 ;
        RECT 185.645 74.760 185.995 75.410 ;
        RECT 186.165 74.590 186.395 75.580 ;
        RECT 185.645 74.420 186.395 74.590 ;
        RECT 185.165 73.870 185.410 74.330 ;
        RECT 185.645 74.130 185.900 74.420 ;
        RECT 186.070 73.870 186.400 74.250 ;
        RECT 186.570 74.130 186.740 76.250 ;
        RECT 186.910 75.450 187.235 76.235 ;
        RECT 187.405 75.960 187.655 76.420 ;
        RECT 187.825 75.920 188.075 76.250 ;
        RECT 188.290 75.920 188.970 76.250 ;
        RECT 187.825 75.790 187.995 75.920 ;
        RECT 187.600 75.620 187.995 75.790 ;
        RECT 186.970 74.400 187.430 75.450 ;
        RECT 187.600 74.260 187.770 75.620 ;
        RECT 188.165 75.360 188.630 75.750 ;
        RECT 187.940 74.550 188.290 75.170 ;
        RECT 188.460 74.770 188.630 75.360 ;
        RECT 188.800 75.140 188.970 75.920 ;
        RECT 189.140 75.820 189.310 76.160 ;
        RECT 189.545 75.990 189.875 76.420 ;
        RECT 190.045 75.820 190.215 76.160 ;
        RECT 190.510 75.960 190.880 76.420 ;
        RECT 189.140 75.650 190.215 75.820 ;
        RECT 191.050 75.790 191.220 76.250 ;
        RECT 191.455 75.910 192.325 76.250 ;
        RECT 192.495 75.960 192.745 76.420 ;
        RECT 190.660 75.620 191.220 75.790 ;
        RECT 190.660 75.480 190.830 75.620 ;
        RECT 189.330 75.310 190.830 75.480 ;
        RECT 191.525 75.450 191.985 75.740 ;
        RECT 188.800 74.970 190.490 75.140 ;
        RECT 188.460 74.550 188.815 74.770 ;
        RECT 188.985 74.260 189.155 74.970 ;
        RECT 189.360 74.550 190.150 74.800 ;
        RECT 190.320 74.790 190.490 74.970 ;
        RECT 190.660 74.620 190.830 75.310 ;
        RECT 187.100 73.870 187.430 74.230 ;
        RECT 187.600 74.090 188.095 74.260 ;
        RECT 188.300 74.090 189.155 74.260 ;
        RECT 190.030 73.870 190.360 74.330 ;
        RECT 190.570 74.230 190.830 74.620 ;
        RECT 191.020 75.440 191.985 75.450 ;
        RECT 192.155 75.530 192.325 75.910 ;
        RECT 192.915 75.870 193.085 76.160 ;
        RECT 193.265 76.040 193.595 76.420 ;
        RECT 192.915 75.700 193.715 75.870 ;
        RECT 191.020 75.280 191.695 75.440 ;
        RECT 192.155 75.360 193.375 75.530 ;
        RECT 191.020 74.490 191.230 75.280 ;
        RECT 192.155 75.270 192.325 75.360 ;
        RECT 191.400 74.490 191.750 75.110 ;
        RECT 191.920 75.100 192.325 75.270 ;
        RECT 191.920 74.320 192.090 75.100 ;
        RECT 192.260 74.650 192.480 74.930 ;
        RECT 192.660 74.820 193.200 75.190 ;
        RECT 193.545 75.110 193.715 75.700 ;
        RECT 193.935 75.280 194.240 76.420 ;
        RECT 194.410 75.230 194.660 76.110 ;
        RECT 194.830 75.280 195.080 76.420 ;
        RECT 195.305 75.280 195.640 76.250 ;
        RECT 195.810 75.280 195.980 76.420 ;
        RECT 196.150 76.080 198.180 76.250 ;
        RECT 193.545 75.080 194.285 75.110 ;
        RECT 192.260 74.480 192.790 74.650 ;
        RECT 190.570 74.060 190.920 74.230 ;
        RECT 191.140 74.040 192.090 74.320 ;
        RECT 192.260 73.870 192.450 74.310 ;
        RECT 192.620 74.250 192.790 74.480 ;
        RECT 192.960 74.420 193.200 74.820 ;
        RECT 193.370 74.780 194.285 75.080 ;
        RECT 193.370 74.605 193.695 74.780 ;
        RECT 193.370 74.250 193.690 74.605 ;
        RECT 194.455 74.580 194.660 75.230 ;
        RECT 192.620 74.080 193.690 74.250 ;
        RECT 193.935 73.870 194.240 74.330 ;
        RECT 194.410 74.050 194.660 74.580 ;
        RECT 194.830 73.870 195.080 74.625 ;
        RECT 195.305 74.610 195.475 75.280 ;
        RECT 196.150 75.110 196.320 76.080 ;
        RECT 195.645 74.780 195.900 75.110 ;
        RECT 196.125 74.780 196.320 75.110 ;
        RECT 196.490 75.740 197.615 75.910 ;
        RECT 195.730 74.610 195.900 74.780 ;
        RECT 196.490 74.610 196.660 75.740 ;
        RECT 195.305 74.040 195.560 74.610 ;
        RECT 195.730 74.440 196.660 74.610 ;
        RECT 196.830 75.400 197.840 75.570 ;
        RECT 196.830 74.600 197.000 75.400 ;
        RECT 196.485 74.405 196.660 74.440 ;
        RECT 195.730 73.870 196.060 74.270 ;
        RECT 196.485 74.040 197.015 74.405 ;
        RECT 197.205 74.380 197.480 75.200 ;
        RECT 197.200 74.210 197.480 74.380 ;
        RECT 197.205 74.040 197.480 74.210 ;
        RECT 197.650 74.040 197.840 75.400 ;
        RECT 198.010 75.415 198.180 76.080 ;
        RECT 198.350 75.660 198.520 76.420 ;
        RECT 198.755 75.660 199.270 76.070 ;
        RECT 198.010 75.225 198.760 75.415 ;
        RECT 198.930 74.850 199.270 75.660 ;
        RECT 198.040 74.680 199.270 74.850 ;
        RECT 199.440 75.345 199.710 76.250 ;
        RECT 199.880 75.660 200.210 76.420 ;
        RECT 200.390 75.490 200.560 76.250 ;
        RECT 198.020 73.870 198.530 74.405 ;
        RECT 198.750 74.075 198.995 74.680 ;
        RECT 199.440 74.545 199.610 75.345 ;
        RECT 199.895 75.320 200.560 75.490 ;
        RECT 199.895 75.175 200.065 75.320 ;
        RECT 200.820 75.255 201.110 76.420 ;
        RECT 201.280 75.450 201.590 76.250 ;
        RECT 201.760 75.620 202.070 76.420 ;
        RECT 202.240 75.790 202.500 76.250 ;
        RECT 202.670 75.960 202.925 76.420 ;
        RECT 203.100 75.790 203.360 76.250 ;
        RECT 202.240 75.620 203.360 75.790 ;
        RECT 201.280 75.280 202.310 75.450 ;
        RECT 199.780 74.845 200.065 75.175 ;
        RECT 199.895 74.590 200.065 74.845 ;
        RECT 200.300 74.770 200.630 75.140 ;
        RECT 199.440 74.040 199.700 74.545 ;
        RECT 199.895 74.420 200.560 74.590 ;
        RECT 199.880 73.870 200.210 74.250 ;
        RECT 200.390 74.040 200.560 74.420 ;
        RECT 200.820 73.870 201.110 74.595 ;
        RECT 201.280 74.370 201.450 75.280 ;
        RECT 201.620 74.540 201.970 75.110 ;
        RECT 202.140 75.030 202.310 75.280 ;
        RECT 203.100 75.370 203.360 75.620 ;
        RECT 203.530 75.550 203.815 76.420 ;
        RECT 203.100 75.200 203.855 75.370 ;
        RECT 204.040 75.330 206.630 76.420 ;
        RECT 202.140 74.860 203.280 75.030 ;
        RECT 203.450 74.690 203.855 75.200 ;
        RECT 202.205 74.520 203.855 74.690 ;
        RECT 204.040 74.640 205.250 75.160 ;
        RECT 205.420 74.810 206.630 75.330 ;
        RECT 206.890 75.410 207.060 76.250 ;
        RECT 207.230 76.080 208.400 76.250 ;
        RECT 207.230 75.580 207.560 76.080 ;
        RECT 208.070 76.040 208.400 76.080 ;
        RECT 208.590 76.000 208.945 76.420 ;
        RECT 207.730 75.820 207.960 75.910 ;
        RECT 209.115 75.820 209.365 76.250 ;
        RECT 207.730 75.580 209.365 75.820 ;
        RECT 209.535 75.660 209.865 76.420 ;
        RECT 210.035 75.580 210.290 76.250 ;
        RECT 210.080 75.570 210.290 75.580 ;
        RECT 206.890 75.240 209.950 75.410 ;
        RECT 206.805 74.860 207.155 75.070 ;
        RECT 207.325 74.860 207.770 75.060 ;
        RECT 207.940 74.860 208.415 75.060 ;
        RECT 201.280 74.040 201.580 74.370 ;
        RECT 201.750 73.870 202.025 74.350 ;
        RECT 202.205 74.130 202.500 74.520 ;
        RECT 202.670 73.870 202.925 74.350 ;
        RECT 203.100 74.130 203.360 74.520 ;
        RECT 203.530 73.870 203.810 74.350 ;
        RECT 204.040 73.870 206.630 74.640 ;
        RECT 206.890 74.520 207.955 74.690 ;
        RECT 206.890 74.040 207.060 74.520 ;
        RECT 207.230 73.870 207.560 74.350 ;
        RECT 207.785 74.290 207.955 74.520 ;
        RECT 208.135 74.460 208.415 74.860 ;
        RECT 208.685 74.860 209.015 75.060 ;
        RECT 209.185 74.860 209.550 75.060 ;
        RECT 208.685 74.460 208.970 74.860 ;
        RECT 209.780 74.690 209.950 75.240 ;
        RECT 209.150 74.520 209.950 74.690 ;
        RECT 209.150 74.290 209.320 74.520 ;
        RECT 210.120 74.450 210.290 75.570 ;
        RECT 210.480 75.330 213.990 76.420 ;
        RECT 210.105 74.370 210.290 74.450 ;
        RECT 207.785 74.040 209.320 74.290 ;
        RECT 209.490 73.870 209.820 74.350 ;
        RECT 210.035 74.040 210.290 74.370 ;
        RECT 210.480 74.640 212.130 75.160 ;
        RECT 212.300 74.810 213.990 75.330 ;
        RECT 210.480 73.870 213.990 74.640 ;
        RECT 214.160 74.040 214.910 76.250 ;
        RECT 216.085 75.800 216.260 76.250 ;
        RECT 216.430 75.980 216.760 76.420 ;
        RECT 217.065 75.830 217.235 76.250 ;
        RECT 217.470 76.010 218.140 76.420 ;
        RECT 218.355 75.830 218.525 76.250 ;
        RECT 218.725 76.010 219.055 76.420 ;
        RECT 216.085 75.630 216.715 75.800 ;
        RECT 216.000 74.780 216.365 75.460 ;
        RECT 216.545 75.110 216.715 75.630 ;
        RECT 217.065 75.660 219.080 75.830 ;
        RECT 216.545 74.780 216.895 75.110 ;
        RECT 216.545 74.610 216.715 74.780 ;
        RECT 216.085 74.440 216.715 74.610 ;
        RECT 216.085 74.040 216.260 74.440 ;
        RECT 217.065 74.370 217.235 75.660 ;
        RECT 216.430 73.870 216.760 74.250 ;
        RECT 217.005 74.040 217.235 74.370 ;
        RECT 217.435 74.205 217.715 75.480 ;
        RECT 217.940 74.380 218.210 75.480 ;
        RECT 218.400 74.450 218.740 75.480 ;
        RECT 218.910 75.110 219.080 75.660 ;
        RECT 219.250 75.280 219.510 76.250 ;
        RECT 218.910 74.780 219.170 75.110 ;
        RECT 219.340 74.590 219.510 75.280 ;
        RECT 219.705 75.410 220.000 76.250 ;
        RECT 220.170 75.580 220.420 76.420 ;
        RECT 220.590 75.750 220.840 76.250 ;
        RECT 221.010 75.920 221.260 76.420 ;
        RECT 221.430 75.750 221.680 76.250 ;
        RECT 221.850 75.920 222.100 76.420 ;
        RECT 222.370 76.080 225.980 76.250 ;
        RECT 222.370 75.920 222.620 76.080 ;
        RECT 223.210 75.920 223.460 76.080 ;
        RECT 222.790 75.750 223.040 75.910 ;
        RECT 223.630 75.750 223.880 75.910 ;
        RECT 220.590 75.580 223.880 75.750 ;
        RECT 224.050 75.580 224.300 76.080 ;
        RECT 224.470 75.410 224.720 75.910 ;
        RECT 224.890 75.580 225.140 76.080 ;
        RECT 225.310 75.410 225.560 75.910 ;
        RECT 225.730 75.580 225.980 76.080 ;
        RECT 226.150 75.410 226.355 76.200 ;
        RECT 219.705 75.240 224.300 75.410 ;
        RECT 224.470 75.240 226.355 75.410 ;
        RECT 226.580 75.255 226.870 76.420 ;
        RECT 227.040 75.910 228.230 76.200 ;
        RECT 227.060 75.570 228.230 75.740 ;
        RECT 228.400 75.620 228.680 76.420 ;
        RECT 227.060 75.280 227.385 75.570 ;
        RECT 228.060 75.450 228.230 75.570 ;
        RECT 219.705 74.860 220.040 75.070 ;
        RECT 220.210 74.690 220.380 75.240 ;
        RECT 224.130 75.070 224.300 75.240 ;
        RECT 220.630 74.860 222.285 75.070 ;
        RECT 222.630 74.860 223.895 75.070 ;
        RECT 224.130 74.860 225.720 75.070 ;
        RECT 226.015 74.690 226.355 75.240 ;
        RECT 227.555 75.110 227.750 75.400 ;
        RECT 228.060 75.280 228.720 75.450 ;
        RECT 228.890 75.280 229.165 76.250 ;
        RECT 229.340 75.330 232.850 76.420 ;
        RECT 234.025 75.800 234.200 76.250 ;
        RECT 234.370 75.980 234.700 76.420 ;
        RECT 235.005 75.830 235.175 76.250 ;
        RECT 235.410 76.010 236.080 76.420 ;
        RECT 236.295 75.830 236.465 76.250 ;
        RECT 236.665 76.010 236.995 76.420 ;
        RECT 234.025 75.630 234.655 75.800 ;
        RECT 228.550 75.110 228.720 75.280 ;
        RECT 227.040 74.780 227.385 75.110 ;
        RECT 227.555 74.780 228.380 75.110 ;
        RECT 228.550 74.780 228.825 75.110 ;
        RECT 217.900 74.210 218.210 74.380 ;
        RECT 217.940 74.205 218.210 74.210 ;
        RECT 218.670 73.870 219.000 74.250 ;
        RECT 219.170 74.125 219.510 74.590 ;
        RECT 219.705 74.520 220.380 74.690 ;
        RECT 219.170 74.080 219.505 74.125 ;
        RECT 219.705 74.040 220.040 74.520 ;
        RECT 220.550 74.510 226.355 74.690 ;
        RECT 228.550 74.610 228.720 74.780 ;
        RECT 220.210 73.870 220.380 74.340 ;
        RECT 220.550 74.040 220.880 74.510 ;
        RECT 221.050 73.870 221.220 74.340 ;
        RECT 221.390 74.040 221.720 74.510 ;
        RECT 221.890 73.870 222.580 74.340 ;
        RECT 222.750 74.040 223.080 74.510 ;
        RECT 223.250 73.870 223.420 74.340 ;
        RECT 223.590 74.040 223.920 74.510 ;
        RECT 224.090 73.870 224.260 74.340 ;
        RECT 224.430 74.040 224.760 74.510 ;
        RECT 224.930 73.870 225.100 74.340 ;
        RECT 225.270 74.040 225.600 74.510 ;
        RECT 225.770 73.870 225.940 74.340 ;
        RECT 226.110 74.100 226.355 74.510 ;
        RECT 226.580 73.870 226.870 74.595 ;
        RECT 227.055 74.440 228.720 74.610 ;
        RECT 228.995 74.545 229.165 75.280 ;
        RECT 227.055 74.090 227.310 74.440 ;
        RECT 227.480 73.870 227.810 74.270 ;
        RECT 227.980 74.090 228.150 74.440 ;
        RECT 228.320 73.870 228.700 74.270 ;
        RECT 228.890 74.200 229.165 74.545 ;
        RECT 229.340 74.640 230.990 75.160 ;
        RECT 231.160 74.810 232.850 75.330 ;
        RECT 233.940 74.780 234.305 75.460 ;
        RECT 234.485 75.110 234.655 75.630 ;
        RECT 235.005 75.660 237.020 75.830 ;
        RECT 234.485 74.780 234.835 75.110 ;
        RECT 229.340 73.870 232.850 74.640 ;
        RECT 234.485 74.610 234.655 74.780 ;
        RECT 234.025 74.440 234.655 74.610 ;
        RECT 234.025 74.040 234.200 74.440 ;
        RECT 235.005 74.370 235.175 75.660 ;
        RECT 234.370 73.870 234.700 74.250 ;
        RECT 234.945 74.040 235.175 74.370 ;
        RECT 235.375 74.205 235.655 75.480 ;
        RECT 235.880 74.720 236.150 75.480 ;
        RECT 235.840 74.550 236.150 74.720 ;
        RECT 235.880 74.205 236.150 74.550 ;
        RECT 236.340 74.450 236.680 75.480 ;
        RECT 236.850 75.110 237.020 75.660 ;
        RECT 237.190 75.280 237.450 76.250 ;
        RECT 237.620 75.330 241.130 76.420 ;
        RECT 242.220 75.910 243.410 76.200 ;
        RECT 236.850 74.780 237.110 75.110 ;
        RECT 237.280 74.590 237.450 75.280 ;
        RECT 236.610 73.870 236.940 74.250 ;
        RECT 237.110 74.125 237.450 74.590 ;
        RECT 237.620 74.640 239.270 75.160 ;
        RECT 239.440 74.810 241.130 75.330 ;
        RECT 242.240 75.570 243.410 75.740 ;
        RECT 243.580 75.620 243.860 76.420 ;
        RECT 242.240 75.280 242.565 75.570 ;
        RECT 243.240 75.450 243.410 75.570 ;
        RECT 242.735 75.110 242.930 75.400 ;
        RECT 243.240 75.280 243.900 75.450 ;
        RECT 244.070 75.280 244.345 76.250 ;
        RECT 244.520 75.985 249.865 76.420 ;
        RECT 243.730 75.110 243.900 75.280 ;
        RECT 242.220 74.780 242.565 75.110 ;
        RECT 242.735 74.780 243.560 75.110 ;
        RECT 243.730 74.780 244.005 75.110 ;
        RECT 237.110 74.080 237.445 74.125 ;
        RECT 237.620 73.870 241.130 74.640 ;
        RECT 243.730 74.610 243.900 74.780 ;
        RECT 242.235 74.440 243.900 74.610 ;
        RECT 244.175 74.545 244.345 75.280 ;
        RECT 242.235 74.090 242.490 74.440 ;
        RECT 242.660 73.870 242.990 74.270 ;
        RECT 243.160 74.090 243.330 74.440 ;
        RECT 243.500 73.870 243.880 74.270 ;
        RECT 244.070 74.200 244.345 74.545 ;
        RECT 246.105 74.415 246.445 75.245 ;
        RECT 247.925 74.735 248.275 75.985 ;
        RECT 250.040 75.330 251.710 76.420 ;
        RECT 250.040 74.640 250.790 75.160 ;
        RECT 250.960 74.810 251.710 75.330 ;
        RECT 252.340 75.255 252.630 76.420 ;
        RECT 252.800 75.330 256.310 76.420 ;
        RECT 252.800 74.640 254.450 75.160 ;
        RECT 254.620 74.810 256.310 75.330 ;
        RECT 257.405 76.030 257.740 76.250 ;
        RECT 258.745 76.040 259.100 76.420 ;
        RECT 257.405 75.410 257.660 76.030 ;
        RECT 257.910 75.870 258.140 75.910 ;
        RECT 259.270 75.870 259.520 76.250 ;
        RECT 257.910 75.670 259.520 75.870 ;
        RECT 257.910 75.580 258.095 75.670 ;
        RECT 258.685 75.660 259.520 75.670 ;
        RECT 259.770 75.640 260.020 76.420 ;
        RECT 260.190 75.570 260.450 76.250 ;
        RECT 260.620 75.910 261.810 76.200 ;
        RECT 258.250 75.470 258.580 75.500 ;
        RECT 258.250 75.410 260.050 75.470 ;
        RECT 257.405 75.300 260.110 75.410 ;
        RECT 257.405 75.240 258.580 75.300 ;
        RECT 259.910 75.265 260.110 75.300 ;
        RECT 257.400 74.860 257.890 75.060 ;
        RECT 258.080 74.860 258.555 75.070 ;
        RECT 244.520 73.870 249.865 74.415 ;
        RECT 250.040 73.870 251.710 74.640 ;
        RECT 252.340 73.870 252.630 74.595 ;
        RECT 252.800 73.870 256.310 74.640 ;
        RECT 257.405 73.870 257.860 74.635 ;
        RECT 258.335 74.460 258.555 74.860 ;
        RECT 258.800 74.860 259.130 75.070 ;
        RECT 258.800 74.460 259.010 74.860 ;
        RECT 259.300 74.825 259.710 75.130 ;
        RECT 259.940 74.690 260.110 75.265 ;
        RECT 259.840 74.570 260.110 74.690 ;
        RECT 259.265 74.525 260.110 74.570 ;
        RECT 259.265 74.400 260.020 74.525 ;
        RECT 259.265 74.250 259.435 74.400 ;
        RECT 260.280 74.370 260.450 75.570 ;
        RECT 260.640 75.570 261.810 75.740 ;
        RECT 261.980 75.620 262.260 76.420 ;
        RECT 260.640 75.280 260.965 75.570 ;
        RECT 261.640 75.450 261.810 75.570 ;
        RECT 261.135 75.110 261.330 75.400 ;
        RECT 261.640 75.280 262.300 75.450 ;
        RECT 262.470 75.280 262.745 76.250 ;
        RECT 262.920 75.910 264.110 76.200 ;
        RECT 262.940 75.570 264.110 75.740 ;
        RECT 264.280 75.620 264.560 76.420 ;
        RECT 262.940 75.280 263.265 75.570 ;
        RECT 263.940 75.450 264.110 75.570 ;
        RECT 262.130 75.110 262.300 75.280 ;
        RECT 260.620 74.780 260.965 75.110 ;
        RECT 261.135 74.780 261.960 75.110 ;
        RECT 262.130 74.780 262.405 75.110 ;
        RECT 262.130 74.610 262.300 74.780 ;
        RECT 258.135 74.040 259.435 74.250 ;
        RECT 259.690 73.870 260.020 74.230 ;
        RECT 260.190 74.040 260.450 74.370 ;
        RECT 260.635 74.440 262.300 74.610 ;
        RECT 262.575 74.545 262.745 75.280 ;
        RECT 263.435 75.110 263.630 75.400 ;
        RECT 263.940 75.280 264.600 75.450 ;
        RECT 264.770 75.280 265.045 76.250 ;
        RECT 265.220 75.985 270.565 76.420 ;
        RECT 264.430 75.110 264.600 75.280 ;
        RECT 262.920 74.780 263.265 75.110 ;
        RECT 263.435 74.780 264.260 75.110 ;
        RECT 264.430 74.780 264.705 75.110 ;
        RECT 264.430 74.610 264.600 74.780 ;
        RECT 260.635 74.090 260.890 74.440 ;
        RECT 261.060 73.870 261.390 74.270 ;
        RECT 261.560 74.090 261.730 74.440 ;
        RECT 261.900 73.870 262.280 74.270 ;
        RECT 262.470 74.200 262.745 74.545 ;
        RECT 262.935 74.440 264.600 74.610 ;
        RECT 264.875 74.545 265.045 75.280 ;
        RECT 262.935 74.090 263.190 74.440 ;
        RECT 263.360 73.870 263.690 74.270 ;
        RECT 263.860 74.090 264.030 74.440 ;
        RECT 264.200 73.870 264.580 74.270 ;
        RECT 264.770 74.200 265.045 74.545 ;
        RECT 266.805 74.415 267.145 75.245 ;
        RECT 268.625 74.735 268.975 75.985 ;
        RECT 270.740 75.330 273.330 76.420 ;
        RECT 270.740 74.640 271.950 75.160 ;
        RECT 272.120 74.810 273.330 75.330 ;
        RECT 273.965 75.280 274.300 76.250 ;
        RECT 274.470 75.280 274.640 76.420 ;
        RECT 274.810 76.080 276.840 76.250 ;
        RECT 265.220 73.870 270.565 74.415 ;
        RECT 270.740 73.870 273.330 74.640 ;
        RECT 273.965 74.610 274.135 75.280 ;
        RECT 274.810 75.110 274.980 76.080 ;
        RECT 274.305 74.780 274.560 75.110 ;
        RECT 274.785 74.780 274.980 75.110 ;
        RECT 275.150 75.740 276.275 75.910 ;
        RECT 274.390 74.610 274.560 74.780 ;
        RECT 275.150 74.610 275.320 75.740 ;
        RECT 273.965 74.040 274.220 74.610 ;
        RECT 274.390 74.440 275.320 74.610 ;
        RECT 275.490 75.400 276.500 75.570 ;
        RECT 275.490 74.600 275.660 75.400 ;
        RECT 275.865 75.060 276.140 75.200 ;
        RECT 275.860 74.890 276.140 75.060 ;
        RECT 275.145 74.405 275.320 74.440 ;
        RECT 274.390 73.870 274.720 74.270 ;
        RECT 275.145 74.040 275.675 74.405 ;
        RECT 275.865 74.040 276.140 74.890 ;
        RECT 276.310 74.040 276.500 75.400 ;
        RECT 276.670 75.415 276.840 76.080 ;
        RECT 277.010 75.660 277.180 76.420 ;
        RECT 277.415 75.660 277.930 76.070 ;
        RECT 276.670 75.225 277.420 75.415 ;
        RECT 277.590 74.850 277.930 75.660 ;
        RECT 278.100 75.255 278.390 76.420 ;
        RECT 278.565 75.280 278.900 76.250 ;
        RECT 279.070 75.280 279.240 76.420 ;
        RECT 279.410 76.080 281.440 76.250 ;
        RECT 276.700 74.680 277.930 74.850 ;
        RECT 276.680 73.870 277.190 74.405 ;
        RECT 277.410 74.075 277.655 74.680 ;
        RECT 278.565 74.610 278.735 75.280 ;
        RECT 279.410 75.110 279.580 76.080 ;
        RECT 278.905 74.780 279.160 75.110 ;
        RECT 279.385 74.780 279.580 75.110 ;
        RECT 279.750 75.740 280.875 75.910 ;
        RECT 278.990 74.610 279.160 74.780 ;
        RECT 279.750 74.610 279.920 75.740 ;
        RECT 278.100 73.870 278.390 74.595 ;
        RECT 278.565 74.040 278.820 74.610 ;
        RECT 278.990 74.440 279.920 74.610 ;
        RECT 280.090 75.400 281.100 75.570 ;
        RECT 280.090 74.600 280.260 75.400 ;
        RECT 279.745 74.405 279.920 74.440 ;
        RECT 278.990 73.870 279.320 74.270 ;
        RECT 279.745 74.040 280.275 74.405 ;
        RECT 280.465 74.380 280.740 75.200 ;
        RECT 280.460 74.210 280.740 74.380 ;
        RECT 280.465 74.040 280.740 74.210 ;
        RECT 280.910 74.040 281.100 75.400 ;
        RECT 281.270 75.415 281.440 76.080 ;
        RECT 281.610 75.660 281.780 76.420 ;
        RECT 282.015 75.660 282.530 76.070 ;
        RECT 281.270 75.225 282.020 75.415 ;
        RECT 282.190 74.850 282.530 75.660 ;
        RECT 282.700 75.330 284.370 76.420 ;
        RECT 281.300 74.680 282.530 74.850 ;
        RECT 281.280 73.870 281.790 74.405 ;
        RECT 282.010 74.075 282.255 74.680 ;
        RECT 282.700 74.640 283.450 75.160 ;
        RECT 283.620 74.810 284.370 75.330 ;
        RECT 285.090 75.490 285.260 76.250 ;
        RECT 285.440 75.660 285.770 76.420 ;
        RECT 285.090 75.320 285.755 75.490 ;
        RECT 285.940 75.345 286.210 76.250 ;
        RECT 285.585 75.175 285.755 75.320 ;
        RECT 285.020 74.770 285.350 75.140 ;
        RECT 285.585 74.845 285.870 75.175 ;
        RECT 282.700 73.870 284.370 74.640 ;
        RECT 285.585 74.590 285.755 74.845 ;
        RECT 285.090 74.420 285.755 74.590 ;
        RECT 286.040 74.545 286.210 75.345 ;
        RECT 285.090 74.040 285.260 74.420 ;
        RECT 285.440 73.870 285.770 74.250 ;
        RECT 285.950 74.040 286.210 74.545 ;
        RECT 286.385 75.230 286.640 76.110 ;
        RECT 286.810 75.280 287.115 76.420 ;
        RECT 287.455 76.040 287.785 76.420 ;
        RECT 287.965 75.870 288.135 76.160 ;
        RECT 288.305 75.960 288.555 76.420 ;
        RECT 287.335 75.700 288.135 75.870 ;
        RECT 288.725 75.910 289.595 76.250 ;
        RECT 286.385 74.580 286.595 75.230 ;
        RECT 287.335 75.110 287.505 75.700 ;
        RECT 288.725 75.530 288.895 75.910 ;
        RECT 289.830 75.790 290.000 76.250 ;
        RECT 290.170 75.960 290.540 76.420 ;
        RECT 290.835 75.820 291.005 76.160 ;
        RECT 291.175 75.990 291.505 76.420 ;
        RECT 291.740 75.820 291.910 76.160 ;
        RECT 287.675 75.360 288.895 75.530 ;
        RECT 289.065 75.450 289.525 75.740 ;
        RECT 289.830 75.620 290.390 75.790 ;
        RECT 290.835 75.650 291.910 75.820 ;
        RECT 292.080 75.920 292.760 76.250 ;
        RECT 292.975 75.920 293.225 76.250 ;
        RECT 293.395 75.960 293.645 76.420 ;
        RECT 290.220 75.480 290.390 75.620 ;
        RECT 289.065 75.440 290.030 75.450 ;
        RECT 288.725 75.270 288.895 75.360 ;
        RECT 289.355 75.280 290.030 75.440 ;
        RECT 286.765 75.080 287.505 75.110 ;
        RECT 286.765 74.780 287.680 75.080 ;
        RECT 287.355 74.605 287.680 74.780 ;
        RECT 286.385 74.050 286.640 74.580 ;
        RECT 286.810 73.870 287.115 74.330 ;
        RECT 287.360 74.250 287.680 74.605 ;
        RECT 287.850 74.820 288.390 75.190 ;
        RECT 288.725 75.100 289.130 75.270 ;
        RECT 287.850 74.420 288.090 74.820 ;
        RECT 288.570 74.650 288.790 74.930 ;
        RECT 288.260 74.480 288.790 74.650 ;
        RECT 288.260 74.250 288.430 74.480 ;
        RECT 288.960 74.320 289.130 75.100 ;
        RECT 289.300 74.490 289.650 75.110 ;
        RECT 289.820 74.490 290.030 75.280 ;
        RECT 290.220 75.310 291.720 75.480 ;
        RECT 290.220 74.620 290.390 75.310 ;
        RECT 292.080 75.140 292.250 75.920 ;
        RECT 293.055 75.790 293.225 75.920 ;
        RECT 290.560 74.970 292.250 75.140 ;
        RECT 292.420 75.360 292.885 75.750 ;
        RECT 293.055 75.620 293.450 75.790 ;
        RECT 290.560 74.790 290.730 74.970 ;
        RECT 287.360 74.080 288.430 74.250 ;
        RECT 288.600 73.870 288.790 74.310 ;
        RECT 288.960 74.040 289.910 74.320 ;
        RECT 290.220 74.230 290.480 74.620 ;
        RECT 290.900 74.550 291.690 74.800 ;
        RECT 290.130 74.060 290.480 74.230 ;
        RECT 290.690 73.870 291.020 74.330 ;
        RECT 291.895 74.260 292.065 74.970 ;
        RECT 292.420 74.770 292.590 75.360 ;
        RECT 292.235 74.550 292.590 74.770 ;
        RECT 292.760 74.550 293.110 75.170 ;
        RECT 293.280 74.260 293.450 75.620 ;
        RECT 293.815 75.450 294.140 76.235 ;
        RECT 293.620 74.400 294.080 75.450 ;
        RECT 291.895 74.090 292.750 74.260 ;
        RECT 292.955 74.090 293.450 74.260 ;
        RECT 293.620 73.870 293.950 74.230 ;
        RECT 294.310 74.130 294.480 76.250 ;
        RECT 294.650 75.920 294.980 76.420 ;
        RECT 295.150 75.750 295.405 76.250 ;
        RECT 294.655 75.580 295.405 75.750 ;
        RECT 296.040 75.660 296.555 76.070 ;
        RECT 296.790 75.660 296.960 76.420 ;
        RECT 297.130 76.080 299.160 76.250 ;
        RECT 294.655 74.590 294.885 75.580 ;
        RECT 295.055 74.760 295.405 75.410 ;
        RECT 296.040 74.850 296.380 75.660 ;
        RECT 297.130 75.415 297.300 76.080 ;
        RECT 297.695 75.740 298.820 75.910 ;
        RECT 296.550 75.225 297.300 75.415 ;
        RECT 297.470 75.400 298.480 75.570 ;
        RECT 296.040 74.680 297.270 74.850 ;
        RECT 294.655 74.420 295.405 74.590 ;
        RECT 294.650 73.870 294.980 74.250 ;
        RECT 295.150 74.130 295.405 74.420 ;
        RECT 296.315 74.075 296.560 74.680 ;
        RECT 296.780 73.870 297.290 74.405 ;
        RECT 297.470 74.040 297.660 75.400 ;
        RECT 297.830 74.720 298.105 75.200 ;
        RECT 297.830 74.550 298.110 74.720 ;
        RECT 298.310 74.600 298.480 75.400 ;
        RECT 298.650 74.610 298.820 75.740 ;
        RECT 298.990 75.110 299.160 76.080 ;
        RECT 299.330 75.280 299.500 76.420 ;
        RECT 299.670 75.280 300.005 76.250 ;
        RECT 298.990 74.780 299.185 75.110 ;
        RECT 299.410 74.780 299.665 75.110 ;
        RECT 299.410 74.610 299.580 74.780 ;
        RECT 299.835 74.610 300.005 75.280 ;
        RECT 297.830 74.040 298.105 74.550 ;
        RECT 298.650 74.440 299.580 74.610 ;
        RECT 298.650 74.405 298.825 74.440 ;
        RECT 298.295 74.040 298.825 74.405 ;
        RECT 299.250 73.870 299.580 74.270 ;
        RECT 299.750 74.040 300.005 74.610 ;
        RECT 300.180 75.345 300.450 76.250 ;
        RECT 300.620 75.660 300.950 76.420 ;
        RECT 301.130 75.490 301.300 76.250 ;
        RECT 300.180 74.545 300.350 75.345 ;
        RECT 300.635 75.320 301.300 75.490 ;
        RECT 301.560 75.330 303.230 76.420 ;
        RECT 300.635 75.175 300.805 75.320 ;
        RECT 300.520 74.845 300.805 75.175 ;
        RECT 300.635 74.590 300.805 74.845 ;
        RECT 301.040 74.770 301.370 75.140 ;
        RECT 301.560 74.640 302.310 75.160 ;
        RECT 302.480 74.810 303.230 75.330 ;
        RECT 303.860 75.255 304.150 76.420 ;
        RECT 304.325 75.280 304.660 76.250 ;
        RECT 304.830 75.280 305.000 76.420 ;
        RECT 305.170 76.080 307.200 76.250 ;
        RECT 300.180 74.040 300.440 74.545 ;
        RECT 300.635 74.420 301.300 74.590 ;
        RECT 300.620 73.870 300.950 74.250 ;
        RECT 301.130 74.040 301.300 74.420 ;
        RECT 301.560 73.870 303.230 74.640 ;
        RECT 304.325 74.610 304.495 75.280 ;
        RECT 305.170 75.110 305.340 76.080 ;
        RECT 304.665 74.780 304.920 75.110 ;
        RECT 305.145 74.780 305.340 75.110 ;
        RECT 305.510 75.740 306.635 75.910 ;
        RECT 304.750 74.610 304.920 74.780 ;
        RECT 305.510 74.610 305.680 75.740 ;
        RECT 303.860 73.870 304.150 74.595 ;
        RECT 304.325 74.040 304.580 74.610 ;
        RECT 304.750 74.440 305.680 74.610 ;
        RECT 305.850 75.400 306.860 75.570 ;
        RECT 305.850 74.600 306.020 75.400 ;
        RECT 306.225 75.060 306.500 75.200 ;
        RECT 306.220 74.890 306.500 75.060 ;
        RECT 305.505 74.405 305.680 74.440 ;
        RECT 304.750 73.870 305.080 74.270 ;
        RECT 305.505 74.040 306.035 74.405 ;
        RECT 306.225 74.040 306.500 74.890 ;
        RECT 306.670 74.040 306.860 75.400 ;
        RECT 307.030 75.415 307.200 76.080 ;
        RECT 307.370 75.660 307.540 76.420 ;
        RECT 307.775 75.660 308.290 76.070 ;
        RECT 307.030 75.225 307.780 75.415 ;
        RECT 307.950 74.850 308.290 75.660 ;
        RECT 308.460 75.330 309.670 76.420 ;
        RECT 307.060 74.680 308.290 74.850 ;
        RECT 307.040 73.870 307.550 74.405 ;
        RECT 307.770 74.075 308.015 74.680 ;
        RECT 308.460 74.620 308.980 75.160 ;
        RECT 309.150 74.790 309.670 75.330 ;
        RECT 309.840 75.330 311.050 76.420 ;
        RECT 309.840 74.790 310.360 75.330 ;
        RECT 310.530 74.620 311.050 75.160 ;
        RECT 308.460 73.870 309.670 74.620 ;
        RECT 309.840 73.870 311.050 74.620 ;
        RECT 162.095 73.700 311.135 73.870 ;
        RECT 162.180 72.950 163.390 73.700 ;
        RECT 163.560 73.155 168.905 73.700 ;
        RECT 162.180 72.410 162.700 72.950 ;
        RECT 162.870 72.240 163.390 72.780 ;
        RECT 165.145 72.325 165.485 73.155 ;
        RECT 170.000 73.025 170.260 73.530 ;
        RECT 170.440 73.320 170.770 73.700 ;
        RECT 170.950 73.150 171.120 73.530 ;
        RECT 162.180 71.150 163.390 72.240 ;
        RECT 166.965 71.585 167.315 72.835 ;
        RECT 170.000 72.225 170.170 73.025 ;
        RECT 170.455 72.980 171.120 73.150 ;
        RECT 170.455 72.725 170.625 72.980 ;
        RECT 171.380 72.930 173.050 73.700 ;
        RECT 173.225 72.960 173.480 73.530 ;
        RECT 173.650 73.300 173.980 73.700 ;
        RECT 174.405 73.165 174.935 73.530 ;
        RECT 174.405 73.130 174.580 73.165 ;
        RECT 173.650 72.960 174.580 73.130 ;
        RECT 170.340 72.395 170.625 72.725 ;
        RECT 170.860 72.430 171.190 72.800 ;
        RECT 171.380 72.410 172.130 72.930 ;
        RECT 170.455 72.250 170.625 72.395 ;
        RECT 163.560 71.150 168.905 71.585 ;
        RECT 170.000 71.320 170.270 72.225 ;
        RECT 170.455 72.080 171.120 72.250 ;
        RECT 172.300 72.240 173.050 72.760 ;
        RECT 170.440 71.150 170.770 71.910 ;
        RECT 170.950 71.320 171.120 72.080 ;
        RECT 171.380 71.150 173.050 72.240 ;
        RECT 173.225 72.290 173.395 72.960 ;
        RECT 173.650 72.790 173.820 72.960 ;
        RECT 173.565 72.460 173.820 72.790 ;
        RECT 174.045 72.460 174.240 72.790 ;
        RECT 173.225 71.320 173.560 72.290 ;
        RECT 173.730 71.150 173.900 72.290 ;
        RECT 174.070 71.490 174.240 72.460 ;
        RECT 174.410 71.830 174.580 72.960 ;
        RECT 174.750 72.170 174.920 72.970 ;
        RECT 175.125 72.680 175.400 73.530 ;
        RECT 175.120 72.510 175.400 72.680 ;
        RECT 175.125 72.370 175.400 72.510 ;
        RECT 175.570 72.170 175.760 73.530 ;
        RECT 175.940 73.165 176.450 73.700 ;
        RECT 176.670 72.890 176.915 73.495 ;
        RECT 177.365 72.960 177.620 73.530 ;
        RECT 177.790 73.300 178.120 73.700 ;
        RECT 178.545 73.165 179.075 73.530 ;
        RECT 179.265 73.360 179.540 73.530 ;
        RECT 179.260 73.190 179.540 73.360 ;
        RECT 178.545 73.130 178.720 73.165 ;
        RECT 177.790 72.960 178.720 73.130 ;
        RECT 175.960 72.720 177.190 72.890 ;
        RECT 174.750 72.000 175.760 72.170 ;
        RECT 175.930 72.155 176.680 72.345 ;
        RECT 174.410 71.660 175.535 71.830 ;
        RECT 175.930 71.490 176.100 72.155 ;
        RECT 176.850 71.910 177.190 72.720 ;
        RECT 174.070 71.320 176.100 71.490 ;
        RECT 176.270 71.150 176.440 71.910 ;
        RECT 176.675 71.500 177.190 71.910 ;
        RECT 177.365 72.290 177.535 72.960 ;
        RECT 177.790 72.790 177.960 72.960 ;
        RECT 177.705 72.460 177.960 72.790 ;
        RECT 178.185 72.460 178.380 72.790 ;
        RECT 177.365 71.320 177.700 72.290 ;
        RECT 177.870 71.150 178.040 72.290 ;
        RECT 178.210 71.490 178.380 72.460 ;
        RECT 178.550 71.830 178.720 72.960 ;
        RECT 178.890 72.170 179.060 72.970 ;
        RECT 179.265 72.370 179.540 73.190 ;
        RECT 179.710 72.170 179.900 73.530 ;
        RECT 180.080 73.165 180.590 73.700 ;
        RECT 180.810 72.890 181.055 73.495 ;
        RECT 181.500 72.930 183.170 73.700 ;
        RECT 180.100 72.720 181.330 72.890 ;
        RECT 178.890 72.000 179.900 72.170 ;
        RECT 180.070 72.155 180.820 72.345 ;
        RECT 178.550 71.660 179.675 71.830 ;
        RECT 180.070 71.490 180.240 72.155 ;
        RECT 180.990 71.910 181.330 72.720 ;
        RECT 181.500 72.410 182.250 72.930 ;
        RECT 184.075 72.890 184.320 73.495 ;
        RECT 184.540 73.165 185.050 73.700 ;
        RECT 182.420 72.240 183.170 72.760 ;
        RECT 178.210 71.320 180.240 71.490 ;
        RECT 180.410 71.150 180.580 71.910 ;
        RECT 180.815 71.500 181.330 71.910 ;
        RECT 181.500 71.150 183.170 72.240 ;
        RECT 183.800 72.720 185.030 72.890 ;
        RECT 183.800 71.910 184.140 72.720 ;
        RECT 184.310 72.155 185.060 72.345 ;
        RECT 183.800 71.500 184.315 71.910 ;
        RECT 184.550 71.150 184.720 71.910 ;
        RECT 184.890 71.490 185.060 72.155 ;
        RECT 185.230 72.170 185.420 73.530 ;
        RECT 185.590 72.680 185.865 73.530 ;
        RECT 186.055 73.165 186.585 73.530 ;
        RECT 187.010 73.300 187.340 73.700 ;
        RECT 186.410 73.130 186.585 73.165 ;
        RECT 185.590 72.510 185.870 72.680 ;
        RECT 185.590 72.370 185.865 72.510 ;
        RECT 186.070 72.170 186.240 72.970 ;
        RECT 185.230 72.000 186.240 72.170 ;
        RECT 186.410 72.960 187.340 73.130 ;
        RECT 187.510 72.960 187.765 73.530 ;
        RECT 187.940 72.975 188.230 73.700 ;
        RECT 188.645 73.220 188.945 73.700 ;
        RECT 189.115 73.050 189.375 73.505 ;
        RECT 189.545 73.220 189.805 73.700 ;
        RECT 189.975 73.050 190.235 73.505 ;
        RECT 190.405 73.220 190.665 73.700 ;
        RECT 190.835 73.050 191.095 73.505 ;
        RECT 191.265 73.220 191.525 73.700 ;
        RECT 191.695 73.050 191.955 73.505 ;
        RECT 192.125 73.175 192.385 73.700 ;
        RECT 186.410 71.830 186.580 72.960 ;
        RECT 187.170 72.790 187.340 72.960 ;
        RECT 185.455 71.660 186.580 71.830 ;
        RECT 186.750 72.460 186.945 72.790 ;
        RECT 187.170 72.460 187.425 72.790 ;
        RECT 186.750 71.490 186.920 72.460 ;
        RECT 187.595 72.290 187.765 72.960 ;
        RECT 188.645 72.880 191.955 73.050 ;
        RECT 184.890 71.320 186.920 71.490 ;
        RECT 187.090 71.150 187.260 72.290 ;
        RECT 187.430 71.320 187.765 72.290 ;
        RECT 187.940 71.150 188.230 72.315 ;
        RECT 188.645 72.290 189.615 72.880 ;
        RECT 192.555 72.710 192.805 73.520 ;
        RECT 192.985 73.240 193.230 73.700 ;
        RECT 193.925 73.150 194.180 73.440 ;
        RECT 194.350 73.320 194.680 73.700 ;
        RECT 189.785 72.460 192.805 72.710 ;
        RECT 192.975 72.460 193.290 73.070 ;
        RECT 193.925 72.980 194.675 73.150 ;
        RECT 188.645 72.050 191.955 72.290 ;
        RECT 188.650 71.150 188.945 71.880 ;
        RECT 189.115 71.325 189.375 72.050 ;
        RECT 189.545 71.150 189.805 71.880 ;
        RECT 189.975 71.325 190.235 72.050 ;
        RECT 190.405 71.150 190.665 71.880 ;
        RECT 190.835 71.325 191.095 72.050 ;
        RECT 191.265 71.150 191.525 71.880 ;
        RECT 191.695 71.325 191.955 72.050 ;
        RECT 192.125 71.150 192.385 72.260 ;
        RECT 192.555 71.325 192.805 72.460 ;
        RECT 192.985 71.150 193.280 72.260 ;
        RECT 193.925 72.160 194.275 72.810 ;
        RECT 194.445 71.990 194.675 72.980 ;
        RECT 193.925 71.820 194.675 71.990 ;
        RECT 193.925 71.320 194.180 71.820 ;
        RECT 194.350 71.150 194.680 71.650 ;
        RECT 194.850 71.320 195.020 73.440 ;
        RECT 195.380 73.340 195.710 73.700 ;
        RECT 195.880 73.310 196.375 73.480 ;
        RECT 196.580 73.310 197.435 73.480 ;
        RECT 195.250 72.120 195.710 73.170 ;
        RECT 195.190 71.335 195.515 72.120 ;
        RECT 195.880 71.950 196.050 73.310 ;
        RECT 196.220 72.400 196.570 73.020 ;
        RECT 196.740 72.800 197.095 73.020 ;
        RECT 196.740 72.210 196.910 72.800 ;
        RECT 197.265 72.600 197.435 73.310 ;
        RECT 198.310 73.240 198.640 73.700 ;
        RECT 198.850 73.340 199.200 73.510 ;
        RECT 197.640 72.770 198.430 73.020 ;
        RECT 198.850 72.950 199.110 73.340 ;
        RECT 199.420 73.250 200.370 73.530 ;
        RECT 200.540 73.260 200.730 73.700 ;
        RECT 200.900 73.320 201.970 73.490 ;
        RECT 198.600 72.600 198.770 72.780 ;
        RECT 195.880 71.780 196.275 71.950 ;
        RECT 196.445 71.820 196.910 72.210 ;
        RECT 197.080 72.430 198.770 72.600 ;
        RECT 196.105 71.650 196.275 71.780 ;
        RECT 197.080 71.650 197.250 72.430 ;
        RECT 198.940 72.260 199.110 72.950 ;
        RECT 197.610 72.090 199.110 72.260 ;
        RECT 199.300 72.290 199.510 73.080 ;
        RECT 199.680 72.460 200.030 73.080 ;
        RECT 200.200 72.470 200.370 73.250 ;
        RECT 200.900 73.090 201.070 73.320 ;
        RECT 200.540 72.920 201.070 73.090 ;
        RECT 200.540 72.640 200.760 72.920 ;
        RECT 201.240 72.750 201.480 73.150 ;
        RECT 200.200 72.300 200.605 72.470 ;
        RECT 200.940 72.380 201.480 72.750 ;
        RECT 201.650 72.965 201.970 73.320 ;
        RECT 202.215 73.240 202.520 73.700 ;
        RECT 202.690 72.990 202.940 73.520 ;
        RECT 201.650 72.790 201.975 72.965 ;
        RECT 201.650 72.490 202.565 72.790 ;
        RECT 201.825 72.460 202.565 72.490 ;
        RECT 199.300 72.130 199.975 72.290 ;
        RECT 200.435 72.210 200.605 72.300 ;
        RECT 199.300 72.120 200.265 72.130 ;
        RECT 198.940 71.950 199.110 72.090 ;
        RECT 195.685 71.150 195.935 71.610 ;
        RECT 196.105 71.320 196.355 71.650 ;
        RECT 196.570 71.320 197.250 71.650 ;
        RECT 197.420 71.750 198.495 71.920 ;
        RECT 198.940 71.780 199.500 71.950 ;
        RECT 199.805 71.830 200.265 72.120 ;
        RECT 200.435 72.040 201.655 72.210 ;
        RECT 197.420 71.410 197.590 71.750 ;
        RECT 197.825 71.150 198.155 71.580 ;
        RECT 198.325 71.410 198.495 71.750 ;
        RECT 198.790 71.150 199.160 71.610 ;
        RECT 199.330 71.320 199.500 71.780 ;
        RECT 200.435 71.660 200.605 72.040 ;
        RECT 201.825 71.870 201.995 72.460 ;
        RECT 202.735 72.340 202.940 72.990 ;
        RECT 203.110 72.945 203.360 73.700 ;
        RECT 199.735 71.320 200.605 71.660 ;
        RECT 201.195 71.700 201.995 71.870 ;
        RECT 200.775 71.150 201.025 71.610 ;
        RECT 201.195 71.410 201.365 71.700 ;
        RECT 201.545 71.150 201.875 71.530 ;
        RECT 202.215 71.150 202.520 72.290 ;
        RECT 202.690 71.460 202.940 72.340 ;
        RECT 203.580 72.755 203.920 73.530 ;
        RECT 204.090 73.240 204.260 73.700 ;
        RECT 204.500 73.265 204.860 73.530 ;
        RECT 204.500 73.260 204.855 73.265 ;
        RECT 204.500 73.250 204.850 73.260 ;
        RECT 204.500 73.245 204.845 73.250 ;
        RECT 204.500 73.235 204.840 73.245 ;
        RECT 205.490 73.240 205.660 73.700 ;
        RECT 204.500 73.230 204.835 73.235 ;
        RECT 204.500 73.220 204.825 73.230 ;
        RECT 204.500 73.210 204.815 73.220 ;
        RECT 204.500 73.070 204.800 73.210 ;
        RECT 204.090 72.880 204.800 73.070 ;
        RECT 204.990 73.070 205.320 73.150 ;
        RECT 205.830 73.070 206.170 73.530 ;
        RECT 206.340 73.155 211.685 73.700 ;
        RECT 204.990 72.880 206.170 73.070 ;
        RECT 203.110 71.150 203.360 72.290 ;
        RECT 203.580 71.320 203.860 72.755 ;
        RECT 204.090 72.310 204.375 72.880 ;
        RECT 204.560 72.480 205.030 72.710 ;
        RECT 205.200 72.690 205.530 72.710 ;
        RECT 205.200 72.510 205.650 72.690 ;
        RECT 205.840 72.510 206.170 72.710 ;
        RECT 204.090 72.095 205.240 72.310 ;
        RECT 204.030 71.150 204.740 71.925 ;
        RECT 204.910 71.320 205.240 72.095 ;
        RECT 205.435 71.395 205.650 72.510 ;
        RECT 205.940 72.170 206.170 72.510 ;
        RECT 207.925 72.325 208.265 73.155 ;
        RECT 211.860 72.930 213.530 73.700 ;
        RECT 213.700 72.975 213.990 73.700 ;
        RECT 214.160 73.155 219.505 73.700 ;
        RECT 220.600 73.210 220.870 73.700 ;
        RECT 205.830 71.150 206.160 71.870 ;
        RECT 209.745 71.585 210.095 72.835 ;
        RECT 211.860 72.410 212.610 72.930 ;
        RECT 212.780 72.240 213.530 72.760 ;
        RECT 215.745 72.325 216.085 73.155 ;
        RECT 206.340 71.150 211.685 71.585 ;
        RECT 211.860 71.150 213.530 72.240 ;
        RECT 213.700 71.150 213.990 72.315 ;
        RECT 217.565 71.585 217.915 72.835 ;
        RECT 220.660 72.460 220.925 73.040 ;
        RECT 221.095 72.770 221.370 73.480 ;
        RECT 221.570 73.215 222.355 73.480 ;
        RECT 221.095 72.540 221.930 72.770 ;
        RECT 214.160 71.150 219.505 71.585 ;
        RECT 220.600 71.150 220.915 72.210 ;
        RECT 221.095 71.880 221.370 72.540 ;
        RECT 222.100 72.360 222.355 73.215 ;
        RECT 222.525 73.020 222.735 73.480 ;
        RECT 222.925 73.205 223.255 73.700 ;
        RECT 223.430 73.070 223.675 73.530 ;
        RECT 222.525 72.540 222.935 73.020 ;
        RECT 223.505 72.860 223.675 73.070 ;
        RECT 223.845 73.040 224.110 73.700 ;
        RECT 224.280 73.155 229.625 73.700 ;
        RECT 229.800 73.155 235.145 73.700 ;
        RECT 223.105 72.360 223.335 72.790 ;
        RECT 221.565 72.190 223.335 72.360 ;
        RECT 223.505 72.340 224.110 72.860 ;
        RECT 221.565 71.825 221.800 72.190 ;
        RECT 221.970 71.830 222.300 72.020 ;
        RECT 222.525 71.895 222.715 72.190 ;
        RECT 221.970 71.655 222.160 71.830 ;
        RECT 221.545 71.150 222.160 71.655 ;
        RECT 222.330 71.320 222.805 71.660 ;
        RECT 222.975 71.150 223.190 71.995 ;
        RECT 223.505 71.990 223.675 72.340 ;
        RECT 225.865 72.325 226.205 73.155 ;
        RECT 223.390 71.320 223.675 71.990 ;
        RECT 223.845 71.150 224.110 72.160 ;
        RECT 227.685 71.585 228.035 72.835 ;
        RECT 231.385 72.325 231.725 73.155 ;
        RECT 235.320 72.930 238.830 73.700 ;
        RECT 239.460 72.975 239.750 73.700 ;
        RECT 240.010 73.050 240.180 73.530 ;
        RECT 240.350 73.220 240.680 73.700 ;
        RECT 240.905 73.280 242.440 73.530 ;
        RECT 240.905 73.050 241.075 73.280 ;
        RECT 233.205 71.585 233.555 72.835 ;
        RECT 235.320 72.410 236.970 72.930 ;
        RECT 240.010 72.880 241.075 73.050 ;
        RECT 237.140 72.240 238.830 72.760 ;
        RECT 241.255 72.710 241.535 73.110 ;
        RECT 239.925 72.500 240.275 72.710 ;
        RECT 240.445 72.510 240.890 72.710 ;
        RECT 241.060 72.510 241.535 72.710 ;
        RECT 241.805 72.710 242.090 73.110 ;
        RECT 242.270 73.050 242.440 73.280 ;
        RECT 242.610 73.220 242.940 73.700 ;
        RECT 243.155 73.200 243.410 73.530 ;
        RECT 243.200 73.190 243.410 73.200 ;
        RECT 243.225 73.120 243.410 73.190 ;
        RECT 243.600 73.155 248.945 73.700 ;
        RECT 249.120 73.155 254.465 73.700 ;
        RECT 242.270 72.880 243.070 73.050 ;
        RECT 241.805 72.510 242.135 72.710 ;
        RECT 242.305 72.680 242.670 72.710 ;
        RECT 242.305 72.510 242.680 72.680 ;
        RECT 242.900 72.330 243.070 72.880 ;
        RECT 224.280 71.150 229.625 71.585 ;
        RECT 229.800 71.150 235.145 71.585 ;
        RECT 235.320 71.150 238.830 72.240 ;
        RECT 239.460 71.150 239.750 72.315 ;
        RECT 240.010 72.160 243.070 72.330 ;
        RECT 240.010 71.320 240.180 72.160 ;
        RECT 243.240 71.990 243.410 73.120 ;
        RECT 245.185 72.325 245.525 73.155 ;
        RECT 240.350 71.490 240.680 71.990 ;
        RECT 240.850 71.750 242.485 71.990 ;
        RECT 240.850 71.660 241.080 71.750 ;
        RECT 241.190 71.490 241.520 71.530 ;
        RECT 240.350 71.320 241.520 71.490 ;
        RECT 241.710 71.150 242.065 71.570 ;
        RECT 242.235 71.320 242.485 71.750 ;
        RECT 242.655 71.150 242.985 71.910 ;
        RECT 243.155 71.320 243.410 71.990 ;
        RECT 247.005 71.585 247.355 72.835 ;
        RECT 250.705 72.325 251.045 73.155 ;
        RECT 255.190 73.050 255.360 73.530 ;
        RECT 255.530 73.220 255.860 73.700 ;
        RECT 256.085 73.280 257.620 73.530 ;
        RECT 256.085 73.050 256.255 73.280 ;
        RECT 255.190 72.880 256.255 73.050 ;
        RECT 252.525 71.585 252.875 72.835 ;
        RECT 256.435 72.710 256.715 73.110 ;
        RECT 255.105 72.500 255.455 72.710 ;
        RECT 255.625 72.510 256.070 72.710 ;
        RECT 256.240 72.510 256.715 72.710 ;
        RECT 256.985 72.710 257.270 73.110 ;
        RECT 257.450 73.050 257.620 73.280 ;
        RECT 257.790 73.220 258.120 73.700 ;
        RECT 258.335 73.200 258.590 73.530 ;
        RECT 258.380 73.190 258.590 73.200 ;
        RECT 258.405 73.120 258.590 73.190 ;
        RECT 258.780 73.155 264.125 73.700 ;
        RECT 257.450 72.880 258.250 73.050 ;
        RECT 256.985 72.510 257.315 72.710 ;
        RECT 257.485 72.510 257.850 72.710 ;
        RECT 258.080 72.330 258.250 72.880 ;
        RECT 255.190 72.160 258.250 72.330 ;
        RECT 243.600 71.150 248.945 71.585 ;
        RECT 249.120 71.150 254.465 71.585 ;
        RECT 255.190 71.320 255.360 72.160 ;
        RECT 258.420 71.990 258.590 73.120 ;
        RECT 260.365 72.325 260.705 73.155 ;
        RECT 265.220 72.975 265.510 73.700 ;
        RECT 265.680 73.155 271.025 73.700 ;
        RECT 271.200 73.155 276.545 73.700 ;
        RECT 255.530 71.490 255.860 71.990 ;
        RECT 256.030 71.750 257.665 71.990 ;
        RECT 256.030 71.660 256.260 71.750 ;
        RECT 256.370 71.490 256.700 71.530 ;
        RECT 255.530 71.320 256.700 71.490 ;
        RECT 256.890 71.150 257.245 71.570 ;
        RECT 257.415 71.320 257.665 71.750 ;
        RECT 257.835 71.150 258.165 71.910 ;
        RECT 258.335 71.320 258.590 71.990 ;
        RECT 262.185 71.585 262.535 72.835 ;
        RECT 267.265 72.325 267.605 73.155 ;
        RECT 258.780 71.150 264.125 71.585 ;
        RECT 265.220 71.150 265.510 72.315 ;
        RECT 269.085 71.585 269.435 72.835 ;
        RECT 272.785 72.325 273.125 73.155 ;
        RECT 276.720 72.930 278.390 73.700 ;
        RECT 278.560 73.070 278.900 73.530 ;
        RECT 279.070 73.240 279.240 73.700 ;
        RECT 279.870 73.265 280.230 73.530 ;
        RECT 279.875 73.260 280.230 73.265 ;
        RECT 279.880 73.250 280.230 73.260 ;
        RECT 279.885 73.245 280.230 73.250 ;
        RECT 279.890 73.235 280.230 73.245 ;
        RECT 280.470 73.240 280.640 73.700 ;
        RECT 279.895 73.230 280.230 73.235 ;
        RECT 279.905 73.220 280.230 73.230 ;
        RECT 279.915 73.210 280.230 73.220 ;
        RECT 279.410 73.070 279.740 73.150 ;
        RECT 274.605 71.585 274.955 72.835 ;
        RECT 276.720 72.410 277.470 72.930 ;
        RECT 278.560 72.880 279.740 73.070 ;
        RECT 279.930 73.070 280.230 73.210 ;
        RECT 279.930 72.880 280.640 73.070 ;
        RECT 277.640 72.240 278.390 72.760 ;
        RECT 265.680 71.150 271.025 71.585 ;
        RECT 271.200 71.150 276.545 71.585 ;
        RECT 276.720 71.150 278.390 72.240 ;
        RECT 278.560 72.510 278.890 72.710 ;
        RECT 279.200 72.690 279.530 72.710 ;
        RECT 279.080 72.510 279.530 72.690 ;
        RECT 278.560 72.170 278.790 72.510 ;
        RECT 278.570 71.150 278.900 71.870 ;
        RECT 279.080 71.395 279.295 72.510 ;
        RECT 279.700 72.480 280.170 72.710 ;
        RECT 280.355 72.310 280.640 72.880 ;
        RECT 280.810 72.755 281.150 73.530 ;
        RECT 279.490 72.095 280.640 72.310 ;
        RECT 279.490 71.320 279.820 72.095 ;
        RECT 279.990 71.150 280.700 71.925 ;
        RECT 280.870 71.320 281.150 72.755 ;
        RECT 281.320 72.930 284.830 73.700 ;
        RECT 285.980 73.240 286.225 73.700 ;
        RECT 281.320 72.410 282.970 72.930 ;
        RECT 283.140 72.240 284.830 72.760 ;
        RECT 285.920 72.460 286.235 73.070 ;
        RECT 286.405 72.710 286.655 73.520 ;
        RECT 286.825 73.175 287.085 73.700 ;
        RECT 287.255 73.050 287.515 73.505 ;
        RECT 287.685 73.220 287.945 73.700 ;
        RECT 288.115 73.050 288.375 73.505 ;
        RECT 288.545 73.220 288.805 73.700 ;
        RECT 288.975 73.050 289.235 73.505 ;
        RECT 289.405 73.220 289.665 73.700 ;
        RECT 289.835 73.050 290.095 73.505 ;
        RECT 290.265 73.220 290.565 73.700 ;
        RECT 287.255 72.880 290.565 73.050 ;
        RECT 290.980 72.975 291.270 73.700 ;
        RECT 286.405 72.460 289.425 72.710 ;
        RECT 281.320 71.150 284.830 72.240 ;
        RECT 285.930 71.150 286.225 72.260 ;
        RECT 286.405 71.325 286.655 72.460 ;
        RECT 289.595 72.290 290.565 72.880 ;
        RECT 291.440 72.930 293.110 73.700 ;
        RECT 293.830 73.150 294.000 73.530 ;
        RECT 294.180 73.320 294.510 73.700 ;
        RECT 293.830 72.980 294.495 73.150 ;
        RECT 294.690 73.025 294.950 73.530 ;
        RECT 291.440 72.410 292.190 72.930 ;
        RECT 286.825 71.150 287.085 72.260 ;
        RECT 287.255 72.050 290.565 72.290 ;
        RECT 287.255 71.325 287.515 72.050 ;
        RECT 287.685 71.150 287.945 71.880 ;
        RECT 288.115 71.325 288.375 72.050 ;
        RECT 288.545 71.150 288.805 71.880 ;
        RECT 288.975 71.325 289.235 72.050 ;
        RECT 289.405 71.150 289.665 71.880 ;
        RECT 289.835 71.325 290.095 72.050 ;
        RECT 290.265 71.150 290.560 71.880 ;
        RECT 290.980 71.150 291.270 72.315 ;
        RECT 292.360 72.240 293.110 72.760 ;
        RECT 293.760 72.430 294.090 72.800 ;
        RECT 294.325 72.725 294.495 72.980 ;
        RECT 294.325 72.395 294.610 72.725 ;
        RECT 294.325 72.250 294.495 72.395 ;
        RECT 291.440 71.150 293.110 72.240 ;
        RECT 293.830 72.080 294.495 72.250 ;
        RECT 294.780 72.225 294.950 73.025 ;
        RECT 295.125 73.150 295.380 73.440 ;
        RECT 295.550 73.320 295.880 73.700 ;
        RECT 295.125 72.980 295.875 73.150 ;
        RECT 293.830 71.320 294.000 72.080 ;
        RECT 294.180 71.150 294.510 71.910 ;
        RECT 294.680 71.320 294.950 72.225 ;
        RECT 295.125 72.160 295.475 72.810 ;
        RECT 295.645 71.990 295.875 72.980 ;
        RECT 295.125 71.820 295.875 71.990 ;
        RECT 295.125 71.320 295.380 71.820 ;
        RECT 295.550 71.150 295.880 71.650 ;
        RECT 296.050 71.320 296.220 73.440 ;
        RECT 296.580 73.340 296.910 73.700 ;
        RECT 297.080 73.310 297.575 73.480 ;
        RECT 297.780 73.310 298.635 73.480 ;
        RECT 296.450 72.120 296.910 73.170 ;
        RECT 296.390 71.335 296.715 72.120 ;
        RECT 297.080 71.950 297.250 73.310 ;
        RECT 297.420 72.400 297.770 73.020 ;
        RECT 297.940 72.800 298.295 73.020 ;
        RECT 297.940 72.210 298.110 72.800 ;
        RECT 298.465 72.600 298.635 73.310 ;
        RECT 299.510 73.240 299.840 73.700 ;
        RECT 300.050 73.340 300.400 73.510 ;
        RECT 298.840 72.770 299.630 73.020 ;
        RECT 300.050 72.950 300.310 73.340 ;
        RECT 300.620 73.250 301.570 73.530 ;
        RECT 301.740 73.260 301.930 73.700 ;
        RECT 302.100 73.320 303.170 73.490 ;
        RECT 299.800 72.600 299.970 72.780 ;
        RECT 297.080 71.780 297.475 71.950 ;
        RECT 297.645 71.820 298.110 72.210 ;
        RECT 298.280 72.430 299.970 72.600 ;
        RECT 297.305 71.650 297.475 71.780 ;
        RECT 298.280 71.650 298.450 72.430 ;
        RECT 300.140 72.260 300.310 72.950 ;
        RECT 298.810 72.090 300.310 72.260 ;
        RECT 300.500 72.290 300.710 73.080 ;
        RECT 300.880 72.460 301.230 73.080 ;
        RECT 301.400 72.470 301.570 73.250 ;
        RECT 302.100 73.090 302.270 73.320 ;
        RECT 301.740 72.920 302.270 73.090 ;
        RECT 301.740 72.640 301.960 72.920 ;
        RECT 302.440 72.750 302.680 73.150 ;
        RECT 301.400 72.300 301.805 72.470 ;
        RECT 302.140 72.380 302.680 72.750 ;
        RECT 302.850 72.965 303.170 73.320 ;
        RECT 303.415 73.240 303.720 73.700 ;
        RECT 303.890 72.990 304.140 73.520 ;
        RECT 302.850 72.790 303.175 72.965 ;
        RECT 302.850 72.490 303.765 72.790 ;
        RECT 303.025 72.460 303.765 72.490 ;
        RECT 300.500 72.130 301.175 72.290 ;
        RECT 301.635 72.210 301.805 72.300 ;
        RECT 300.500 72.120 301.465 72.130 ;
        RECT 300.140 71.950 300.310 72.090 ;
        RECT 296.885 71.150 297.135 71.610 ;
        RECT 297.305 71.320 297.555 71.650 ;
        RECT 297.770 71.320 298.450 71.650 ;
        RECT 298.620 71.750 299.695 71.920 ;
        RECT 300.140 71.780 300.700 71.950 ;
        RECT 301.005 71.830 301.465 72.120 ;
        RECT 301.635 72.040 302.855 72.210 ;
        RECT 298.620 71.410 298.790 71.750 ;
        RECT 299.025 71.150 299.355 71.580 ;
        RECT 299.525 71.410 299.695 71.750 ;
        RECT 299.990 71.150 300.360 71.610 ;
        RECT 300.530 71.320 300.700 71.780 ;
        RECT 301.635 71.660 301.805 72.040 ;
        RECT 303.025 71.870 303.195 72.460 ;
        RECT 303.935 72.340 304.140 72.990 ;
        RECT 304.310 72.945 304.560 73.700 ;
        RECT 304.780 72.930 308.290 73.700 ;
        RECT 308.460 72.950 309.670 73.700 ;
        RECT 309.840 72.950 311.050 73.700 ;
        RECT 304.780 72.410 306.430 72.930 ;
        RECT 300.935 71.320 301.805 71.660 ;
        RECT 302.395 71.700 303.195 71.870 ;
        RECT 301.975 71.150 302.225 71.610 ;
        RECT 302.395 71.410 302.565 71.700 ;
        RECT 302.745 71.150 303.075 71.530 ;
        RECT 303.415 71.150 303.720 72.290 ;
        RECT 303.890 71.460 304.140 72.340 ;
        RECT 304.310 71.150 304.560 72.290 ;
        RECT 306.600 72.240 308.290 72.760 ;
        RECT 308.460 72.410 308.980 72.950 ;
        RECT 309.150 72.240 309.670 72.780 ;
        RECT 304.780 71.150 308.290 72.240 ;
        RECT 308.460 71.150 309.670 72.240 ;
        RECT 309.840 72.240 310.360 72.780 ;
        RECT 310.530 72.410 311.050 72.950 ;
        RECT 309.840 71.150 311.050 72.240 ;
        RECT 162.095 70.980 311.135 71.150 ;
        RECT 162.180 69.890 163.390 70.980 ;
        RECT 163.560 69.890 165.230 70.980 ;
        RECT 165.405 70.310 165.660 70.810 ;
        RECT 165.830 70.480 166.160 70.980 ;
        RECT 165.405 70.140 166.155 70.310 ;
        RECT 162.180 69.180 162.700 69.720 ;
        RECT 162.870 69.350 163.390 69.890 ;
        RECT 163.560 69.200 164.310 69.720 ;
        RECT 164.480 69.370 165.230 69.890 ;
        RECT 165.405 69.320 165.755 69.970 ;
        RECT 162.180 68.430 163.390 69.180 ;
        RECT 163.560 68.430 165.230 69.200 ;
        RECT 165.925 69.150 166.155 70.140 ;
        RECT 165.405 68.980 166.155 69.150 ;
        RECT 165.405 68.690 165.660 68.980 ;
        RECT 165.830 68.430 166.160 68.810 ;
        RECT 166.330 68.690 166.500 70.810 ;
        RECT 166.670 70.010 166.995 70.795 ;
        RECT 167.165 70.520 167.415 70.980 ;
        RECT 167.585 70.480 167.835 70.810 ;
        RECT 168.050 70.480 168.730 70.810 ;
        RECT 167.585 70.350 167.755 70.480 ;
        RECT 167.360 70.180 167.755 70.350 ;
        RECT 166.730 68.960 167.190 70.010 ;
        RECT 167.360 68.820 167.530 70.180 ;
        RECT 167.925 69.920 168.390 70.310 ;
        RECT 167.700 69.110 168.050 69.730 ;
        RECT 168.220 69.330 168.390 69.920 ;
        RECT 168.560 69.700 168.730 70.480 ;
        RECT 168.900 70.380 169.070 70.720 ;
        RECT 169.305 70.550 169.635 70.980 ;
        RECT 169.805 70.380 169.975 70.720 ;
        RECT 170.270 70.520 170.640 70.980 ;
        RECT 168.900 70.210 169.975 70.380 ;
        RECT 170.810 70.350 170.980 70.810 ;
        RECT 171.215 70.470 172.085 70.810 ;
        RECT 172.255 70.520 172.505 70.980 ;
        RECT 170.420 70.180 170.980 70.350 ;
        RECT 170.420 70.040 170.590 70.180 ;
        RECT 169.090 69.870 170.590 70.040 ;
        RECT 171.285 70.010 171.745 70.300 ;
        RECT 168.560 69.530 170.250 69.700 ;
        RECT 168.220 69.110 168.575 69.330 ;
        RECT 168.745 68.820 168.915 69.530 ;
        RECT 169.120 69.110 169.910 69.360 ;
        RECT 170.080 69.350 170.250 69.530 ;
        RECT 170.420 69.180 170.590 69.870 ;
        RECT 166.860 68.430 167.190 68.790 ;
        RECT 167.360 68.650 167.855 68.820 ;
        RECT 168.060 68.650 168.915 68.820 ;
        RECT 169.790 68.430 170.120 68.890 ;
        RECT 170.330 68.790 170.590 69.180 ;
        RECT 170.780 70.000 171.745 70.010 ;
        RECT 171.915 70.090 172.085 70.470 ;
        RECT 172.675 70.430 172.845 70.720 ;
        RECT 173.025 70.600 173.355 70.980 ;
        RECT 172.675 70.260 173.475 70.430 ;
        RECT 170.780 69.840 171.455 70.000 ;
        RECT 171.915 69.920 173.135 70.090 ;
        RECT 170.780 69.050 170.990 69.840 ;
        RECT 171.915 69.830 172.085 69.920 ;
        RECT 171.160 69.050 171.510 69.670 ;
        RECT 171.680 69.660 172.085 69.830 ;
        RECT 171.680 68.880 171.850 69.660 ;
        RECT 172.020 69.210 172.240 69.490 ;
        RECT 172.420 69.380 172.960 69.750 ;
        RECT 173.305 69.670 173.475 70.260 ;
        RECT 173.695 69.840 174.000 70.980 ;
        RECT 174.170 69.790 174.420 70.670 ;
        RECT 174.590 69.840 174.840 70.980 ;
        RECT 175.060 69.815 175.350 70.980 ;
        RECT 176.445 69.840 176.780 70.810 ;
        RECT 176.950 69.840 177.120 70.980 ;
        RECT 177.290 70.640 179.320 70.810 ;
        RECT 173.305 69.640 174.045 69.670 ;
        RECT 172.020 69.040 172.550 69.210 ;
        RECT 170.330 68.620 170.680 68.790 ;
        RECT 170.900 68.600 171.850 68.880 ;
        RECT 172.020 68.430 172.210 68.870 ;
        RECT 172.380 68.810 172.550 69.040 ;
        RECT 172.720 68.980 172.960 69.380 ;
        RECT 173.130 69.340 174.045 69.640 ;
        RECT 173.130 69.165 173.455 69.340 ;
        RECT 173.130 68.810 173.450 69.165 ;
        RECT 174.215 69.140 174.420 69.790 ;
        RECT 172.380 68.640 173.450 68.810 ;
        RECT 173.695 68.430 174.000 68.890 ;
        RECT 174.170 68.610 174.420 69.140 ;
        RECT 174.590 68.430 174.840 69.185 ;
        RECT 176.445 69.170 176.615 69.840 ;
        RECT 177.290 69.670 177.460 70.640 ;
        RECT 176.785 69.340 177.040 69.670 ;
        RECT 177.265 69.340 177.460 69.670 ;
        RECT 177.630 70.300 178.755 70.470 ;
        RECT 176.870 69.170 177.040 69.340 ;
        RECT 177.630 69.170 177.800 70.300 ;
        RECT 175.060 68.430 175.350 69.155 ;
        RECT 176.445 68.600 176.700 69.170 ;
        RECT 176.870 69.000 177.800 69.170 ;
        RECT 177.970 69.960 178.980 70.130 ;
        RECT 177.970 69.160 178.140 69.960 ;
        RECT 178.345 69.280 178.620 69.760 ;
        RECT 178.340 69.110 178.620 69.280 ;
        RECT 177.625 68.965 177.800 69.000 ;
        RECT 176.870 68.430 177.200 68.830 ;
        RECT 177.625 68.600 178.155 68.965 ;
        RECT 178.345 68.600 178.620 69.110 ;
        RECT 178.790 68.600 178.980 69.960 ;
        RECT 179.150 69.975 179.320 70.640 ;
        RECT 179.490 70.220 179.660 70.980 ;
        RECT 179.895 70.220 180.410 70.630 ;
        RECT 180.580 70.545 185.925 70.980 ;
        RECT 179.150 69.785 179.900 69.975 ;
        RECT 180.070 69.410 180.410 70.220 ;
        RECT 179.180 69.240 180.410 69.410 ;
        RECT 179.160 68.430 179.670 68.965 ;
        RECT 179.890 68.635 180.135 69.240 ;
        RECT 182.165 68.975 182.505 69.805 ;
        RECT 183.985 69.295 184.335 70.545 ;
        RECT 186.100 69.890 187.770 70.980 ;
        RECT 186.100 69.200 186.850 69.720 ;
        RECT 187.020 69.370 187.770 69.890 ;
        RECT 188.400 69.905 188.670 70.810 ;
        RECT 188.840 70.220 189.170 70.980 ;
        RECT 189.350 70.050 189.520 70.810 ;
        RECT 180.580 68.430 185.925 68.975 ;
        RECT 186.100 68.430 187.770 69.200 ;
        RECT 188.400 69.105 188.570 69.905 ;
        RECT 188.855 69.880 189.520 70.050 ;
        RECT 188.855 69.735 189.025 69.880 ;
        RECT 188.740 69.405 189.025 69.735 ;
        RECT 189.785 69.840 190.120 70.810 ;
        RECT 190.290 69.840 190.460 70.980 ;
        RECT 190.630 70.640 192.660 70.810 ;
        RECT 188.855 69.150 189.025 69.405 ;
        RECT 189.260 69.330 189.590 69.700 ;
        RECT 189.785 69.170 189.955 69.840 ;
        RECT 190.630 69.670 190.800 70.640 ;
        RECT 190.125 69.340 190.380 69.670 ;
        RECT 190.605 69.340 190.800 69.670 ;
        RECT 190.970 70.300 192.095 70.470 ;
        RECT 190.210 69.170 190.380 69.340 ;
        RECT 190.970 69.170 191.140 70.300 ;
        RECT 188.400 68.600 188.660 69.105 ;
        RECT 188.855 68.980 189.520 69.150 ;
        RECT 188.840 68.430 189.170 68.810 ;
        RECT 189.350 68.600 189.520 68.980 ;
        RECT 189.785 68.600 190.040 69.170 ;
        RECT 190.210 69.000 191.140 69.170 ;
        RECT 191.310 69.960 192.320 70.130 ;
        RECT 191.310 69.160 191.480 69.960 ;
        RECT 190.965 68.965 191.140 69.000 ;
        RECT 190.210 68.430 190.540 68.830 ;
        RECT 190.965 68.600 191.495 68.965 ;
        RECT 191.685 68.940 191.960 69.760 ;
        RECT 191.680 68.770 191.960 68.940 ;
        RECT 191.685 68.600 191.960 68.770 ;
        RECT 192.130 68.600 192.320 69.960 ;
        RECT 192.490 69.975 192.660 70.640 ;
        RECT 192.830 70.220 193.000 70.980 ;
        RECT 193.235 70.220 193.750 70.630 ;
        RECT 192.490 69.785 193.240 69.975 ;
        RECT 193.410 69.410 193.750 70.220 ;
        RECT 193.925 69.830 194.185 70.980 ;
        RECT 194.360 69.905 194.615 70.810 ;
        RECT 194.785 70.220 195.115 70.980 ;
        RECT 195.330 70.050 195.500 70.810 ;
        RECT 192.520 69.240 193.750 69.410 ;
        RECT 192.500 68.430 193.010 68.965 ;
        RECT 193.230 68.635 193.475 69.240 ;
        RECT 193.925 68.430 194.185 69.270 ;
        RECT 194.360 69.175 194.530 69.905 ;
        RECT 194.785 69.880 195.500 70.050 ;
        RECT 196.220 70.220 196.735 70.630 ;
        RECT 196.970 70.220 197.140 70.980 ;
        RECT 197.310 70.640 199.340 70.810 ;
        RECT 194.785 69.670 194.955 69.880 ;
        RECT 194.700 69.340 194.955 69.670 ;
        RECT 194.360 68.600 194.615 69.175 ;
        RECT 194.785 69.150 194.955 69.340 ;
        RECT 195.235 69.330 195.590 69.700 ;
        RECT 196.220 69.410 196.560 70.220 ;
        RECT 197.310 69.975 197.480 70.640 ;
        RECT 197.875 70.300 199.000 70.470 ;
        RECT 196.730 69.785 197.480 69.975 ;
        RECT 197.650 69.960 198.660 70.130 ;
        RECT 196.220 69.240 197.450 69.410 ;
        RECT 194.785 68.980 195.500 69.150 ;
        RECT 194.785 68.430 195.115 68.810 ;
        RECT 195.330 68.600 195.500 68.980 ;
        RECT 196.495 68.635 196.740 69.240 ;
        RECT 196.960 68.430 197.470 68.965 ;
        RECT 197.650 68.600 197.840 69.960 ;
        RECT 198.010 68.940 198.285 69.760 ;
        RECT 198.490 69.160 198.660 69.960 ;
        RECT 198.830 69.170 199.000 70.300 ;
        RECT 199.170 69.670 199.340 70.640 ;
        RECT 199.510 69.840 199.680 70.980 ;
        RECT 199.850 69.840 200.185 70.810 ;
        RECT 199.170 69.340 199.365 69.670 ;
        RECT 199.590 69.340 199.845 69.670 ;
        RECT 199.590 69.170 199.760 69.340 ;
        RECT 200.015 69.170 200.185 69.840 ;
        RECT 200.820 69.815 201.110 70.980 ;
        RECT 201.280 69.890 202.950 70.980 ;
        RECT 203.130 69.915 203.440 70.980 ;
        RECT 203.610 70.310 203.845 70.810 ;
        RECT 204.015 70.520 204.345 70.980 ;
        RECT 204.540 70.640 205.650 70.810 ;
        RECT 204.540 70.480 204.730 70.640 ;
        RECT 204.960 70.310 205.260 70.470 ;
        RECT 203.610 70.130 205.260 70.310 ;
        RECT 205.430 70.130 205.650 70.640 ;
        RECT 205.820 70.130 206.150 70.980 ;
        RECT 198.830 69.000 199.760 69.170 ;
        RECT 198.830 68.965 199.005 69.000 ;
        RECT 198.010 68.770 198.290 68.940 ;
        RECT 198.010 68.600 198.285 68.770 ;
        RECT 198.475 68.600 199.005 68.965 ;
        RECT 199.430 68.430 199.760 68.830 ;
        RECT 199.930 68.600 200.185 69.170 ;
        RECT 201.280 69.200 202.030 69.720 ;
        RECT 202.200 69.370 202.950 69.890 ;
        RECT 200.820 68.430 201.110 69.155 ;
        RECT 201.280 68.430 202.950 69.200 ;
        RECT 203.125 69.110 203.440 69.745 ;
        RECT 203.610 68.940 203.820 70.130 ;
        RECT 204.160 69.790 206.135 69.960 ;
        RECT 206.350 69.915 206.660 70.980 ;
        RECT 206.830 70.310 207.065 70.810 ;
        RECT 207.235 70.520 207.565 70.980 ;
        RECT 207.760 70.640 208.870 70.810 ;
        RECT 207.760 70.480 207.950 70.640 ;
        RECT 208.180 70.310 208.480 70.470 ;
        RECT 206.830 70.130 208.480 70.310 ;
        RECT 208.650 70.130 208.870 70.640 ;
        RECT 209.040 70.130 209.370 70.980 ;
        RECT 204.160 69.620 204.655 69.790 ;
        RECT 204.100 69.450 204.655 69.620 ;
        RECT 204.160 69.420 204.655 69.450 ;
        RECT 204.835 69.420 205.635 69.620 ;
        RECT 205.805 69.400 206.135 69.790 ;
        RECT 203.990 69.060 206.150 69.230 ;
        RECT 206.345 69.110 206.660 69.745 ;
        RECT 203.130 68.770 203.440 68.940 ;
        RECT 203.990 68.770 204.320 69.060 ;
        RECT 203.130 68.600 204.320 68.770 ;
        RECT 204.560 68.430 204.730 68.890 ;
        RECT 204.960 68.600 205.290 69.060 ;
        RECT 205.470 68.430 205.640 68.890 ;
        RECT 205.820 68.600 206.150 69.060 ;
        RECT 206.830 68.940 207.040 70.130 ;
        RECT 209.560 70.010 209.870 70.810 ;
        RECT 210.040 70.180 210.350 70.980 ;
        RECT 210.520 70.350 210.780 70.810 ;
        RECT 210.950 70.520 211.205 70.980 ;
        RECT 211.380 70.350 211.640 70.810 ;
        RECT 210.520 70.180 211.640 70.350 ;
        RECT 207.380 69.790 209.355 69.960 ;
        RECT 207.380 69.620 207.875 69.790 ;
        RECT 207.320 69.450 207.875 69.620 ;
        RECT 207.380 69.420 207.875 69.450 ;
        RECT 208.055 69.420 208.855 69.620 ;
        RECT 209.025 69.400 209.355 69.790 ;
        RECT 209.560 69.840 210.590 70.010 ;
        RECT 207.210 69.060 209.370 69.230 ;
        RECT 206.350 68.770 206.660 68.940 ;
        RECT 207.210 68.770 207.540 69.060 ;
        RECT 206.350 68.600 207.540 68.770 ;
        RECT 207.780 68.430 207.950 68.890 ;
        RECT 208.180 68.600 208.510 69.060 ;
        RECT 208.690 68.430 208.860 68.890 ;
        RECT 209.040 68.600 209.370 69.060 ;
        RECT 209.560 68.930 209.730 69.840 ;
        RECT 209.900 69.100 210.250 69.670 ;
        RECT 210.420 69.590 210.590 69.840 ;
        RECT 211.380 69.930 211.640 70.180 ;
        RECT 211.810 70.110 212.095 70.980 ;
        RECT 212.320 70.010 212.590 70.780 ;
        RECT 212.760 70.200 213.090 70.980 ;
        RECT 213.295 70.375 213.480 70.780 ;
        RECT 213.650 70.555 213.985 70.980 ;
        RECT 214.160 70.545 219.505 70.980 ;
        RECT 219.680 70.545 225.025 70.980 ;
        RECT 213.295 70.200 213.960 70.375 ;
        RECT 211.380 69.760 212.135 69.930 ;
        RECT 210.420 69.420 211.560 69.590 ;
        RECT 211.730 69.250 212.135 69.760 ;
        RECT 210.485 69.080 212.135 69.250 ;
        RECT 212.320 69.840 213.450 70.010 ;
        RECT 209.560 68.600 209.860 68.930 ;
        RECT 210.030 68.430 210.305 68.910 ;
        RECT 210.485 68.690 210.780 69.080 ;
        RECT 210.950 68.430 211.205 68.910 ;
        RECT 211.380 68.690 211.640 69.080 ;
        RECT 212.320 68.930 212.490 69.840 ;
        RECT 212.660 69.090 213.020 69.670 ;
        RECT 213.200 69.340 213.450 69.840 ;
        RECT 213.620 69.170 213.960 70.200 ;
        RECT 213.275 69.000 213.960 69.170 ;
        RECT 211.810 68.430 212.090 68.910 ;
        RECT 212.320 68.600 212.580 68.930 ;
        RECT 212.790 68.430 213.065 68.910 ;
        RECT 213.275 68.600 213.480 69.000 ;
        RECT 215.745 68.975 216.085 69.805 ;
        RECT 217.565 69.295 217.915 70.545 ;
        RECT 221.265 68.975 221.605 69.805 ;
        RECT 223.085 69.295 223.435 70.545 ;
        RECT 225.200 69.890 226.410 70.980 ;
        RECT 225.200 69.180 225.720 69.720 ;
        RECT 225.890 69.350 226.410 69.890 ;
        RECT 226.580 69.815 226.870 70.980 ;
        RECT 227.130 69.970 227.300 70.810 ;
        RECT 227.470 70.640 228.640 70.810 ;
        RECT 227.470 70.140 227.800 70.640 ;
        RECT 228.310 70.600 228.640 70.640 ;
        RECT 228.830 70.560 229.185 70.980 ;
        RECT 227.970 70.380 228.200 70.470 ;
        RECT 229.355 70.380 229.605 70.810 ;
        RECT 227.970 70.140 229.605 70.380 ;
        RECT 229.775 70.220 230.105 70.980 ;
        RECT 230.275 70.140 230.530 70.810 ;
        RECT 227.130 69.800 230.190 69.970 ;
        RECT 227.045 69.420 227.395 69.630 ;
        RECT 227.565 69.420 228.010 69.620 ;
        RECT 228.180 69.420 228.655 69.620 ;
        RECT 213.650 68.430 213.985 68.830 ;
        RECT 214.160 68.430 219.505 68.975 ;
        RECT 219.680 68.430 225.025 68.975 ;
        RECT 225.200 68.430 226.410 69.180 ;
        RECT 226.580 68.430 226.870 69.155 ;
        RECT 227.130 69.080 228.195 69.250 ;
        RECT 227.130 68.600 227.300 69.080 ;
        RECT 227.470 68.430 227.800 68.910 ;
        RECT 228.025 68.850 228.195 69.080 ;
        RECT 228.375 69.020 228.655 69.420 ;
        RECT 228.925 69.420 229.255 69.620 ;
        RECT 229.425 69.450 229.800 69.620 ;
        RECT 229.425 69.420 229.790 69.450 ;
        RECT 228.925 69.020 229.210 69.420 ;
        RECT 230.020 69.250 230.190 69.800 ;
        RECT 229.390 69.080 230.190 69.250 ;
        RECT 229.390 68.850 229.560 69.080 ;
        RECT 230.360 69.010 230.530 70.140 ;
        RECT 230.720 69.890 231.930 70.980 ;
        RECT 230.345 68.940 230.530 69.010 ;
        RECT 230.320 68.930 230.530 68.940 ;
        RECT 228.025 68.600 229.560 68.850 ;
        RECT 229.730 68.430 230.060 68.910 ;
        RECT 230.275 68.600 230.530 68.930 ;
        RECT 230.720 69.180 231.240 69.720 ;
        RECT 231.410 69.350 231.930 69.890 ;
        RECT 230.720 68.430 231.930 69.180 ;
        RECT 232.100 68.600 232.850 70.810 ;
        RECT 234.025 70.360 234.200 70.810 ;
        RECT 234.370 70.540 234.700 70.980 ;
        RECT 235.005 70.390 235.175 70.810 ;
        RECT 235.410 70.570 236.080 70.980 ;
        RECT 236.295 70.390 236.465 70.810 ;
        RECT 236.665 70.570 236.995 70.980 ;
        RECT 234.025 70.190 234.655 70.360 ;
        RECT 233.940 69.340 234.305 70.020 ;
        RECT 234.485 69.670 234.655 70.190 ;
        RECT 235.005 70.220 237.020 70.390 ;
        RECT 234.485 69.340 234.835 69.670 ;
        RECT 234.485 69.170 234.655 69.340 ;
        RECT 234.025 69.000 234.655 69.170 ;
        RECT 234.025 68.600 234.200 69.000 ;
        RECT 235.005 68.930 235.175 70.220 ;
        RECT 234.370 68.430 234.700 68.810 ;
        RECT 234.945 68.600 235.175 68.930 ;
        RECT 235.375 68.765 235.655 70.040 ;
        RECT 235.880 69.960 236.150 70.040 ;
        RECT 235.840 69.790 236.150 69.960 ;
        RECT 235.880 68.765 236.150 69.790 ;
        RECT 236.340 69.010 236.680 70.040 ;
        RECT 236.850 69.670 237.020 70.220 ;
        RECT 237.190 69.840 237.450 70.810 ;
        RECT 237.620 70.545 242.965 70.980 ;
        RECT 243.145 70.600 243.480 70.980 ;
        RECT 236.850 69.340 237.110 69.670 ;
        RECT 237.280 69.150 237.450 69.840 ;
        RECT 236.610 68.430 236.940 68.810 ;
        RECT 237.110 68.685 237.450 69.150 ;
        RECT 239.205 68.975 239.545 69.805 ;
        RECT 241.025 69.295 241.375 70.545 ;
        RECT 243.140 69.110 243.380 70.420 ;
        RECT 243.650 70.010 243.900 70.810 ;
        RECT 244.120 70.260 244.450 70.980 ;
        RECT 244.635 70.010 244.885 70.810 ;
        RECT 245.350 70.180 245.680 70.980 ;
        RECT 245.850 70.550 246.190 70.810 ;
        RECT 243.550 69.840 245.740 70.010 ;
        RECT 237.110 68.640 237.445 68.685 ;
        RECT 237.620 68.430 242.965 68.975 ;
        RECT 243.550 68.930 243.720 69.840 ;
        RECT 245.425 69.670 245.740 69.840 ;
        RECT 243.225 68.600 243.720 68.930 ;
        RECT 243.940 68.705 244.290 69.670 ;
        RECT 244.470 68.700 244.770 69.670 ;
        RECT 244.950 68.700 245.230 69.670 ;
        RECT 245.425 69.420 245.755 69.670 ;
        RECT 245.410 68.430 245.680 69.230 ;
        RECT 245.930 69.150 246.190 70.550 ;
        RECT 246.360 70.545 251.705 70.980 ;
        RECT 245.850 68.640 246.190 69.150 ;
        RECT 247.945 68.975 248.285 69.805 ;
        RECT 249.765 69.295 250.115 70.545 ;
        RECT 252.340 69.815 252.630 70.980 ;
        RECT 252.890 69.970 253.060 70.810 ;
        RECT 253.230 70.640 254.400 70.810 ;
        RECT 253.230 70.140 253.560 70.640 ;
        RECT 254.070 70.600 254.400 70.640 ;
        RECT 254.590 70.560 254.945 70.980 ;
        RECT 253.730 70.380 253.960 70.470 ;
        RECT 255.115 70.380 255.365 70.810 ;
        RECT 253.730 70.140 255.365 70.380 ;
        RECT 255.535 70.220 255.865 70.980 ;
        RECT 256.035 70.140 256.290 70.810 ;
        RECT 257.600 70.310 257.880 70.980 ;
        RECT 252.890 69.800 255.950 69.970 ;
        RECT 252.805 69.420 253.155 69.630 ;
        RECT 253.325 69.420 253.770 69.620 ;
        RECT 253.940 69.420 254.415 69.620 ;
        RECT 246.360 68.430 251.705 68.975 ;
        RECT 252.340 68.430 252.630 69.155 ;
        RECT 252.890 69.080 253.955 69.250 ;
        RECT 252.890 68.600 253.060 69.080 ;
        RECT 253.230 68.430 253.560 68.910 ;
        RECT 253.785 68.850 253.955 69.080 ;
        RECT 254.135 69.020 254.415 69.420 ;
        RECT 254.685 69.420 255.015 69.620 ;
        RECT 255.185 69.420 255.550 69.620 ;
        RECT 254.685 69.020 254.970 69.420 ;
        RECT 255.780 69.250 255.950 69.800 ;
        RECT 255.150 69.080 255.950 69.250 ;
        RECT 255.150 68.850 255.320 69.080 ;
        RECT 256.120 69.010 256.290 70.140 ;
        RECT 258.050 70.090 258.350 70.640 ;
        RECT 258.550 70.260 258.880 70.980 ;
        RECT 259.070 70.260 259.530 70.810 ;
        RECT 259.700 70.545 265.045 70.980 ;
        RECT 265.220 70.545 270.565 70.980 ;
        RECT 257.415 69.670 257.680 70.030 ;
        RECT 258.050 69.920 258.990 70.090 ;
        RECT 258.820 69.670 258.990 69.920 ;
        RECT 257.415 69.420 258.090 69.670 ;
        RECT 258.310 69.420 258.650 69.670 ;
        RECT 258.820 69.340 259.110 69.670 ;
        RECT 258.820 69.250 258.990 69.340 ;
        RECT 256.105 68.940 256.290 69.010 ;
        RECT 256.080 68.930 256.290 68.940 ;
        RECT 253.785 68.600 255.320 68.850 ;
        RECT 255.490 68.430 255.820 68.910 ;
        RECT 256.035 68.600 256.290 68.930 ;
        RECT 257.600 69.060 258.990 69.250 ;
        RECT 257.600 68.700 257.930 69.060 ;
        RECT 259.280 68.890 259.530 70.260 ;
        RECT 261.285 68.975 261.625 69.805 ;
        RECT 263.105 69.295 263.455 70.545 ;
        RECT 266.805 68.975 267.145 69.805 ;
        RECT 268.625 69.295 268.975 70.545 ;
        RECT 270.740 69.890 272.410 70.980 ;
        RECT 270.740 69.200 271.490 69.720 ;
        RECT 271.660 69.370 272.410 69.890 ;
        RECT 272.585 69.840 272.920 70.810 ;
        RECT 273.090 69.840 273.260 70.980 ;
        RECT 273.430 70.640 275.460 70.810 ;
        RECT 258.550 68.430 258.800 68.890 ;
        RECT 258.970 68.600 259.530 68.890 ;
        RECT 259.700 68.430 265.045 68.975 ;
        RECT 265.220 68.430 270.565 68.975 ;
        RECT 270.740 68.430 272.410 69.200 ;
        RECT 272.585 69.170 272.755 69.840 ;
        RECT 273.430 69.670 273.600 70.640 ;
        RECT 272.925 69.340 273.180 69.670 ;
        RECT 273.405 69.340 273.600 69.670 ;
        RECT 273.770 70.300 274.895 70.470 ;
        RECT 273.010 69.170 273.180 69.340 ;
        RECT 273.770 69.170 273.940 70.300 ;
        RECT 272.585 68.600 272.840 69.170 ;
        RECT 273.010 69.000 273.940 69.170 ;
        RECT 274.110 69.960 275.120 70.130 ;
        RECT 274.110 69.160 274.280 69.960 ;
        RECT 274.485 69.280 274.760 69.760 ;
        RECT 274.480 69.110 274.760 69.280 ;
        RECT 273.765 68.965 273.940 69.000 ;
        RECT 273.010 68.430 273.340 68.830 ;
        RECT 273.765 68.600 274.295 68.965 ;
        RECT 274.485 68.600 274.760 69.110 ;
        RECT 274.930 68.600 275.120 69.960 ;
        RECT 275.290 69.975 275.460 70.640 ;
        RECT 275.630 70.220 275.800 70.980 ;
        RECT 276.035 70.220 276.550 70.630 ;
        RECT 275.290 69.785 276.040 69.975 ;
        RECT 276.210 69.410 276.550 70.220 ;
        RECT 276.720 69.890 277.930 70.980 ;
        RECT 275.320 69.240 276.550 69.410 ;
        RECT 275.300 68.430 275.810 68.965 ;
        RECT 276.030 68.635 276.275 69.240 ;
        RECT 276.720 69.180 277.240 69.720 ;
        RECT 277.410 69.350 277.930 69.890 ;
        RECT 278.100 69.815 278.390 70.980 ;
        RECT 278.570 70.260 278.900 70.980 ;
        RECT 278.560 69.620 278.790 69.960 ;
        RECT 279.080 69.620 279.295 70.735 ;
        RECT 279.490 70.035 279.820 70.810 ;
        RECT 279.990 70.205 280.700 70.980 ;
        RECT 279.490 69.820 280.640 70.035 ;
        RECT 278.560 69.420 278.890 69.620 ;
        RECT 279.080 69.440 279.530 69.620 ;
        RECT 279.200 69.420 279.530 69.440 ;
        RECT 279.700 69.420 280.170 69.650 ;
        RECT 280.355 69.250 280.640 69.820 ;
        RECT 280.870 69.375 281.150 70.810 ;
        RECT 276.720 68.430 277.930 69.180 ;
        RECT 278.100 68.430 278.390 69.155 ;
        RECT 278.560 69.060 279.740 69.250 ;
        RECT 278.560 68.600 278.900 69.060 ;
        RECT 279.410 68.980 279.740 69.060 ;
        RECT 279.930 69.060 280.640 69.250 ;
        RECT 279.930 68.920 280.230 69.060 ;
        RECT 279.915 68.910 280.230 68.920 ;
        RECT 279.905 68.900 280.230 68.910 ;
        RECT 279.895 68.895 280.230 68.900 ;
        RECT 279.070 68.430 279.240 68.890 ;
        RECT 279.890 68.885 280.230 68.895 ;
        RECT 279.885 68.880 280.230 68.885 ;
        RECT 279.880 68.870 280.230 68.880 ;
        RECT 279.875 68.865 280.230 68.870 ;
        RECT 279.870 68.600 280.230 68.865 ;
        RECT 280.470 68.430 280.640 68.890 ;
        RECT 280.810 68.600 281.150 69.375 ;
        RECT 281.320 69.905 281.590 70.810 ;
        RECT 281.760 70.220 282.090 70.980 ;
        RECT 282.270 70.050 282.440 70.810 ;
        RECT 281.320 69.105 281.490 69.905 ;
        RECT 281.775 69.880 282.440 70.050 ;
        RECT 281.775 69.735 281.945 69.880 ;
        RECT 281.660 69.405 281.945 69.735 ;
        RECT 282.705 69.840 283.040 70.810 ;
        RECT 283.210 69.840 283.380 70.980 ;
        RECT 283.550 70.640 285.580 70.810 ;
        RECT 281.775 69.150 281.945 69.405 ;
        RECT 282.180 69.330 282.510 69.700 ;
        RECT 282.705 69.170 282.875 69.840 ;
        RECT 283.550 69.670 283.720 70.640 ;
        RECT 283.045 69.340 283.300 69.670 ;
        RECT 283.525 69.340 283.720 69.670 ;
        RECT 283.890 70.300 285.015 70.470 ;
        RECT 283.130 69.170 283.300 69.340 ;
        RECT 283.890 69.170 284.060 70.300 ;
        RECT 281.320 68.600 281.580 69.105 ;
        RECT 281.775 68.980 282.440 69.150 ;
        RECT 281.760 68.430 282.090 68.810 ;
        RECT 282.270 68.600 282.440 68.980 ;
        RECT 282.705 68.600 282.960 69.170 ;
        RECT 283.130 69.000 284.060 69.170 ;
        RECT 284.230 69.960 285.240 70.130 ;
        RECT 284.230 69.160 284.400 69.960 ;
        RECT 284.605 69.620 284.880 69.760 ;
        RECT 284.600 69.450 284.880 69.620 ;
        RECT 283.885 68.965 284.060 69.000 ;
        RECT 283.130 68.430 283.460 68.830 ;
        RECT 283.885 68.600 284.415 68.965 ;
        RECT 284.605 68.600 284.880 69.450 ;
        RECT 285.050 68.600 285.240 69.960 ;
        RECT 285.410 69.975 285.580 70.640 ;
        RECT 285.750 70.220 285.920 70.980 ;
        RECT 286.155 70.220 286.670 70.630 ;
        RECT 285.410 69.785 286.160 69.975 ;
        RECT 286.330 69.410 286.670 70.220 ;
        RECT 285.440 69.240 286.670 69.410 ;
        RECT 286.845 69.840 287.180 70.810 ;
        RECT 287.350 69.840 287.520 70.980 ;
        RECT 287.690 70.640 289.720 70.810 ;
        RECT 285.420 68.430 285.930 68.965 ;
        RECT 286.150 68.635 286.395 69.240 ;
        RECT 286.845 69.170 287.015 69.840 ;
        RECT 287.690 69.670 287.860 70.640 ;
        RECT 287.185 69.340 287.440 69.670 ;
        RECT 287.665 69.340 287.860 69.670 ;
        RECT 288.030 70.300 289.155 70.470 ;
        RECT 287.270 69.170 287.440 69.340 ;
        RECT 288.030 69.170 288.200 70.300 ;
        RECT 286.845 68.600 287.100 69.170 ;
        RECT 287.270 69.000 288.200 69.170 ;
        RECT 288.370 69.960 289.380 70.130 ;
        RECT 288.370 69.160 288.540 69.960 ;
        RECT 288.745 69.620 289.020 69.760 ;
        RECT 288.740 69.450 289.020 69.620 ;
        RECT 288.025 68.965 288.200 69.000 ;
        RECT 287.270 68.430 287.600 68.830 ;
        RECT 288.025 68.600 288.555 68.965 ;
        RECT 288.745 68.600 289.020 69.450 ;
        RECT 289.190 68.600 289.380 69.960 ;
        RECT 289.550 69.975 289.720 70.640 ;
        RECT 289.890 70.220 290.060 70.980 ;
        RECT 290.295 70.220 290.810 70.630 ;
        RECT 289.550 69.785 290.300 69.975 ;
        RECT 290.470 69.410 290.810 70.220 ;
        RECT 290.980 69.890 293.570 70.980 ;
        RECT 294.205 70.310 294.460 70.810 ;
        RECT 294.630 70.480 294.960 70.980 ;
        RECT 294.205 70.140 294.955 70.310 ;
        RECT 289.580 69.240 290.810 69.410 ;
        RECT 289.560 68.430 290.070 68.965 ;
        RECT 290.290 68.635 290.535 69.240 ;
        RECT 290.980 69.200 292.190 69.720 ;
        RECT 292.360 69.370 293.570 69.890 ;
        RECT 294.205 69.320 294.555 69.970 ;
        RECT 290.980 68.430 293.570 69.200 ;
        RECT 294.725 69.150 294.955 70.140 ;
        RECT 294.205 68.980 294.955 69.150 ;
        RECT 294.205 68.690 294.460 68.980 ;
        RECT 294.630 68.430 294.960 68.810 ;
        RECT 295.130 68.690 295.300 70.810 ;
        RECT 295.470 70.010 295.795 70.795 ;
        RECT 295.965 70.520 296.215 70.980 ;
        RECT 296.385 70.480 296.635 70.810 ;
        RECT 296.850 70.480 297.530 70.810 ;
        RECT 296.385 70.350 296.555 70.480 ;
        RECT 296.160 70.180 296.555 70.350 ;
        RECT 295.530 68.960 295.990 70.010 ;
        RECT 296.160 68.820 296.330 70.180 ;
        RECT 296.725 69.920 297.190 70.310 ;
        RECT 296.500 69.110 296.850 69.730 ;
        RECT 297.020 69.330 297.190 69.920 ;
        RECT 297.360 69.700 297.530 70.480 ;
        RECT 297.700 70.380 297.870 70.720 ;
        RECT 298.105 70.550 298.435 70.980 ;
        RECT 298.605 70.380 298.775 70.720 ;
        RECT 299.070 70.520 299.440 70.980 ;
        RECT 297.700 70.210 298.775 70.380 ;
        RECT 299.610 70.350 299.780 70.810 ;
        RECT 300.015 70.470 300.885 70.810 ;
        RECT 301.055 70.520 301.305 70.980 ;
        RECT 299.220 70.180 299.780 70.350 ;
        RECT 299.220 70.040 299.390 70.180 ;
        RECT 297.890 69.870 299.390 70.040 ;
        RECT 300.085 70.010 300.545 70.300 ;
        RECT 297.360 69.530 299.050 69.700 ;
        RECT 297.020 69.110 297.375 69.330 ;
        RECT 297.545 68.820 297.715 69.530 ;
        RECT 297.920 69.110 298.710 69.360 ;
        RECT 298.880 69.350 299.050 69.530 ;
        RECT 299.220 69.180 299.390 69.870 ;
        RECT 295.660 68.430 295.990 68.790 ;
        RECT 296.160 68.650 296.655 68.820 ;
        RECT 296.860 68.650 297.715 68.820 ;
        RECT 298.590 68.430 298.920 68.890 ;
        RECT 299.130 68.790 299.390 69.180 ;
        RECT 299.580 70.000 300.545 70.010 ;
        RECT 300.715 70.090 300.885 70.470 ;
        RECT 301.475 70.430 301.645 70.720 ;
        RECT 301.825 70.600 302.155 70.980 ;
        RECT 301.475 70.260 302.275 70.430 ;
        RECT 299.580 69.840 300.255 70.000 ;
        RECT 300.715 69.920 301.935 70.090 ;
        RECT 299.580 69.050 299.790 69.840 ;
        RECT 300.715 69.830 300.885 69.920 ;
        RECT 299.960 69.050 300.310 69.670 ;
        RECT 300.480 69.660 300.885 69.830 ;
        RECT 300.480 68.880 300.650 69.660 ;
        RECT 300.820 69.210 301.040 69.490 ;
        RECT 301.220 69.380 301.760 69.750 ;
        RECT 302.105 69.670 302.275 70.260 ;
        RECT 302.495 69.840 302.800 70.980 ;
        RECT 302.970 69.790 303.220 70.670 ;
        RECT 303.390 69.840 303.640 70.980 ;
        RECT 303.860 69.815 304.150 70.980 ;
        RECT 304.410 70.050 304.580 70.810 ;
        RECT 304.795 70.220 305.125 70.980 ;
        RECT 304.410 69.880 305.125 70.050 ;
        RECT 305.295 69.905 305.550 70.810 ;
        RECT 302.105 69.640 302.845 69.670 ;
        RECT 300.820 69.040 301.350 69.210 ;
        RECT 299.130 68.620 299.480 68.790 ;
        RECT 299.700 68.600 300.650 68.880 ;
        RECT 300.820 68.430 301.010 68.870 ;
        RECT 301.180 68.810 301.350 69.040 ;
        RECT 301.520 68.980 301.760 69.380 ;
        RECT 301.930 69.340 302.845 69.640 ;
        RECT 301.930 69.165 302.255 69.340 ;
        RECT 301.930 68.810 302.250 69.165 ;
        RECT 303.015 69.140 303.220 69.790 ;
        RECT 304.320 69.330 304.675 69.700 ;
        RECT 304.955 69.670 305.125 69.880 ;
        RECT 304.955 69.340 305.210 69.670 ;
        RECT 301.180 68.640 302.250 68.810 ;
        RECT 302.495 68.430 302.800 68.890 ;
        RECT 302.970 68.610 303.220 69.140 ;
        RECT 303.390 68.430 303.640 69.185 ;
        RECT 303.860 68.430 304.150 69.155 ;
        RECT 304.955 69.150 305.125 69.340 ;
        RECT 305.380 69.175 305.550 69.905 ;
        RECT 305.725 69.830 305.985 70.980 ;
        RECT 306.160 69.890 307.830 70.980 ;
        RECT 304.410 68.980 305.125 69.150 ;
        RECT 304.410 68.600 304.580 68.980 ;
        RECT 304.795 68.430 305.125 68.810 ;
        RECT 305.295 68.600 305.550 69.175 ;
        RECT 305.725 68.430 305.985 69.270 ;
        RECT 306.160 69.200 306.910 69.720 ;
        RECT 307.080 69.370 307.830 69.890 ;
        RECT 308.460 69.905 308.730 70.810 ;
        RECT 308.900 70.220 309.230 70.980 ;
        RECT 309.410 70.050 309.580 70.810 ;
        RECT 306.160 68.430 307.830 69.200 ;
        RECT 308.460 69.105 308.630 69.905 ;
        RECT 308.915 69.880 309.580 70.050 ;
        RECT 309.840 69.890 311.050 70.980 ;
        RECT 308.915 69.735 309.085 69.880 ;
        RECT 308.800 69.405 309.085 69.735 ;
        RECT 308.915 69.150 309.085 69.405 ;
        RECT 309.320 69.330 309.650 69.700 ;
        RECT 309.840 69.350 310.360 69.890 ;
        RECT 310.530 69.180 311.050 69.720 ;
        RECT 308.460 68.600 308.720 69.105 ;
        RECT 308.915 68.980 309.580 69.150 ;
        RECT 308.900 68.430 309.230 68.810 ;
        RECT 309.410 68.600 309.580 68.980 ;
        RECT 309.840 68.430 311.050 69.180 ;
        RECT 162.095 68.260 311.135 68.430 ;
        RECT 162.180 67.510 163.390 68.260 ;
        RECT 163.560 67.715 168.905 68.260 ;
        RECT 162.180 66.970 162.700 67.510 ;
        RECT 162.870 66.800 163.390 67.340 ;
        RECT 165.145 66.885 165.485 67.715 ;
        RECT 169.080 67.585 169.340 68.090 ;
        RECT 169.520 67.880 169.850 68.260 ;
        RECT 170.030 67.710 170.200 68.090 ;
        RECT 162.180 65.710 163.390 66.800 ;
        RECT 166.965 66.145 167.315 67.395 ;
        RECT 169.080 66.785 169.250 67.585 ;
        RECT 169.535 67.540 170.200 67.710 ;
        RECT 170.550 67.710 170.720 68.090 ;
        RECT 170.900 67.880 171.230 68.260 ;
        RECT 170.550 67.540 171.215 67.710 ;
        RECT 171.410 67.585 171.670 68.090 ;
        RECT 169.535 67.285 169.705 67.540 ;
        RECT 169.420 66.955 169.705 67.285 ;
        RECT 169.940 66.990 170.270 67.360 ;
        RECT 170.480 66.990 170.810 67.360 ;
        RECT 171.045 67.285 171.215 67.540 ;
        RECT 169.535 66.810 169.705 66.955 ;
        RECT 171.045 66.955 171.330 67.285 ;
        RECT 171.045 66.810 171.215 66.955 ;
        RECT 163.560 65.710 168.905 66.145 ;
        RECT 169.080 65.880 169.350 66.785 ;
        RECT 169.535 66.640 170.200 66.810 ;
        RECT 169.520 65.710 169.850 66.470 ;
        RECT 170.030 65.880 170.200 66.640 ;
        RECT 170.550 66.640 171.215 66.810 ;
        RECT 171.500 66.785 171.670 67.585 ;
        RECT 171.845 67.710 172.100 68.000 ;
        RECT 172.270 67.880 172.600 68.260 ;
        RECT 171.845 67.540 172.595 67.710 ;
        RECT 170.550 65.880 170.720 66.640 ;
        RECT 170.900 65.710 171.230 66.470 ;
        RECT 171.400 65.880 171.670 66.785 ;
        RECT 171.845 66.720 172.195 67.370 ;
        RECT 172.365 66.550 172.595 67.540 ;
        RECT 171.845 66.380 172.595 66.550 ;
        RECT 171.845 65.880 172.100 66.380 ;
        RECT 172.270 65.710 172.600 66.210 ;
        RECT 172.770 65.880 172.940 68.000 ;
        RECT 173.300 67.900 173.630 68.260 ;
        RECT 173.800 67.870 174.295 68.040 ;
        RECT 174.500 67.870 175.355 68.040 ;
        RECT 173.170 66.680 173.630 67.730 ;
        RECT 173.110 65.895 173.435 66.680 ;
        RECT 173.800 66.510 173.970 67.870 ;
        RECT 174.140 66.960 174.490 67.580 ;
        RECT 174.660 67.360 175.015 67.580 ;
        RECT 174.660 66.770 174.830 67.360 ;
        RECT 175.185 67.160 175.355 67.870 ;
        RECT 176.230 67.800 176.560 68.260 ;
        RECT 176.770 67.900 177.120 68.070 ;
        RECT 175.560 67.330 176.350 67.580 ;
        RECT 176.770 67.510 177.030 67.900 ;
        RECT 177.340 67.810 178.290 68.090 ;
        RECT 178.460 67.820 178.650 68.260 ;
        RECT 178.820 67.880 179.890 68.050 ;
        RECT 176.520 67.160 176.690 67.340 ;
        RECT 173.800 66.340 174.195 66.510 ;
        RECT 174.365 66.380 174.830 66.770 ;
        RECT 175.000 66.990 176.690 67.160 ;
        RECT 174.025 66.210 174.195 66.340 ;
        RECT 175.000 66.210 175.170 66.990 ;
        RECT 176.860 66.820 177.030 67.510 ;
        RECT 175.530 66.650 177.030 66.820 ;
        RECT 177.220 66.850 177.430 67.640 ;
        RECT 177.600 67.020 177.950 67.640 ;
        RECT 178.120 67.030 178.290 67.810 ;
        RECT 178.820 67.650 178.990 67.880 ;
        RECT 178.460 67.480 178.990 67.650 ;
        RECT 178.460 67.200 178.680 67.480 ;
        RECT 179.160 67.310 179.400 67.710 ;
        RECT 178.120 66.860 178.525 67.030 ;
        RECT 178.860 66.940 179.400 67.310 ;
        RECT 179.570 67.525 179.890 67.880 ;
        RECT 180.135 67.800 180.440 68.260 ;
        RECT 180.610 67.550 180.860 68.080 ;
        RECT 179.570 67.350 179.895 67.525 ;
        RECT 179.570 67.050 180.485 67.350 ;
        RECT 179.745 67.020 180.485 67.050 ;
        RECT 177.220 66.690 177.895 66.850 ;
        RECT 178.355 66.770 178.525 66.860 ;
        RECT 177.220 66.680 178.185 66.690 ;
        RECT 176.860 66.510 177.030 66.650 ;
        RECT 173.605 65.710 173.855 66.170 ;
        RECT 174.025 65.880 174.275 66.210 ;
        RECT 174.490 65.880 175.170 66.210 ;
        RECT 175.340 66.310 176.415 66.480 ;
        RECT 176.860 66.340 177.420 66.510 ;
        RECT 177.725 66.390 178.185 66.680 ;
        RECT 178.355 66.600 179.575 66.770 ;
        RECT 175.340 65.970 175.510 66.310 ;
        RECT 175.745 65.710 176.075 66.140 ;
        RECT 176.245 65.970 176.415 66.310 ;
        RECT 176.710 65.710 177.080 66.170 ;
        RECT 177.250 65.880 177.420 66.340 ;
        RECT 178.355 66.220 178.525 66.600 ;
        RECT 179.745 66.430 179.915 67.020 ;
        RECT 180.655 66.900 180.860 67.550 ;
        RECT 181.030 67.505 181.280 68.260 ;
        RECT 181.500 67.490 185.010 68.260 ;
        RECT 185.270 67.710 185.440 68.090 ;
        RECT 185.620 67.880 185.950 68.260 ;
        RECT 185.270 67.540 185.935 67.710 ;
        RECT 186.130 67.585 186.390 68.090 ;
        RECT 181.500 66.970 183.150 67.490 ;
        RECT 177.655 65.880 178.525 66.220 ;
        RECT 179.115 66.260 179.915 66.430 ;
        RECT 178.695 65.710 178.945 66.170 ;
        RECT 179.115 65.970 179.285 66.260 ;
        RECT 179.465 65.710 179.795 66.090 ;
        RECT 180.135 65.710 180.440 66.850 ;
        RECT 180.610 66.020 180.860 66.900 ;
        RECT 181.030 65.710 181.280 66.850 ;
        RECT 183.320 66.800 185.010 67.320 ;
        RECT 185.200 66.990 185.530 67.360 ;
        RECT 185.765 67.285 185.935 67.540 ;
        RECT 185.765 66.955 186.050 67.285 ;
        RECT 185.765 66.810 185.935 66.955 ;
        RECT 181.500 65.710 185.010 66.800 ;
        RECT 185.270 66.640 185.935 66.810 ;
        RECT 186.220 66.785 186.390 67.585 ;
        RECT 186.650 67.710 186.820 68.090 ;
        RECT 187.000 67.880 187.330 68.260 ;
        RECT 186.650 67.540 187.315 67.710 ;
        RECT 187.510 67.585 187.770 68.090 ;
        RECT 186.580 66.990 186.910 67.360 ;
        RECT 187.145 67.285 187.315 67.540 ;
        RECT 187.145 66.955 187.430 67.285 ;
        RECT 187.145 66.810 187.315 66.955 ;
        RECT 185.270 65.880 185.440 66.640 ;
        RECT 185.620 65.710 185.950 66.470 ;
        RECT 186.120 65.880 186.390 66.785 ;
        RECT 186.650 66.640 187.315 66.810 ;
        RECT 187.600 66.785 187.770 67.585 ;
        RECT 187.940 67.535 188.230 68.260 ;
        RECT 188.405 67.710 188.660 68.000 ;
        RECT 188.830 67.880 189.160 68.260 ;
        RECT 188.405 67.540 189.155 67.710 ;
        RECT 186.650 65.880 186.820 66.640 ;
        RECT 187.000 65.710 187.330 66.470 ;
        RECT 187.500 65.880 187.770 66.785 ;
        RECT 187.940 65.710 188.230 66.875 ;
        RECT 188.405 66.720 188.755 67.370 ;
        RECT 188.925 66.550 189.155 67.540 ;
        RECT 188.405 66.380 189.155 66.550 ;
        RECT 188.405 65.880 188.660 66.380 ;
        RECT 188.830 65.710 189.160 66.210 ;
        RECT 189.330 65.880 189.500 68.000 ;
        RECT 189.860 67.900 190.190 68.260 ;
        RECT 190.360 67.870 190.855 68.040 ;
        RECT 191.060 67.870 191.915 68.040 ;
        RECT 189.730 66.680 190.190 67.730 ;
        RECT 189.670 65.895 189.995 66.680 ;
        RECT 190.360 66.510 190.530 67.870 ;
        RECT 190.700 66.960 191.050 67.580 ;
        RECT 191.220 67.360 191.575 67.580 ;
        RECT 191.220 66.770 191.390 67.360 ;
        RECT 191.745 67.160 191.915 67.870 ;
        RECT 192.790 67.800 193.120 68.260 ;
        RECT 193.330 67.900 193.680 68.070 ;
        RECT 192.120 67.330 192.910 67.580 ;
        RECT 193.330 67.510 193.590 67.900 ;
        RECT 193.900 67.810 194.850 68.090 ;
        RECT 195.020 67.820 195.210 68.260 ;
        RECT 195.380 67.880 196.450 68.050 ;
        RECT 193.080 67.160 193.250 67.340 ;
        RECT 190.360 66.340 190.755 66.510 ;
        RECT 190.925 66.380 191.390 66.770 ;
        RECT 191.560 66.990 193.250 67.160 ;
        RECT 190.585 66.210 190.755 66.340 ;
        RECT 191.560 66.210 191.730 66.990 ;
        RECT 193.420 66.820 193.590 67.510 ;
        RECT 192.090 66.650 193.590 66.820 ;
        RECT 193.780 66.850 193.990 67.640 ;
        RECT 194.160 67.020 194.510 67.640 ;
        RECT 194.680 67.030 194.850 67.810 ;
        RECT 195.380 67.650 195.550 67.880 ;
        RECT 195.020 67.480 195.550 67.650 ;
        RECT 195.020 67.200 195.240 67.480 ;
        RECT 195.720 67.310 195.960 67.710 ;
        RECT 194.680 66.860 195.085 67.030 ;
        RECT 195.420 66.940 195.960 67.310 ;
        RECT 196.130 67.525 196.450 67.880 ;
        RECT 196.695 67.800 197.000 68.260 ;
        RECT 197.170 67.550 197.420 68.080 ;
        RECT 196.130 67.350 196.455 67.525 ;
        RECT 196.130 67.050 197.045 67.350 ;
        RECT 196.305 67.020 197.045 67.050 ;
        RECT 193.780 66.690 194.455 66.850 ;
        RECT 194.915 66.770 195.085 66.860 ;
        RECT 193.780 66.680 194.745 66.690 ;
        RECT 193.420 66.510 193.590 66.650 ;
        RECT 190.165 65.710 190.415 66.170 ;
        RECT 190.585 65.880 190.835 66.210 ;
        RECT 191.050 65.880 191.730 66.210 ;
        RECT 191.900 66.310 192.975 66.480 ;
        RECT 193.420 66.340 193.980 66.510 ;
        RECT 194.285 66.390 194.745 66.680 ;
        RECT 194.915 66.600 196.135 66.770 ;
        RECT 191.900 65.970 192.070 66.310 ;
        RECT 192.305 65.710 192.635 66.140 ;
        RECT 192.805 65.970 192.975 66.310 ;
        RECT 193.270 65.710 193.640 66.170 ;
        RECT 193.810 65.880 193.980 66.340 ;
        RECT 194.915 66.220 195.085 66.600 ;
        RECT 196.305 66.430 196.475 67.020 ;
        RECT 197.215 66.900 197.420 67.550 ;
        RECT 197.590 67.505 197.840 68.260 ;
        RECT 198.065 67.520 198.320 68.090 ;
        RECT 198.490 67.860 198.820 68.260 ;
        RECT 199.245 67.725 199.775 68.090 ;
        RECT 199.965 67.920 200.240 68.090 ;
        RECT 199.960 67.750 200.240 67.920 ;
        RECT 199.245 67.690 199.420 67.725 ;
        RECT 198.490 67.520 199.420 67.690 ;
        RECT 194.215 65.880 195.085 66.220 ;
        RECT 195.675 66.260 196.475 66.430 ;
        RECT 195.255 65.710 195.505 66.170 ;
        RECT 195.675 65.970 195.845 66.260 ;
        RECT 196.025 65.710 196.355 66.090 ;
        RECT 196.695 65.710 197.000 66.850 ;
        RECT 197.170 66.020 197.420 66.900 ;
        RECT 198.065 66.850 198.235 67.520 ;
        RECT 198.490 67.350 198.660 67.520 ;
        RECT 198.405 67.020 198.660 67.350 ;
        RECT 198.885 67.020 199.080 67.350 ;
        RECT 197.590 65.710 197.840 66.850 ;
        RECT 198.065 65.880 198.400 66.850 ;
        RECT 198.570 65.710 198.740 66.850 ;
        RECT 198.910 66.050 199.080 67.020 ;
        RECT 199.250 66.390 199.420 67.520 ;
        RECT 199.590 66.730 199.760 67.530 ;
        RECT 199.965 66.930 200.240 67.750 ;
        RECT 200.410 66.730 200.600 68.090 ;
        RECT 200.780 67.725 201.290 68.260 ;
        RECT 201.510 67.450 201.755 68.055 ;
        RECT 202.200 67.490 203.870 68.260 ;
        RECT 204.510 67.520 204.800 68.260 ;
        RECT 200.800 67.280 202.030 67.450 ;
        RECT 199.590 66.560 200.600 66.730 ;
        RECT 200.770 66.715 201.520 66.905 ;
        RECT 199.250 66.220 200.375 66.390 ;
        RECT 200.770 66.050 200.940 66.715 ;
        RECT 201.690 66.470 202.030 67.280 ;
        RECT 202.200 66.970 202.950 67.490 ;
        RECT 204.970 67.440 205.325 67.965 ;
        RECT 205.535 67.450 205.740 68.260 ;
        RECT 205.910 67.620 206.240 68.090 ;
        RECT 206.410 67.790 207.140 68.260 ;
        RECT 207.310 67.620 207.640 68.090 ;
        RECT 207.810 67.790 207.980 68.260 ;
        RECT 208.150 67.620 208.480 68.090 ;
        RECT 205.910 67.440 208.480 67.620 ;
        RECT 208.650 67.440 208.925 68.260 ;
        RECT 209.110 67.520 209.400 68.260 ;
        RECT 209.570 67.440 209.925 67.965 ;
        RECT 210.135 67.450 210.340 68.260 ;
        RECT 210.510 67.620 210.840 68.090 ;
        RECT 211.010 67.790 211.740 68.260 ;
        RECT 211.910 67.620 212.240 68.090 ;
        RECT 212.410 67.790 212.580 68.260 ;
        RECT 212.750 67.620 213.080 68.090 ;
        RECT 210.510 67.440 213.080 67.620 ;
        RECT 213.250 67.440 213.525 68.260 ;
        RECT 213.700 67.535 213.990 68.260 ;
        RECT 214.160 67.760 214.460 68.090 ;
        RECT 214.630 67.780 214.905 68.260 ;
        RECT 203.120 66.800 203.870 67.320 ;
        RECT 205.155 67.270 205.325 67.440 ;
        RECT 204.500 67.060 204.985 67.270 ;
        RECT 205.155 67.060 205.780 67.270 ;
        RECT 205.155 66.890 205.325 67.060 ;
        RECT 198.910 65.880 200.940 66.050 ;
        RECT 201.110 65.710 201.280 66.470 ;
        RECT 201.515 66.060 202.030 66.470 ;
        RECT 202.200 65.710 203.870 66.800 ;
        RECT 204.550 65.710 204.800 66.805 ;
        RECT 204.970 66.475 205.325 66.890 ;
        RECT 205.535 66.050 205.780 66.890 ;
        RECT 205.950 66.220 206.200 67.440 ;
        RECT 209.755 67.270 209.925 67.440 ;
        RECT 206.375 67.060 207.880 67.270 ;
        RECT 208.050 67.060 208.905 67.270 ;
        RECT 209.100 67.060 209.585 67.270 ;
        RECT 209.755 67.060 210.380 67.270 ;
        RECT 209.755 66.890 209.925 67.060 ;
        RECT 206.370 66.050 206.640 66.890 ;
        RECT 206.930 66.720 208.925 66.890 ;
        RECT 206.930 66.220 207.180 66.720 ;
        RECT 207.350 66.050 207.600 66.550 ;
        RECT 205.535 65.880 207.600 66.050 ;
        RECT 207.770 65.880 208.020 66.720 ;
        RECT 208.190 65.710 208.440 66.550 ;
        RECT 208.610 65.880 208.925 66.720 ;
        RECT 209.150 65.710 209.400 66.805 ;
        RECT 209.570 66.475 209.925 66.890 ;
        RECT 210.135 66.050 210.380 66.890 ;
        RECT 210.550 66.220 210.800 67.440 ;
        RECT 210.975 67.060 212.480 67.270 ;
        RECT 212.650 67.060 213.505 67.270 ;
        RECT 210.970 66.050 211.240 66.890 ;
        RECT 211.530 66.720 213.525 66.890 ;
        RECT 211.530 66.220 211.780 66.720 ;
        RECT 211.950 66.050 212.200 66.550 ;
        RECT 210.135 65.880 212.200 66.050 ;
        RECT 212.370 65.880 212.620 66.720 ;
        RECT 212.790 65.710 213.040 66.550 ;
        RECT 213.210 65.880 213.525 66.720 ;
        RECT 213.700 65.710 213.990 66.875 ;
        RECT 214.160 66.850 214.330 67.760 ;
        RECT 215.085 67.610 215.380 68.000 ;
        RECT 215.550 67.780 215.805 68.260 ;
        RECT 215.980 67.610 216.240 68.000 ;
        RECT 216.410 67.780 216.690 68.260 ;
        RECT 214.500 67.020 214.850 67.590 ;
        RECT 215.085 67.440 216.735 67.610 ;
        RECT 215.020 67.100 216.160 67.270 ;
        RECT 215.020 66.850 215.190 67.100 ;
        RECT 216.330 66.930 216.735 67.440 ;
        RECT 216.920 67.490 220.430 68.260 ;
        RECT 216.920 66.970 218.570 67.490 ;
        RECT 214.160 66.680 215.190 66.850 ;
        RECT 215.980 66.760 216.735 66.930 ;
        RECT 218.740 66.800 220.430 67.320 ;
        RECT 214.160 65.880 214.470 66.680 ;
        RECT 215.980 66.510 216.240 66.760 ;
        RECT 214.640 65.710 214.950 66.510 ;
        RECT 215.120 66.340 216.240 66.510 ;
        RECT 215.120 65.880 215.380 66.340 ;
        RECT 215.550 65.710 215.805 66.170 ;
        RECT 215.980 65.880 216.240 66.340 ;
        RECT 216.410 65.710 216.695 66.580 ;
        RECT 216.920 65.710 220.430 66.800 ;
        RECT 221.540 66.680 221.770 68.020 ;
        RECT 221.950 67.180 222.180 68.080 ;
        RECT 222.380 67.480 222.625 68.260 ;
        RECT 222.795 67.720 223.225 68.080 ;
        RECT 223.805 67.890 224.535 68.260 ;
        RECT 222.795 67.530 224.535 67.720 ;
        RECT 222.795 67.300 223.015 67.530 ;
        RECT 221.950 66.500 222.290 67.180 ;
        RECT 221.540 66.300 222.290 66.500 ;
        RECT 222.470 67.000 223.015 67.300 ;
        RECT 221.540 65.910 221.780 66.300 ;
        RECT 221.950 65.710 222.300 66.120 ;
        RECT 222.470 65.890 222.800 67.000 ;
        RECT 223.185 66.730 223.610 67.350 ;
        RECT 223.805 66.730 224.065 67.350 ;
        RECT 224.275 67.020 224.535 67.530 ;
        RECT 222.970 66.360 223.995 66.560 ;
        RECT 222.970 65.890 223.150 66.360 ;
        RECT 223.320 65.710 223.650 66.190 ;
        RECT 223.825 65.890 223.995 66.360 ;
        RECT 224.260 65.710 224.545 66.850 ;
        RECT 224.735 65.890 225.015 68.080 ;
        RECT 225.205 67.495 225.660 68.260 ;
        RECT 225.935 67.880 227.235 68.090 ;
        RECT 227.490 67.900 227.820 68.260 ;
        RECT 227.065 67.730 227.235 67.880 ;
        RECT 227.990 67.760 228.250 68.090 ;
        RECT 228.020 67.750 228.250 67.760 ;
        RECT 226.135 67.270 226.355 67.670 ;
        RECT 225.200 67.070 225.690 67.270 ;
        RECT 225.880 67.060 226.355 67.270 ;
        RECT 226.600 67.270 226.810 67.670 ;
        RECT 227.065 67.605 227.820 67.730 ;
        RECT 227.065 67.560 227.910 67.605 ;
        RECT 227.640 67.440 227.910 67.560 ;
        RECT 226.600 67.060 226.930 67.270 ;
        RECT 227.100 67.000 227.510 67.305 ;
        RECT 225.205 66.830 226.380 66.890 ;
        RECT 227.740 66.865 227.910 67.440 ;
        RECT 227.710 66.830 227.910 66.865 ;
        RECT 225.205 66.720 227.910 66.830 ;
        RECT 225.205 66.100 225.460 66.720 ;
        RECT 226.050 66.660 227.850 66.720 ;
        RECT 226.050 66.630 226.380 66.660 ;
        RECT 228.080 66.560 228.250 67.750 ;
        RECT 225.710 66.460 225.895 66.550 ;
        RECT 226.485 66.460 227.320 66.470 ;
        RECT 225.710 66.260 227.320 66.460 ;
        RECT 225.710 66.220 225.940 66.260 ;
        RECT 225.205 65.880 225.540 66.100 ;
        RECT 226.545 65.710 226.900 66.090 ;
        RECT 227.070 65.880 227.320 66.260 ;
        RECT 227.570 65.710 227.820 66.490 ;
        RECT 227.990 65.880 228.250 66.560 ;
        RECT 228.425 67.585 228.700 67.930 ;
        RECT 228.890 67.860 229.270 68.260 ;
        RECT 229.440 67.690 229.610 68.040 ;
        RECT 229.780 67.860 230.110 68.260 ;
        RECT 230.280 67.690 230.535 68.040 ;
        RECT 230.720 67.715 236.065 68.260 ;
        RECT 228.425 66.850 228.595 67.585 ;
        RECT 228.870 67.520 230.535 67.690 ;
        RECT 228.870 67.350 229.040 67.520 ;
        RECT 228.765 67.020 229.040 67.350 ;
        RECT 229.210 67.020 230.035 67.350 ;
        RECT 230.205 67.020 230.550 67.350 ;
        RECT 228.870 66.850 229.040 67.020 ;
        RECT 228.425 65.880 228.700 66.850 ;
        RECT 228.870 66.680 229.530 66.850 ;
        RECT 229.840 66.730 230.035 67.020 ;
        RECT 232.305 66.885 232.645 67.715 ;
        RECT 236.245 67.495 236.700 68.260 ;
        RECT 236.975 67.880 238.275 68.090 ;
        RECT 238.530 67.900 238.860 68.260 ;
        RECT 238.105 67.730 238.275 67.880 ;
        RECT 239.030 67.760 239.290 68.090 ;
        RECT 229.360 66.560 229.530 66.680 ;
        RECT 230.205 66.560 230.530 66.850 ;
        RECT 228.910 65.710 229.190 66.510 ;
        RECT 229.360 66.390 230.530 66.560 ;
        RECT 229.360 65.930 230.550 66.220 ;
        RECT 234.125 66.145 234.475 67.395 ;
        RECT 237.175 67.270 237.395 67.670 ;
        RECT 236.240 67.070 236.730 67.270 ;
        RECT 236.920 67.060 237.395 67.270 ;
        RECT 237.640 67.270 237.850 67.670 ;
        RECT 238.105 67.605 238.860 67.730 ;
        RECT 238.105 67.560 238.950 67.605 ;
        RECT 238.680 67.440 238.950 67.560 ;
        RECT 237.640 67.060 237.970 67.270 ;
        RECT 238.140 67.000 238.550 67.305 ;
        RECT 236.245 66.830 237.420 66.890 ;
        RECT 238.780 66.865 238.950 67.440 ;
        RECT 238.750 66.830 238.950 66.865 ;
        RECT 236.245 66.720 238.950 66.830 ;
        RECT 230.720 65.710 236.065 66.145 ;
        RECT 236.245 66.100 236.500 66.720 ;
        RECT 237.090 66.660 238.890 66.720 ;
        RECT 237.090 66.630 237.420 66.660 ;
        RECT 239.120 66.560 239.290 67.760 ;
        RECT 239.460 67.535 239.750 68.260 ;
        RECT 240.010 67.780 240.310 68.260 ;
        RECT 240.480 67.610 240.740 68.065 ;
        RECT 240.910 67.780 241.170 68.260 ;
        RECT 241.350 67.610 241.610 68.065 ;
        RECT 241.780 67.780 242.030 68.260 ;
        RECT 242.210 67.610 242.470 68.065 ;
        RECT 242.640 67.780 242.890 68.260 ;
        RECT 243.070 67.610 243.330 68.065 ;
        RECT 243.500 67.780 243.745 68.260 ;
        RECT 243.915 67.610 244.190 68.065 ;
        RECT 244.360 67.780 244.605 68.260 ;
        RECT 244.775 67.610 245.035 68.065 ;
        RECT 245.205 67.780 245.465 68.260 ;
        RECT 245.635 67.610 245.895 68.065 ;
        RECT 246.065 67.780 246.325 68.260 ;
        RECT 246.495 67.610 246.755 68.065 ;
        RECT 246.925 67.700 247.185 68.260 ;
        RECT 240.010 67.440 246.755 67.610 ;
        RECT 236.750 66.460 236.935 66.550 ;
        RECT 237.525 66.460 238.360 66.470 ;
        RECT 236.750 66.260 238.360 66.460 ;
        RECT 236.750 66.220 236.980 66.260 ;
        RECT 236.245 65.880 236.580 66.100 ;
        RECT 237.585 65.710 237.940 66.090 ;
        RECT 238.110 65.880 238.360 66.260 ;
        RECT 238.610 65.710 238.860 66.490 ;
        RECT 239.030 65.880 239.290 66.560 ;
        RECT 239.460 65.710 239.750 66.875 ;
        RECT 240.010 66.850 241.175 67.440 ;
        RECT 247.355 67.270 247.605 68.080 ;
        RECT 247.785 67.735 248.045 68.260 ;
        RECT 248.215 67.270 248.465 68.080 ;
        RECT 248.645 67.750 248.950 68.260 ;
        RECT 249.120 67.715 254.465 68.260 ;
        RECT 241.345 67.020 248.465 67.270 ;
        RECT 248.635 67.020 248.950 67.580 ;
        RECT 240.010 66.625 246.755 66.850 ;
        RECT 240.010 65.710 240.280 66.455 ;
        RECT 240.450 65.885 240.740 66.625 ;
        RECT 241.350 66.610 246.755 66.625 ;
        RECT 240.910 65.715 241.165 66.440 ;
        RECT 241.350 65.885 241.610 66.610 ;
        RECT 241.780 65.715 242.025 66.440 ;
        RECT 242.210 65.885 242.470 66.610 ;
        RECT 242.640 65.715 242.885 66.440 ;
        RECT 243.070 65.885 243.330 66.610 ;
        RECT 243.500 65.715 243.745 66.440 ;
        RECT 243.915 65.885 244.175 66.610 ;
        RECT 244.345 65.715 244.605 66.440 ;
        RECT 244.775 65.885 245.035 66.610 ;
        RECT 245.205 65.715 245.465 66.440 ;
        RECT 245.635 65.885 245.895 66.610 ;
        RECT 246.065 65.715 246.325 66.440 ;
        RECT 246.495 65.885 246.755 66.610 ;
        RECT 246.925 65.715 247.185 66.510 ;
        RECT 247.355 65.885 247.605 67.020 ;
        RECT 240.910 65.710 247.185 65.715 ;
        RECT 247.785 65.710 248.045 66.520 ;
        RECT 248.220 65.880 248.465 67.020 ;
        RECT 250.705 66.885 251.045 67.715 ;
        RECT 254.645 67.495 255.100 68.260 ;
        RECT 255.375 67.880 256.675 68.090 ;
        RECT 256.930 67.900 257.260 68.260 ;
        RECT 256.505 67.730 256.675 67.880 ;
        RECT 257.430 67.760 257.690 68.090 ;
        RECT 248.645 65.710 248.940 66.520 ;
        RECT 252.525 66.145 252.875 67.395 ;
        RECT 255.575 67.270 255.795 67.670 ;
        RECT 254.640 67.070 255.130 67.270 ;
        RECT 255.320 67.060 255.795 67.270 ;
        RECT 256.040 67.270 256.250 67.670 ;
        RECT 256.505 67.605 257.260 67.730 ;
        RECT 256.505 67.560 257.350 67.605 ;
        RECT 257.080 67.440 257.350 67.560 ;
        RECT 256.040 67.060 256.370 67.270 ;
        RECT 256.540 67.000 256.950 67.305 ;
        RECT 254.645 66.830 255.820 66.890 ;
        RECT 257.180 66.865 257.350 67.440 ;
        RECT 257.150 66.830 257.350 66.865 ;
        RECT 254.645 66.720 257.350 66.830 ;
        RECT 249.120 65.710 254.465 66.145 ;
        RECT 254.645 66.100 254.900 66.720 ;
        RECT 255.490 66.660 257.290 66.720 ;
        RECT 255.490 66.630 255.820 66.660 ;
        RECT 257.520 66.560 257.690 67.760 ;
        RECT 255.150 66.460 255.335 66.550 ;
        RECT 255.925 66.460 256.760 66.470 ;
        RECT 255.150 66.260 256.760 66.460 ;
        RECT 255.150 66.220 255.380 66.260 ;
        RECT 254.645 65.880 254.980 66.100 ;
        RECT 255.985 65.710 256.340 66.090 ;
        RECT 256.510 65.880 256.760 66.260 ;
        RECT 257.010 65.710 257.260 66.490 ;
        RECT 257.430 65.880 257.690 66.560 ;
        RECT 258.340 67.760 258.595 68.090 ;
        RECT 258.810 67.780 259.140 68.260 ;
        RECT 259.310 67.840 260.845 68.090 ;
        RECT 258.340 67.680 258.525 67.760 ;
        RECT 258.340 66.550 258.510 67.680 ;
        RECT 259.310 67.610 259.480 67.840 ;
        RECT 258.680 67.440 259.480 67.610 ;
        RECT 258.680 66.890 258.850 67.440 ;
        RECT 259.660 67.270 259.945 67.670 ;
        RECT 259.080 67.240 259.445 67.270 ;
        RECT 259.070 67.070 259.445 67.240 ;
        RECT 259.615 67.070 259.945 67.270 ;
        RECT 260.215 67.270 260.495 67.670 ;
        RECT 260.675 67.610 260.845 67.840 ;
        RECT 261.070 67.780 261.400 68.260 ;
        RECT 261.570 67.610 261.740 68.090 ;
        RECT 260.675 67.440 261.740 67.610 ;
        RECT 262.000 67.760 262.260 68.090 ;
        RECT 262.430 67.900 262.760 68.260 ;
        RECT 263.015 67.880 264.315 68.090 ;
        RECT 260.215 67.070 260.690 67.270 ;
        RECT 260.860 67.070 261.305 67.270 ;
        RECT 261.475 67.060 261.825 67.270 ;
        RECT 258.680 66.720 261.740 66.890 ;
        RECT 258.340 65.880 258.595 66.550 ;
        RECT 258.765 65.710 259.095 66.470 ;
        RECT 259.265 66.310 260.900 66.550 ;
        RECT 259.265 65.880 259.515 66.310 ;
        RECT 260.670 66.220 260.900 66.310 ;
        RECT 259.685 65.710 260.040 66.130 ;
        RECT 260.230 66.050 260.560 66.090 ;
        RECT 261.070 66.050 261.400 66.550 ;
        RECT 260.230 65.880 261.400 66.050 ;
        RECT 261.570 65.880 261.740 66.720 ;
        RECT 262.000 66.560 262.170 67.760 ;
        RECT 263.015 67.730 263.185 67.880 ;
        RECT 262.430 67.605 263.185 67.730 ;
        RECT 262.340 67.560 263.185 67.605 ;
        RECT 262.340 67.440 262.610 67.560 ;
        RECT 262.340 66.865 262.510 67.440 ;
        RECT 262.740 67.000 263.150 67.305 ;
        RECT 263.440 67.270 263.650 67.670 ;
        RECT 263.320 67.060 263.650 67.270 ;
        RECT 263.895 67.270 264.115 67.670 ;
        RECT 264.590 67.495 265.045 68.260 ;
        RECT 265.220 67.535 265.510 68.260 ;
        RECT 265.680 67.490 268.270 68.260 ;
        RECT 268.990 67.710 269.160 68.090 ;
        RECT 269.340 67.880 269.670 68.260 ;
        RECT 268.990 67.540 269.655 67.710 ;
        RECT 269.850 67.585 270.110 68.090 ;
        RECT 263.895 67.060 264.370 67.270 ;
        RECT 264.560 67.070 265.050 67.270 ;
        RECT 265.680 66.970 266.890 67.490 ;
        RECT 262.340 66.830 262.540 66.865 ;
        RECT 263.870 66.830 265.045 66.890 ;
        RECT 262.340 66.720 265.045 66.830 ;
        RECT 262.400 66.660 264.200 66.720 ;
        RECT 263.870 66.630 264.200 66.660 ;
        RECT 262.000 65.880 262.260 66.560 ;
        RECT 262.430 65.710 262.680 66.490 ;
        RECT 262.930 66.460 263.765 66.470 ;
        RECT 264.355 66.460 264.540 66.550 ;
        RECT 262.930 66.260 264.540 66.460 ;
        RECT 262.930 65.880 263.180 66.260 ;
        RECT 264.310 66.220 264.540 66.260 ;
        RECT 264.790 66.100 265.045 66.720 ;
        RECT 263.350 65.710 263.705 66.090 ;
        RECT 264.710 65.880 265.045 66.100 ;
        RECT 265.220 65.710 265.510 66.875 ;
        RECT 267.060 66.800 268.270 67.320 ;
        RECT 268.920 66.990 269.250 67.360 ;
        RECT 269.485 67.285 269.655 67.540 ;
        RECT 269.485 66.955 269.770 67.285 ;
        RECT 269.485 66.810 269.655 66.955 ;
        RECT 265.680 65.710 268.270 66.800 ;
        RECT 268.990 66.640 269.655 66.810 ;
        RECT 269.940 66.785 270.110 67.585 ;
        RECT 270.285 67.710 270.540 68.000 ;
        RECT 270.710 67.880 271.040 68.260 ;
        RECT 270.285 67.540 271.035 67.710 ;
        RECT 268.990 65.880 269.160 66.640 ;
        RECT 269.340 65.710 269.670 66.470 ;
        RECT 269.840 65.880 270.110 66.785 ;
        RECT 270.285 66.720 270.635 67.370 ;
        RECT 270.805 66.550 271.035 67.540 ;
        RECT 270.285 66.380 271.035 66.550 ;
        RECT 270.285 65.880 270.540 66.380 ;
        RECT 270.710 65.710 271.040 66.210 ;
        RECT 271.210 65.880 271.380 68.000 ;
        RECT 271.740 67.900 272.070 68.260 ;
        RECT 272.240 67.870 272.735 68.040 ;
        RECT 272.940 67.870 273.795 68.040 ;
        RECT 271.610 66.680 272.070 67.730 ;
        RECT 271.550 65.895 271.875 66.680 ;
        RECT 272.240 66.510 272.410 67.870 ;
        RECT 272.580 66.960 272.930 67.580 ;
        RECT 273.100 67.360 273.455 67.580 ;
        RECT 273.100 66.770 273.270 67.360 ;
        RECT 273.625 67.160 273.795 67.870 ;
        RECT 274.670 67.800 275.000 68.260 ;
        RECT 275.210 67.900 275.560 68.070 ;
        RECT 274.000 67.330 274.790 67.580 ;
        RECT 275.210 67.510 275.470 67.900 ;
        RECT 275.780 67.810 276.730 68.090 ;
        RECT 276.900 67.820 277.090 68.260 ;
        RECT 277.260 67.880 278.330 68.050 ;
        RECT 274.960 67.160 275.130 67.340 ;
        RECT 272.240 66.340 272.635 66.510 ;
        RECT 272.805 66.380 273.270 66.770 ;
        RECT 273.440 66.990 275.130 67.160 ;
        RECT 272.465 66.210 272.635 66.340 ;
        RECT 273.440 66.210 273.610 66.990 ;
        RECT 275.300 66.820 275.470 67.510 ;
        RECT 273.970 66.650 275.470 66.820 ;
        RECT 275.660 66.850 275.870 67.640 ;
        RECT 276.040 67.020 276.390 67.640 ;
        RECT 276.560 67.030 276.730 67.810 ;
        RECT 277.260 67.650 277.430 67.880 ;
        RECT 276.900 67.480 277.430 67.650 ;
        RECT 276.900 67.200 277.120 67.480 ;
        RECT 277.600 67.310 277.840 67.710 ;
        RECT 276.560 66.860 276.965 67.030 ;
        RECT 277.300 66.940 277.840 67.310 ;
        RECT 278.010 67.525 278.330 67.880 ;
        RECT 278.575 67.800 278.880 68.260 ;
        RECT 279.050 67.550 279.300 68.080 ;
        RECT 278.010 67.350 278.335 67.525 ;
        RECT 278.010 67.050 278.925 67.350 ;
        RECT 278.185 67.020 278.925 67.050 ;
        RECT 275.660 66.690 276.335 66.850 ;
        RECT 276.795 66.770 276.965 66.860 ;
        RECT 275.660 66.680 276.625 66.690 ;
        RECT 275.300 66.510 275.470 66.650 ;
        RECT 272.045 65.710 272.295 66.170 ;
        RECT 272.465 65.880 272.715 66.210 ;
        RECT 272.930 65.880 273.610 66.210 ;
        RECT 273.780 66.310 274.855 66.480 ;
        RECT 275.300 66.340 275.860 66.510 ;
        RECT 276.165 66.390 276.625 66.680 ;
        RECT 276.795 66.600 278.015 66.770 ;
        RECT 273.780 65.970 273.950 66.310 ;
        RECT 274.185 65.710 274.515 66.140 ;
        RECT 274.685 65.970 274.855 66.310 ;
        RECT 275.150 65.710 275.520 66.170 ;
        RECT 275.690 65.880 275.860 66.340 ;
        RECT 276.795 66.220 276.965 66.600 ;
        RECT 278.185 66.430 278.355 67.020 ;
        RECT 279.095 66.900 279.300 67.550 ;
        RECT 279.470 67.505 279.720 68.260 ;
        RECT 280.405 67.710 280.660 68.000 ;
        RECT 280.830 67.880 281.160 68.260 ;
        RECT 280.405 67.540 281.155 67.710 ;
        RECT 276.095 65.880 276.965 66.220 ;
        RECT 277.555 66.260 278.355 66.430 ;
        RECT 277.135 65.710 277.385 66.170 ;
        RECT 277.555 65.970 277.725 66.260 ;
        RECT 277.905 65.710 278.235 66.090 ;
        RECT 278.575 65.710 278.880 66.850 ;
        RECT 279.050 66.020 279.300 66.900 ;
        RECT 279.470 65.710 279.720 66.850 ;
        RECT 280.405 66.720 280.755 67.370 ;
        RECT 280.925 66.550 281.155 67.540 ;
        RECT 280.405 66.380 281.155 66.550 ;
        RECT 280.405 65.880 280.660 66.380 ;
        RECT 280.830 65.710 281.160 66.210 ;
        RECT 281.330 65.880 281.500 68.000 ;
        RECT 281.860 67.900 282.190 68.260 ;
        RECT 282.360 67.870 282.855 68.040 ;
        RECT 283.060 67.870 283.915 68.040 ;
        RECT 281.730 66.680 282.190 67.730 ;
        RECT 281.670 65.895 281.995 66.680 ;
        RECT 282.360 66.510 282.530 67.870 ;
        RECT 282.700 66.960 283.050 67.580 ;
        RECT 283.220 67.360 283.575 67.580 ;
        RECT 283.220 66.770 283.390 67.360 ;
        RECT 283.745 67.160 283.915 67.870 ;
        RECT 284.790 67.800 285.120 68.260 ;
        RECT 285.330 67.900 285.680 68.070 ;
        RECT 284.120 67.330 284.910 67.580 ;
        RECT 285.330 67.510 285.590 67.900 ;
        RECT 285.900 67.810 286.850 68.090 ;
        RECT 287.020 67.820 287.210 68.260 ;
        RECT 287.380 67.880 288.450 68.050 ;
        RECT 285.080 67.160 285.250 67.340 ;
        RECT 282.360 66.340 282.755 66.510 ;
        RECT 282.925 66.380 283.390 66.770 ;
        RECT 283.560 66.990 285.250 67.160 ;
        RECT 282.585 66.210 282.755 66.340 ;
        RECT 283.560 66.210 283.730 66.990 ;
        RECT 285.420 66.820 285.590 67.510 ;
        RECT 284.090 66.650 285.590 66.820 ;
        RECT 285.780 66.850 285.990 67.640 ;
        RECT 286.160 67.020 286.510 67.640 ;
        RECT 286.680 67.030 286.850 67.810 ;
        RECT 287.380 67.650 287.550 67.880 ;
        RECT 287.020 67.480 287.550 67.650 ;
        RECT 287.020 67.200 287.240 67.480 ;
        RECT 287.720 67.310 287.960 67.710 ;
        RECT 286.680 66.860 287.085 67.030 ;
        RECT 287.420 66.940 287.960 67.310 ;
        RECT 288.130 67.525 288.450 67.880 ;
        RECT 288.695 67.800 289.000 68.260 ;
        RECT 289.170 67.550 289.425 68.080 ;
        RECT 288.130 67.350 288.455 67.525 ;
        RECT 288.130 67.050 289.045 67.350 ;
        RECT 288.305 67.020 289.045 67.050 ;
        RECT 285.780 66.690 286.455 66.850 ;
        RECT 286.915 66.770 287.085 66.860 ;
        RECT 285.780 66.680 286.745 66.690 ;
        RECT 285.420 66.510 285.590 66.650 ;
        RECT 282.165 65.710 282.415 66.170 ;
        RECT 282.585 65.880 282.835 66.210 ;
        RECT 283.050 65.880 283.730 66.210 ;
        RECT 283.900 66.310 284.975 66.480 ;
        RECT 285.420 66.340 285.980 66.510 ;
        RECT 286.285 66.390 286.745 66.680 ;
        RECT 286.915 66.600 288.135 66.770 ;
        RECT 283.900 65.970 284.070 66.310 ;
        RECT 284.305 65.710 284.635 66.140 ;
        RECT 284.805 65.970 284.975 66.310 ;
        RECT 285.270 65.710 285.640 66.170 ;
        RECT 285.810 65.880 285.980 66.340 ;
        RECT 286.915 66.220 287.085 66.600 ;
        RECT 288.305 66.430 288.475 67.020 ;
        RECT 289.215 66.900 289.425 67.550 ;
        RECT 289.600 67.510 290.810 68.260 ;
        RECT 290.980 67.535 291.270 68.260 ;
        RECT 289.600 66.970 290.120 67.510 ;
        RECT 291.440 67.490 293.110 68.260 ;
        RECT 293.830 67.710 294.000 68.090 ;
        RECT 294.180 67.880 294.510 68.260 ;
        RECT 293.830 67.540 294.495 67.710 ;
        RECT 294.690 67.585 294.950 68.090 ;
        RECT 286.215 65.880 287.085 66.220 ;
        RECT 287.675 66.260 288.475 66.430 ;
        RECT 287.255 65.710 287.505 66.170 ;
        RECT 287.675 65.970 287.845 66.260 ;
        RECT 288.025 65.710 288.355 66.090 ;
        RECT 288.695 65.710 289.000 66.850 ;
        RECT 289.170 66.020 289.425 66.900 ;
        RECT 290.290 66.800 290.810 67.340 ;
        RECT 291.440 66.970 292.190 67.490 ;
        RECT 289.600 65.710 290.810 66.800 ;
        RECT 290.980 65.710 291.270 66.875 ;
        RECT 292.360 66.800 293.110 67.320 ;
        RECT 293.760 66.990 294.090 67.360 ;
        RECT 294.325 67.285 294.495 67.540 ;
        RECT 294.325 66.955 294.610 67.285 ;
        RECT 294.325 66.810 294.495 66.955 ;
        RECT 291.440 65.710 293.110 66.800 ;
        RECT 293.830 66.640 294.495 66.810 ;
        RECT 294.780 66.785 294.950 67.585 ;
        RECT 295.125 67.710 295.380 68.000 ;
        RECT 295.550 67.880 295.880 68.260 ;
        RECT 295.125 67.540 295.875 67.710 ;
        RECT 293.830 65.880 294.000 66.640 ;
        RECT 294.180 65.710 294.510 66.470 ;
        RECT 294.680 65.880 294.950 66.785 ;
        RECT 295.125 66.720 295.475 67.370 ;
        RECT 295.645 66.550 295.875 67.540 ;
        RECT 295.125 66.380 295.875 66.550 ;
        RECT 295.125 65.880 295.380 66.380 ;
        RECT 295.550 65.710 295.880 66.210 ;
        RECT 296.050 65.880 296.220 68.000 ;
        RECT 296.580 67.900 296.910 68.260 ;
        RECT 297.080 67.870 297.575 68.040 ;
        RECT 297.780 67.870 298.635 68.040 ;
        RECT 296.450 66.680 296.910 67.730 ;
        RECT 296.390 65.895 296.715 66.680 ;
        RECT 297.080 66.510 297.250 67.870 ;
        RECT 297.420 66.960 297.770 67.580 ;
        RECT 297.940 67.360 298.295 67.580 ;
        RECT 297.940 66.770 298.110 67.360 ;
        RECT 298.465 67.160 298.635 67.870 ;
        RECT 299.510 67.800 299.840 68.260 ;
        RECT 300.050 67.900 300.400 68.070 ;
        RECT 298.840 67.330 299.630 67.580 ;
        RECT 300.050 67.510 300.310 67.900 ;
        RECT 300.620 67.810 301.570 68.090 ;
        RECT 301.740 67.820 301.930 68.260 ;
        RECT 302.100 67.880 303.170 68.050 ;
        RECT 299.800 67.160 299.970 67.340 ;
        RECT 297.080 66.340 297.475 66.510 ;
        RECT 297.645 66.380 298.110 66.770 ;
        RECT 298.280 66.990 299.970 67.160 ;
        RECT 297.305 66.210 297.475 66.340 ;
        RECT 298.280 66.210 298.450 66.990 ;
        RECT 300.140 66.820 300.310 67.510 ;
        RECT 298.810 66.650 300.310 66.820 ;
        RECT 300.500 66.850 300.710 67.640 ;
        RECT 300.880 67.020 301.230 67.640 ;
        RECT 301.400 67.030 301.570 67.810 ;
        RECT 302.100 67.650 302.270 67.880 ;
        RECT 301.740 67.480 302.270 67.650 ;
        RECT 301.740 67.200 301.960 67.480 ;
        RECT 302.440 67.310 302.680 67.710 ;
        RECT 301.400 66.860 301.805 67.030 ;
        RECT 302.140 66.940 302.680 67.310 ;
        RECT 302.850 67.525 303.170 67.880 ;
        RECT 303.415 67.800 303.720 68.260 ;
        RECT 303.890 67.550 304.140 68.080 ;
        RECT 302.850 67.350 303.175 67.525 ;
        RECT 302.850 67.050 303.765 67.350 ;
        RECT 303.025 67.020 303.765 67.050 ;
        RECT 300.500 66.690 301.175 66.850 ;
        RECT 301.635 66.770 301.805 66.860 ;
        RECT 300.500 66.680 301.465 66.690 ;
        RECT 300.140 66.510 300.310 66.650 ;
        RECT 296.885 65.710 297.135 66.170 ;
        RECT 297.305 65.880 297.555 66.210 ;
        RECT 297.770 65.880 298.450 66.210 ;
        RECT 298.620 66.310 299.695 66.480 ;
        RECT 300.140 66.340 300.700 66.510 ;
        RECT 301.005 66.390 301.465 66.680 ;
        RECT 301.635 66.600 302.855 66.770 ;
        RECT 298.620 65.970 298.790 66.310 ;
        RECT 299.025 65.710 299.355 66.140 ;
        RECT 299.525 65.970 299.695 66.310 ;
        RECT 299.990 65.710 300.360 66.170 ;
        RECT 300.530 65.880 300.700 66.340 ;
        RECT 301.635 66.220 301.805 66.600 ;
        RECT 303.025 66.430 303.195 67.020 ;
        RECT 303.935 66.900 304.140 67.550 ;
        RECT 304.310 67.505 304.560 68.260 ;
        RECT 304.840 67.780 305.120 68.260 ;
        RECT 305.290 67.610 305.550 68.000 ;
        RECT 305.725 67.780 305.980 68.260 ;
        RECT 306.150 67.610 306.445 68.000 ;
        RECT 306.625 67.780 306.900 68.260 ;
        RECT 307.070 67.760 307.370 68.090 ;
        RECT 300.935 65.880 301.805 66.220 ;
        RECT 302.395 66.260 303.195 66.430 ;
        RECT 301.975 65.710 302.225 66.170 ;
        RECT 302.395 65.970 302.565 66.260 ;
        RECT 302.745 65.710 303.075 66.090 ;
        RECT 303.415 65.710 303.720 66.850 ;
        RECT 303.890 66.020 304.140 66.900 ;
        RECT 304.795 67.440 306.445 67.610 ;
        RECT 304.795 66.930 305.200 67.440 ;
        RECT 305.370 67.100 306.510 67.270 ;
        RECT 304.310 65.710 304.560 66.850 ;
        RECT 304.795 66.760 305.550 66.930 ;
        RECT 304.835 65.710 305.120 66.580 ;
        RECT 305.290 66.510 305.550 66.760 ;
        RECT 306.340 66.850 306.510 67.100 ;
        RECT 306.680 67.020 307.030 67.590 ;
        RECT 307.200 66.850 307.370 67.760 ;
        RECT 307.540 67.490 309.210 68.260 ;
        RECT 309.840 67.510 311.050 68.260 ;
        RECT 307.540 66.970 308.290 67.490 ;
        RECT 306.340 66.680 307.370 66.850 ;
        RECT 308.460 66.800 309.210 67.320 ;
        RECT 305.290 66.340 306.410 66.510 ;
        RECT 305.290 65.880 305.550 66.340 ;
        RECT 305.725 65.710 305.980 66.170 ;
        RECT 306.150 65.880 306.410 66.340 ;
        RECT 306.580 65.710 306.890 66.510 ;
        RECT 307.060 65.880 307.370 66.680 ;
        RECT 307.540 65.710 309.210 66.800 ;
        RECT 309.840 66.800 310.360 67.340 ;
        RECT 310.530 66.970 311.050 67.510 ;
        RECT 309.840 65.710 311.050 66.800 ;
        RECT 162.095 65.540 311.135 65.710 ;
        RECT 162.180 64.450 163.390 65.540 ;
        RECT 163.560 64.450 165.230 65.540 ;
        RECT 165.405 64.870 165.660 65.370 ;
        RECT 165.830 65.040 166.160 65.540 ;
        RECT 165.405 64.700 166.155 64.870 ;
        RECT 162.180 63.740 162.700 64.280 ;
        RECT 162.870 63.910 163.390 64.450 ;
        RECT 163.560 63.760 164.310 64.280 ;
        RECT 164.480 63.930 165.230 64.450 ;
        RECT 165.405 63.880 165.755 64.530 ;
        RECT 162.180 62.990 163.390 63.740 ;
        RECT 163.560 62.990 165.230 63.760 ;
        RECT 165.925 63.710 166.155 64.700 ;
        RECT 165.405 63.540 166.155 63.710 ;
        RECT 165.405 63.250 165.660 63.540 ;
        RECT 165.830 62.990 166.160 63.370 ;
        RECT 166.330 63.250 166.500 65.370 ;
        RECT 166.670 64.570 166.995 65.355 ;
        RECT 167.165 65.080 167.415 65.540 ;
        RECT 167.585 65.040 167.835 65.370 ;
        RECT 168.050 65.040 168.730 65.370 ;
        RECT 167.585 64.910 167.755 65.040 ;
        RECT 167.360 64.740 167.755 64.910 ;
        RECT 166.730 63.520 167.190 64.570 ;
        RECT 167.360 63.380 167.530 64.740 ;
        RECT 167.925 64.480 168.390 64.870 ;
        RECT 167.700 63.670 168.050 64.290 ;
        RECT 168.220 63.890 168.390 64.480 ;
        RECT 168.560 64.260 168.730 65.040 ;
        RECT 168.900 64.940 169.070 65.280 ;
        RECT 169.305 65.110 169.635 65.540 ;
        RECT 169.805 64.940 169.975 65.280 ;
        RECT 170.270 65.080 170.640 65.540 ;
        RECT 168.900 64.770 169.975 64.940 ;
        RECT 170.810 64.910 170.980 65.370 ;
        RECT 171.215 65.030 172.085 65.370 ;
        RECT 172.255 65.080 172.505 65.540 ;
        RECT 170.420 64.740 170.980 64.910 ;
        RECT 170.420 64.600 170.590 64.740 ;
        RECT 169.090 64.430 170.590 64.600 ;
        RECT 171.285 64.570 171.745 64.860 ;
        RECT 168.560 64.090 170.250 64.260 ;
        RECT 168.220 63.670 168.575 63.890 ;
        RECT 168.745 63.380 168.915 64.090 ;
        RECT 169.120 63.670 169.910 63.920 ;
        RECT 170.080 63.910 170.250 64.090 ;
        RECT 170.420 63.740 170.590 64.430 ;
        RECT 166.860 62.990 167.190 63.350 ;
        RECT 167.360 63.210 167.855 63.380 ;
        RECT 168.060 63.210 168.915 63.380 ;
        RECT 169.790 62.990 170.120 63.450 ;
        RECT 170.330 63.350 170.590 63.740 ;
        RECT 170.780 64.560 171.745 64.570 ;
        RECT 171.915 64.650 172.085 65.030 ;
        RECT 172.675 64.990 172.845 65.280 ;
        RECT 173.025 65.160 173.355 65.540 ;
        RECT 172.675 64.820 173.475 64.990 ;
        RECT 170.780 64.400 171.455 64.560 ;
        RECT 171.915 64.480 173.135 64.650 ;
        RECT 170.780 63.610 170.990 64.400 ;
        RECT 171.915 64.390 172.085 64.480 ;
        RECT 171.160 63.610 171.510 64.230 ;
        RECT 171.680 64.220 172.085 64.390 ;
        RECT 171.680 63.440 171.850 64.220 ;
        RECT 172.020 63.770 172.240 64.050 ;
        RECT 172.420 63.940 172.960 64.310 ;
        RECT 173.305 64.230 173.475 64.820 ;
        RECT 173.695 64.400 174.000 65.540 ;
        RECT 174.170 64.350 174.420 65.230 ;
        RECT 174.590 64.400 174.840 65.540 ;
        RECT 175.060 64.375 175.350 65.540 ;
        RECT 175.525 64.400 175.860 65.370 ;
        RECT 176.030 64.400 176.200 65.540 ;
        RECT 176.370 65.200 178.400 65.370 ;
        RECT 173.305 64.200 174.045 64.230 ;
        RECT 172.020 63.600 172.550 63.770 ;
        RECT 170.330 63.180 170.680 63.350 ;
        RECT 170.900 63.160 171.850 63.440 ;
        RECT 172.020 62.990 172.210 63.430 ;
        RECT 172.380 63.370 172.550 63.600 ;
        RECT 172.720 63.540 172.960 63.940 ;
        RECT 173.130 63.900 174.045 64.200 ;
        RECT 173.130 63.725 173.455 63.900 ;
        RECT 173.130 63.370 173.450 63.725 ;
        RECT 174.215 63.700 174.420 64.350 ;
        RECT 172.380 63.200 173.450 63.370 ;
        RECT 173.695 62.990 174.000 63.450 ;
        RECT 174.170 63.170 174.420 63.700 ;
        RECT 174.590 62.990 174.840 63.745 ;
        RECT 175.525 63.730 175.695 64.400 ;
        RECT 176.370 64.230 176.540 65.200 ;
        RECT 175.865 63.900 176.120 64.230 ;
        RECT 176.345 63.900 176.540 64.230 ;
        RECT 176.710 64.860 177.835 65.030 ;
        RECT 175.950 63.730 176.120 63.900 ;
        RECT 176.710 63.730 176.880 64.860 ;
        RECT 175.060 62.990 175.350 63.715 ;
        RECT 175.525 63.160 175.780 63.730 ;
        RECT 175.950 63.560 176.880 63.730 ;
        RECT 177.050 64.520 178.060 64.690 ;
        RECT 177.050 63.720 177.220 64.520 ;
        RECT 177.425 64.180 177.700 64.320 ;
        RECT 177.420 64.010 177.700 64.180 ;
        RECT 176.705 63.525 176.880 63.560 ;
        RECT 175.950 62.990 176.280 63.390 ;
        RECT 176.705 63.160 177.235 63.525 ;
        RECT 177.425 63.160 177.700 64.010 ;
        RECT 177.870 63.160 178.060 64.520 ;
        RECT 178.230 64.535 178.400 65.200 ;
        RECT 178.570 64.780 178.740 65.540 ;
        RECT 178.975 64.780 179.490 65.190 ;
        RECT 179.660 65.105 185.005 65.540 ;
        RECT 178.230 64.345 178.980 64.535 ;
        RECT 179.150 63.970 179.490 64.780 ;
        RECT 178.260 63.800 179.490 63.970 ;
        RECT 178.240 62.990 178.750 63.525 ;
        RECT 178.970 63.195 179.215 63.800 ;
        RECT 181.245 63.535 181.585 64.365 ;
        RECT 183.065 63.855 183.415 65.105 ;
        RECT 186.105 64.870 186.360 65.370 ;
        RECT 186.530 65.040 186.860 65.540 ;
        RECT 186.105 64.700 186.855 64.870 ;
        RECT 186.105 63.880 186.455 64.530 ;
        RECT 186.625 63.710 186.855 64.700 ;
        RECT 186.105 63.540 186.855 63.710 ;
        RECT 179.660 62.990 185.005 63.535 ;
        RECT 186.105 63.250 186.360 63.540 ;
        RECT 186.530 62.990 186.860 63.370 ;
        RECT 187.030 63.250 187.200 65.370 ;
        RECT 187.370 64.570 187.695 65.355 ;
        RECT 187.865 65.080 188.115 65.540 ;
        RECT 188.285 65.040 188.535 65.370 ;
        RECT 188.750 65.040 189.430 65.370 ;
        RECT 188.285 64.910 188.455 65.040 ;
        RECT 188.060 64.740 188.455 64.910 ;
        RECT 187.430 63.520 187.890 64.570 ;
        RECT 188.060 63.380 188.230 64.740 ;
        RECT 188.625 64.480 189.090 64.870 ;
        RECT 188.400 63.670 188.750 64.290 ;
        RECT 188.920 63.890 189.090 64.480 ;
        RECT 189.260 64.260 189.430 65.040 ;
        RECT 189.600 64.940 189.770 65.280 ;
        RECT 190.005 65.110 190.335 65.540 ;
        RECT 190.505 64.940 190.675 65.280 ;
        RECT 190.970 65.080 191.340 65.540 ;
        RECT 189.600 64.770 190.675 64.940 ;
        RECT 191.510 64.910 191.680 65.370 ;
        RECT 191.915 65.030 192.785 65.370 ;
        RECT 192.955 65.080 193.205 65.540 ;
        RECT 191.120 64.740 191.680 64.910 ;
        RECT 191.120 64.600 191.290 64.740 ;
        RECT 189.790 64.430 191.290 64.600 ;
        RECT 191.985 64.570 192.445 64.860 ;
        RECT 189.260 64.090 190.950 64.260 ;
        RECT 188.920 63.670 189.275 63.890 ;
        RECT 189.445 63.380 189.615 64.090 ;
        RECT 189.820 63.670 190.610 63.920 ;
        RECT 190.780 63.910 190.950 64.090 ;
        RECT 191.120 63.740 191.290 64.430 ;
        RECT 187.560 62.990 187.890 63.350 ;
        RECT 188.060 63.210 188.555 63.380 ;
        RECT 188.760 63.210 189.615 63.380 ;
        RECT 190.490 62.990 190.820 63.450 ;
        RECT 191.030 63.350 191.290 63.740 ;
        RECT 191.480 64.560 192.445 64.570 ;
        RECT 192.615 64.650 192.785 65.030 ;
        RECT 193.375 64.990 193.545 65.280 ;
        RECT 193.725 65.160 194.055 65.540 ;
        RECT 193.375 64.820 194.175 64.990 ;
        RECT 191.480 64.400 192.155 64.560 ;
        RECT 192.615 64.480 193.835 64.650 ;
        RECT 191.480 63.610 191.690 64.400 ;
        RECT 192.615 64.390 192.785 64.480 ;
        RECT 191.860 63.610 192.210 64.230 ;
        RECT 192.380 64.220 192.785 64.390 ;
        RECT 192.380 63.440 192.550 64.220 ;
        RECT 192.720 63.770 192.940 64.050 ;
        RECT 193.120 63.940 193.660 64.310 ;
        RECT 194.005 64.230 194.175 64.820 ;
        RECT 194.395 64.400 194.700 65.540 ;
        RECT 194.870 64.350 195.120 65.230 ;
        RECT 195.290 64.400 195.540 65.540 ;
        RECT 195.760 64.450 199.270 65.540 ;
        RECT 199.440 64.450 200.650 65.540 ;
        RECT 194.005 64.200 194.745 64.230 ;
        RECT 192.720 63.600 193.250 63.770 ;
        RECT 191.030 63.180 191.380 63.350 ;
        RECT 191.600 63.160 192.550 63.440 ;
        RECT 192.720 62.990 192.910 63.430 ;
        RECT 193.080 63.370 193.250 63.600 ;
        RECT 193.420 63.540 193.660 63.940 ;
        RECT 193.830 63.900 194.745 64.200 ;
        RECT 193.830 63.725 194.155 63.900 ;
        RECT 193.830 63.370 194.150 63.725 ;
        RECT 194.915 63.700 195.120 64.350 ;
        RECT 195.760 63.760 197.410 64.280 ;
        RECT 197.580 63.930 199.270 64.450 ;
        RECT 193.080 63.200 194.150 63.370 ;
        RECT 194.395 62.990 194.700 63.450 ;
        RECT 194.870 63.170 195.120 63.700 ;
        RECT 195.290 62.990 195.540 63.745 ;
        RECT 195.760 62.990 199.270 63.760 ;
        RECT 199.440 63.740 199.960 64.280 ;
        RECT 200.130 63.910 200.650 64.450 ;
        RECT 200.820 64.375 201.110 65.540 ;
        RECT 201.280 64.450 202.950 65.540 ;
        RECT 203.580 65.030 203.840 65.540 ;
        RECT 201.280 63.760 202.030 64.280 ;
        RECT 202.200 63.930 202.950 64.450 ;
        RECT 203.580 63.980 203.920 64.860 ;
        RECT 204.090 64.150 204.260 65.370 ;
        RECT 204.500 65.035 205.115 65.540 ;
        RECT 204.500 64.500 204.750 64.865 ;
        RECT 204.920 64.860 205.115 65.035 ;
        RECT 205.285 65.030 205.760 65.370 ;
        RECT 205.930 64.995 206.145 65.540 ;
        RECT 204.920 64.670 205.250 64.860 ;
        RECT 205.470 64.500 206.185 64.795 ;
        RECT 206.355 64.670 206.630 65.370 ;
        RECT 207.445 65.180 207.895 65.540 ;
        RECT 208.460 65.180 208.790 65.540 ;
        RECT 209.360 65.180 209.695 65.540 ;
        RECT 210.220 65.180 210.550 65.540 ;
        RECT 204.500 64.330 206.290 64.500 ;
        RECT 204.090 63.900 204.885 64.150 ;
        RECT 204.090 63.810 204.340 63.900 ;
        RECT 199.440 62.990 200.650 63.740 ;
        RECT 200.820 62.990 201.110 63.715 ;
        RECT 201.280 62.990 202.950 63.760 ;
        RECT 203.580 62.990 203.840 63.810 ;
        RECT 204.010 63.390 204.340 63.810 ;
        RECT 205.055 63.475 205.310 64.330 ;
        RECT 204.520 63.210 205.310 63.475 ;
        RECT 205.480 63.630 205.890 64.150 ;
        RECT 206.060 63.900 206.290 64.330 ;
        RECT 206.460 63.640 206.630 64.670 ;
        RECT 205.480 63.210 205.680 63.630 ;
        RECT 205.870 62.990 206.200 63.450 ;
        RECT 206.370 63.160 206.630 63.640 ;
        RECT 206.865 64.400 207.225 65.070 ;
        RECT 211.400 65.030 211.660 65.540 ;
        RECT 207.395 64.780 211.160 65.010 ;
        RECT 206.865 63.710 207.085 64.400 ;
        RECT 207.395 64.230 207.565 64.780 ;
        RECT 207.995 64.430 208.770 64.600 ;
        RECT 208.940 64.440 210.250 64.610 ;
        RECT 208.600 64.260 208.770 64.430 ;
        RECT 207.255 63.900 207.565 64.230 ;
        RECT 206.865 63.450 207.350 63.710 ;
        RECT 207.735 63.630 207.950 64.245 ;
        RECT 208.240 63.900 208.430 64.245 ;
        RECT 208.600 63.925 209.815 64.260 ;
        RECT 208.600 63.710 208.830 63.925 ;
        RECT 209.985 63.750 210.250 64.440 ;
        RECT 208.135 63.520 208.830 63.710 ;
        RECT 209.000 63.520 210.250 63.750 ;
        RECT 210.430 63.520 210.710 64.610 ;
        RECT 208.135 63.450 208.315 63.520 ;
        RECT 206.865 63.260 208.315 63.450 ;
        RECT 209.000 63.420 209.190 63.520 ;
        RECT 206.865 63.160 207.350 63.260 ;
        RECT 208.495 62.990 208.825 63.350 ;
        RECT 209.360 62.990 209.690 63.350 ;
        RECT 209.860 63.160 210.050 63.520 ;
        RECT 210.220 62.990 210.550 63.350 ;
        RECT 210.880 63.330 211.160 64.780 ;
        RECT 211.400 63.980 211.740 64.860 ;
        RECT 211.910 64.150 212.080 65.370 ;
        RECT 212.320 65.035 212.935 65.540 ;
        RECT 212.320 64.500 212.570 64.865 ;
        RECT 212.740 64.860 212.935 65.035 ;
        RECT 213.105 65.030 213.580 65.370 ;
        RECT 213.750 64.995 213.965 65.540 ;
        RECT 212.740 64.670 213.070 64.860 ;
        RECT 213.290 64.500 214.005 64.795 ;
        RECT 214.175 64.670 214.450 65.370 ;
        RECT 214.620 65.105 219.965 65.540 ;
        RECT 212.320 64.330 214.110 64.500 ;
        RECT 211.910 63.900 212.705 64.150 ;
        RECT 211.910 63.810 212.160 63.900 ;
        RECT 211.400 62.990 211.660 63.810 ;
        RECT 211.830 63.390 212.160 63.810 ;
        RECT 212.875 63.475 213.130 64.330 ;
        RECT 212.340 63.210 213.130 63.475 ;
        RECT 213.300 63.630 213.710 64.150 ;
        RECT 213.880 63.900 214.110 64.330 ;
        RECT 214.280 63.640 214.450 64.670 ;
        RECT 213.300 63.210 213.500 63.630 ;
        RECT 213.690 62.990 214.020 63.450 ;
        RECT 214.190 63.160 214.450 63.640 ;
        RECT 216.205 63.535 216.545 64.365 ;
        RECT 218.025 63.855 218.375 65.105 ;
        RECT 221.090 64.920 221.420 65.370 ;
        RECT 221.590 65.090 221.760 65.540 ;
        RECT 221.930 64.920 222.260 65.370 ;
        RECT 221.090 64.750 222.260 64.920 ;
        RECT 222.430 65.010 222.680 65.370 ;
        RECT 223.285 65.180 223.615 65.540 ;
        RECT 222.430 64.800 223.540 65.010 ;
        RECT 222.430 64.580 222.600 64.800 ;
        RECT 221.095 63.900 221.385 64.520 ;
        RECT 221.555 63.900 221.970 64.520 ;
        RECT 222.140 64.410 222.600 64.580 ;
        RECT 222.790 64.460 223.200 64.630 ;
        RECT 223.370 64.570 223.540 64.800 ;
        RECT 223.805 64.910 224.060 65.330 ;
        RECT 224.230 65.160 224.565 65.540 ;
        RECT 223.805 64.740 224.505 64.910 ;
        RECT 222.140 63.730 222.310 64.410 ;
        RECT 222.790 64.230 222.960 64.460 ;
        RECT 223.370 64.400 224.085 64.570 ;
        RECT 222.480 63.900 222.960 64.230 ;
        RECT 223.130 63.940 223.585 64.230 ;
        RECT 223.755 63.980 224.085 64.400 ;
        RECT 223.130 63.900 223.325 63.940 ;
        RECT 214.620 62.990 219.965 63.535 ;
        RECT 221.090 62.990 221.420 63.730 ;
        RECT 221.915 63.540 222.310 63.730 ;
        RECT 222.790 63.730 222.960 63.900 ;
        RECT 224.275 63.790 224.505 64.740 ;
        RECT 224.740 64.400 225.000 65.540 ;
        RECT 225.170 64.390 225.500 65.370 ;
        RECT 225.670 64.400 225.950 65.540 ;
        RECT 225.260 64.350 225.435 64.390 ;
        RECT 226.580 64.375 226.870 65.540 ;
        RECT 227.040 65.105 232.385 65.540 ;
        RECT 232.560 65.105 237.905 65.540 ;
        RECT 224.760 63.980 225.095 64.230 ;
        RECT 225.265 63.790 225.435 64.350 ;
        RECT 225.605 63.960 225.940 64.230 ;
        RECT 222.790 63.560 223.200 63.730 ;
        RECT 222.350 62.990 222.680 63.370 ;
        RECT 223.435 62.990 223.635 63.770 ;
        RECT 223.805 63.620 224.505 63.790 ;
        RECT 223.805 63.220 224.135 63.620 ;
        RECT 224.310 62.990 224.565 63.450 ;
        RECT 224.740 63.160 225.435 63.790 ;
        RECT 225.640 62.990 225.950 63.790 ;
        RECT 226.580 62.990 226.870 63.715 ;
        RECT 228.625 63.535 228.965 64.365 ;
        RECT 230.445 63.855 230.795 65.105 ;
        RECT 234.145 63.535 234.485 64.365 ;
        RECT 235.965 63.855 236.315 65.105 ;
        RECT 238.080 64.450 239.750 65.540 ;
        RECT 240.005 64.920 240.180 65.370 ;
        RECT 240.350 65.100 240.680 65.540 ;
        RECT 240.985 64.950 241.155 65.370 ;
        RECT 241.390 65.130 242.060 65.540 ;
        RECT 242.275 64.950 242.445 65.370 ;
        RECT 242.645 65.130 242.975 65.540 ;
        RECT 240.005 64.750 240.635 64.920 ;
        RECT 238.080 63.760 238.830 64.280 ;
        RECT 239.000 63.930 239.750 64.450 ;
        RECT 239.920 63.900 240.285 64.580 ;
        RECT 240.465 64.230 240.635 64.750 ;
        RECT 240.985 64.780 243.000 64.950 ;
        RECT 240.465 63.900 240.815 64.230 ;
        RECT 227.040 62.990 232.385 63.535 ;
        RECT 232.560 62.990 237.905 63.535 ;
        RECT 238.080 62.990 239.750 63.760 ;
        RECT 240.465 63.730 240.635 63.900 ;
        RECT 240.005 63.560 240.635 63.730 ;
        RECT 240.005 63.160 240.180 63.560 ;
        RECT 240.985 63.490 241.155 64.780 ;
        RECT 240.350 62.990 240.680 63.370 ;
        RECT 240.925 63.160 241.155 63.490 ;
        RECT 241.355 63.325 241.635 64.600 ;
        RECT 241.860 63.840 242.130 64.600 ;
        RECT 241.820 63.670 242.130 63.840 ;
        RECT 241.860 63.325 242.130 63.670 ;
        RECT 242.320 63.570 242.660 64.600 ;
        RECT 242.830 64.230 243.000 64.780 ;
        RECT 243.170 64.400 243.430 65.370 ;
        RECT 243.600 65.105 248.945 65.540 ;
        RECT 242.830 63.900 243.090 64.230 ;
        RECT 243.260 63.710 243.430 64.400 ;
        RECT 242.590 62.990 242.920 63.370 ;
        RECT 243.090 63.245 243.430 63.710 ;
        RECT 245.185 63.535 245.525 64.365 ;
        RECT 247.005 63.855 247.355 65.105 ;
        RECT 250.040 65.030 251.230 65.320 ;
        RECT 250.060 64.690 251.230 64.860 ;
        RECT 251.400 64.740 251.680 65.540 ;
        RECT 250.060 64.400 250.385 64.690 ;
        RECT 251.060 64.570 251.230 64.690 ;
        RECT 250.555 64.230 250.750 64.520 ;
        RECT 251.060 64.400 251.720 64.570 ;
        RECT 251.890 64.400 252.165 65.370 ;
        RECT 251.550 64.230 251.720 64.400 ;
        RECT 250.040 63.900 250.385 64.230 ;
        RECT 250.555 63.900 251.380 64.230 ;
        RECT 251.550 63.900 251.825 64.230 ;
        RECT 251.550 63.730 251.720 63.900 ;
        RECT 250.055 63.560 251.720 63.730 ;
        RECT 251.995 63.665 252.165 64.400 ;
        RECT 252.340 64.375 252.630 65.540 ;
        RECT 252.820 64.700 253.075 65.370 ;
        RECT 253.245 64.780 253.575 65.540 ;
        RECT 253.745 64.940 253.995 65.370 ;
        RECT 254.165 65.120 254.520 65.540 ;
        RECT 254.710 65.200 255.880 65.370 ;
        RECT 254.710 65.160 255.040 65.200 ;
        RECT 255.150 64.940 255.380 65.030 ;
        RECT 253.745 64.700 255.380 64.940 ;
        RECT 255.550 64.700 255.880 65.200 ;
        RECT 252.820 64.690 253.030 64.700 ;
        RECT 243.090 63.200 243.425 63.245 ;
        RECT 243.600 62.990 248.945 63.535 ;
        RECT 250.055 63.210 250.310 63.560 ;
        RECT 250.480 62.990 250.810 63.390 ;
        RECT 250.980 63.210 251.150 63.560 ;
        RECT 251.320 62.990 251.700 63.390 ;
        RECT 251.890 63.320 252.165 63.665 ;
        RECT 252.340 62.990 252.630 63.715 ;
        RECT 252.820 63.570 252.990 64.690 ;
        RECT 256.050 64.530 256.220 65.370 ;
        RECT 253.160 64.360 256.220 64.530 ;
        RECT 257.405 64.570 257.740 65.355 ;
        RECT 257.405 64.400 257.990 64.570 ;
        RECT 258.345 64.520 258.600 65.355 ;
        RECT 253.160 63.810 253.330 64.360 ;
        RECT 253.560 63.980 253.925 64.180 ;
        RECT 254.095 63.980 254.425 64.180 ;
        RECT 253.160 63.640 253.960 63.810 ;
        RECT 252.820 63.490 253.005 63.570 ;
        RECT 252.820 63.160 253.075 63.490 ;
        RECT 253.290 62.990 253.620 63.470 ;
        RECT 253.790 63.410 253.960 63.640 ;
        RECT 254.140 63.580 254.425 63.980 ;
        RECT 254.695 63.980 255.170 64.180 ;
        RECT 255.340 63.980 255.785 64.180 ;
        RECT 255.955 63.980 256.305 64.190 ;
        RECT 254.695 63.580 254.975 63.980 ;
        RECT 255.155 63.640 256.220 63.810 ;
        RECT 257.400 63.650 257.650 64.230 ;
        RECT 257.820 63.730 257.990 64.400 ;
        RECT 258.160 64.320 258.600 64.520 ;
        RECT 258.160 63.900 258.390 64.320 ;
        RECT 258.770 64.150 259.010 65.355 ;
        RECT 259.270 64.740 259.530 65.540 ;
        RECT 259.700 65.105 265.045 65.540 ;
        RECT 258.560 63.980 259.010 64.150 ;
        RECT 255.155 63.410 255.325 63.640 ;
        RECT 253.790 63.160 255.325 63.410 ;
        RECT 255.550 62.990 255.880 63.470 ;
        RECT 256.050 63.160 256.220 63.640 ;
        RECT 257.820 63.560 259.020 63.730 ;
        RECT 259.270 63.560 259.530 64.570 ;
        RECT 257.820 63.550 258.175 63.560 ;
        RECT 257.400 62.990 257.660 63.480 ;
        RECT 257.910 63.290 258.175 63.550 ;
        RECT 258.350 62.990 258.680 63.390 ;
        RECT 258.850 63.290 259.020 63.560 ;
        RECT 261.285 63.535 261.625 64.365 ;
        RECT 263.105 63.855 263.455 65.105 ;
        RECT 265.220 64.450 266.890 65.540 ;
        RECT 265.220 63.760 265.970 64.280 ;
        RECT 266.140 63.930 266.890 64.450 ;
        RECT 267.150 64.610 267.320 65.370 ;
        RECT 267.500 64.780 267.830 65.540 ;
        RECT 267.150 64.440 267.815 64.610 ;
        RECT 268.000 64.465 268.270 65.370 ;
        RECT 267.645 64.295 267.815 64.440 ;
        RECT 267.080 63.890 267.410 64.260 ;
        RECT 267.645 63.965 267.930 64.295 ;
        RECT 259.190 62.990 259.520 63.390 ;
        RECT 259.700 62.990 265.045 63.535 ;
        RECT 265.220 62.990 266.890 63.760 ;
        RECT 267.645 63.710 267.815 63.965 ;
        RECT 267.150 63.540 267.815 63.710 ;
        RECT 268.100 63.665 268.270 64.465 ;
        RECT 268.490 64.400 268.740 65.540 ;
        RECT 268.910 64.350 269.160 65.230 ;
        RECT 269.330 64.400 269.635 65.540 ;
        RECT 269.975 65.160 270.305 65.540 ;
        RECT 270.485 64.990 270.655 65.280 ;
        RECT 270.825 65.080 271.075 65.540 ;
        RECT 269.855 64.820 270.655 64.990 ;
        RECT 271.245 65.030 272.115 65.370 ;
        RECT 267.150 63.160 267.320 63.540 ;
        RECT 267.500 62.990 267.830 63.370 ;
        RECT 268.010 63.160 268.270 63.665 ;
        RECT 268.490 62.990 268.740 63.745 ;
        RECT 268.910 63.700 269.115 64.350 ;
        RECT 269.855 64.230 270.025 64.820 ;
        RECT 271.245 64.650 271.415 65.030 ;
        RECT 272.350 64.910 272.520 65.370 ;
        RECT 272.690 65.080 273.060 65.540 ;
        RECT 273.355 64.940 273.525 65.280 ;
        RECT 273.695 65.110 274.025 65.540 ;
        RECT 274.260 64.940 274.430 65.280 ;
        RECT 270.195 64.480 271.415 64.650 ;
        RECT 271.585 64.570 272.045 64.860 ;
        RECT 272.350 64.740 272.910 64.910 ;
        RECT 273.355 64.770 274.430 64.940 ;
        RECT 274.600 65.040 275.280 65.370 ;
        RECT 275.495 65.040 275.745 65.370 ;
        RECT 275.915 65.080 276.165 65.540 ;
        RECT 272.740 64.600 272.910 64.740 ;
        RECT 271.585 64.560 272.550 64.570 ;
        RECT 271.245 64.390 271.415 64.480 ;
        RECT 271.875 64.400 272.550 64.560 ;
        RECT 269.285 64.200 270.025 64.230 ;
        RECT 269.285 63.900 270.200 64.200 ;
        RECT 269.875 63.725 270.200 63.900 ;
        RECT 268.910 63.170 269.160 63.700 ;
        RECT 269.330 62.990 269.635 63.450 ;
        RECT 269.880 63.370 270.200 63.725 ;
        RECT 270.370 63.940 270.910 64.310 ;
        RECT 271.245 64.220 271.650 64.390 ;
        RECT 270.370 63.540 270.610 63.940 ;
        RECT 271.090 63.770 271.310 64.050 ;
        RECT 270.780 63.600 271.310 63.770 ;
        RECT 270.780 63.370 270.950 63.600 ;
        RECT 271.480 63.440 271.650 64.220 ;
        RECT 271.820 63.610 272.170 64.230 ;
        RECT 272.340 63.610 272.550 64.400 ;
        RECT 272.740 64.430 274.240 64.600 ;
        RECT 272.740 63.740 272.910 64.430 ;
        RECT 274.600 64.260 274.770 65.040 ;
        RECT 275.575 64.910 275.745 65.040 ;
        RECT 273.080 64.090 274.770 64.260 ;
        RECT 274.940 64.480 275.405 64.870 ;
        RECT 275.575 64.740 275.970 64.910 ;
        RECT 273.080 63.910 273.250 64.090 ;
        RECT 269.880 63.200 270.950 63.370 ;
        RECT 271.120 62.990 271.310 63.430 ;
        RECT 271.480 63.160 272.430 63.440 ;
        RECT 272.740 63.350 273.000 63.740 ;
        RECT 273.420 63.670 274.210 63.920 ;
        RECT 272.650 63.180 273.000 63.350 ;
        RECT 273.210 62.990 273.540 63.450 ;
        RECT 274.415 63.380 274.585 64.090 ;
        RECT 274.940 63.890 275.110 64.480 ;
        RECT 274.755 63.670 275.110 63.890 ;
        RECT 275.280 63.670 275.630 64.290 ;
        RECT 275.800 63.380 275.970 64.740 ;
        RECT 276.335 64.570 276.660 65.355 ;
        RECT 276.140 63.520 276.600 64.570 ;
        RECT 274.415 63.210 275.270 63.380 ;
        RECT 275.475 63.210 275.970 63.380 ;
        RECT 276.140 62.990 276.470 63.350 ;
        RECT 276.830 63.250 277.000 65.370 ;
        RECT 277.170 65.040 277.500 65.540 ;
        RECT 277.670 64.870 277.925 65.370 ;
        RECT 277.175 64.700 277.925 64.870 ;
        RECT 277.175 63.710 277.405 64.700 ;
        RECT 277.575 63.880 277.925 64.530 ;
        RECT 278.100 64.375 278.390 65.540 ;
        RECT 278.560 65.105 283.905 65.540 ;
        RECT 284.080 65.105 289.425 65.540 ;
        RECT 277.175 63.540 277.925 63.710 ;
        RECT 277.170 62.990 277.500 63.370 ;
        RECT 277.670 63.250 277.925 63.540 ;
        RECT 278.100 62.990 278.390 63.715 ;
        RECT 280.145 63.535 280.485 64.365 ;
        RECT 281.965 63.855 282.315 65.105 ;
        RECT 285.665 63.535 286.005 64.365 ;
        RECT 287.485 63.855 287.835 65.105 ;
        RECT 290.520 64.780 291.035 65.190 ;
        RECT 291.270 64.780 291.440 65.540 ;
        RECT 291.610 65.200 293.640 65.370 ;
        RECT 290.520 63.970 290.860 64.780 ;
        RECT 291.610 64.535 291.780 65.200 ;
        RECT 292.175 64.860 293.300 65.030 ;
        RECT 291.030 64.345 291.780 64.535 ;
        RECT 291.950 64.520 292.960 64.690 ;
        RECT 290.520 63.800 291.750 63.970 ;
        RECT 278.560 62.990 283.905 63.535 ;
        RECT 284.080 62.990 289.425 63.535 ;
        RECT 290.795 63.195 291.040 63.800 ;
        RECT 291.260 62.990 291.770 63.525 ;
        RECT 291.950 63.160 292.140 64.520 ;
        RECT 292.310 64.180 292.585 64.320 ;
        RECT 292.310 64.010 292.590 64.180 ;
        RECT 292.310 63.160 292.585 64.010 ;
        RECT 292.790 63.720 292.960 64.520 ;
        RECT 293.130 63.730 293.300 64.860 ;
        RECT 293.470 64.230 293.640 65.200 ;
        RECT 293.810 64.400 293.980 65.540 ;
        RECT 294.150 64.400 294.485 65.370 ;
        RECT 293.470 63.900 293.665 64.230 ;
        RECT 293.890 63.900 294.145 64.230 ;
        RECT 293.890 63.730 294.060 63.900 ;
        RECT 294.315 63.730 294.485 64.400 ;
        RECT 295.580 64.780 296.095 65.190 ;
        RECT 296.330 64.780 296.500 65.540 ;
        RECT 296.670 65.200 298.700 65.370 ;
        RECT 295.580 63.970 295.920 64.780 ;
        RECT 296.670 64.535 296.840 65.200 ;
        RECT 297.235 64.860 298.360 65.030 ;
        RECT 296.090 64.345 296.840 64.535 ;
        RECT 297.010 64.520 298.020 64.690 ;
        RECT 295.580 63.800 296.810 63.970 ;
        RECT 293.130 63.560 294.060 63.730 ;
        RECT 293.130 63.525 293.305 63.560 ;
        RECT 292.775 63.160 293.305 63.525 ;
        RECT 293.730 62.990 294.060 63.390 ;
        RECT 294.230 63.160 294.485 63.730 ;
        RECT 295.855 63.195 296.100 63.800 ;
        RECT 296.320 62.990 296.830 63.525 ;
        RECT 297.010 63.160 297.200 64.520 ;
        RECT 297.370 63.500 297.645 64.320 ;
        RECT 297.850 63.720 298.020 64.520 ;
        RECT 298.190 63.730 298.360 64.860 ;
        RECT 298.530 64.230 298.700 65.200 ;
        RECT 298.870 64.400 299.040 65.540 ;
        RECT 299.210 64.400 299.545 65.370 ;
        RECT 299.720 64.450 303.230 65.540 ;
        RECT 298.530 63.900 298.725 64.230 ;
        RECT 298.950 63.900 299.205 64.230 ;
        RECT 298.950 63.730 299.120 63.900 ;
        RECT 299.375 63.730 299.545 64.400 ;
        RECT 298.190 63.560 299.120 63.730 ;
        RECT 298.190 63.525 298.365 63.560 ;
        RECT 297.370 63.330 297.650 63.500 ;
        RECT 297.370 63.160 297.645 63.330 ;
        RECT 297.835 63.160 298.365 63.525 ;
        RECT 298.790 62.990 299.120 63.390 ;
        RECT 299.290 63.160 299.545 63.730 ;
        RECT 299.720 63.760 301.370 64.280 ;
        RECT 301.540 63.930 303.230 64.450 ;
        RECT 303.860 64.375 304.150 65.540 ;
        RECT 304.320 65.105 309.665 65.540 ;
        RECT 299.720 62.990 303.230 63.760 ;
        RECT 303.860 62.990 304.150 63.715 ;
        RECT 305.905 63.535 306.245 64.365 ;
        RECT 307.725 63.855 308.075 65.105 ;
        RECT 309.840 64.450 311.050 65.540 ;
        RECT 309.840 63.910 310.360 64.450 ;
        RECT 310.530 63.740 311.050 64.280 ;
        RECT 304.320 62.990 309.665 63.535 ;
        RECT 309.840 62.990 311.050 63.740 ;
        RECT 162.095 62.820 311.135 62.990 ;
        RECT 162.180 62.070 163.390 62.820 ;
        RECT 162.180 61.530 162.700 62.070 ;
        RECT 163.565 61.980 163.825 62.820 ;
        RECT 164.000 62.075 164.255 62.650 ;
        RECT 164.425 62.440 164.755 62.820 ;
        RECT 164.970 62.270 165.140 62.650 ;
        RECT 164.425 62.100 165.140 62.270 ;
        RECT 162.870 61.360 163.390 61.900 ;
        RECT 162.180 60.270 163.390 61.360 ;
        RECT 163.565 60.270 163.825 61.420 ;
        RECT 164.000 61.345 164.170 62.075 ;
        RECT 164.425 61.910 164.595 62.100 ;
        RECT 165.400 62.050 167.990 62.820 ;
        RECT 168.620 62.145 168.880 62.650 ;
        RECT 169.060 62.440 169.390 62.820 ;
        RECT 169.570 62.270 169.740 62.650 ;
        RECT 164.340 61.580 164.595 61.910 ;
        RECT 164.425 61.370 164.595 61.580 ;
        RECT 164.875 61.550 165.230 61.920 ;
        RECT 165.400 61.530 166.610 62.050 ;
        RECT 164.000 60.440 164.255 61.345 ;
        RECT 164.425 61.200 165.140 61.370 ;
        RECT 166.780 61.360 167.990 61.880 ;
        RECT 164.425 60.270 164.755 61.030 ;
        RECT 164.970 60.440 165.140 61.200 ;
        RECT 165.400 60.270 167.990 61.360 ;
        RECT 168.620 61.345 168.790 62.145 ;
        RECT 169.075 62.100 169.740 62.270 ;
        RECT 169.075 61.845 169.245 62.100 ;
        RECT 170.000 62.050 171.670 62.820 ;
        RECT 172.305 62.080 172.560 62.650 ;
        RECT 172.730 62.420 173.060 62.820 ;
        RECT 173.485 62.285 174.015 62.650 ;
        RECT 174.205 62.480 174.480 62.650 ;
        RECT 174.200 62.310 174.480 62.480 ;
        RECT 173.485 62.250 173.660 62.285 ;
        RECT 172.730 62.080 173.660 62.250 ;
        RECT 168.960 61.515 169.245 61.845 ;
        RECT 169.480 61.550 169.810 61.920 ;
        RECT 170.000 61.530 170.750 62.050 ;
        RECT 169.075 61.370 169.245 61.515 ;
        RECT 168.620 60.440 168.890 61.345 ;
        RECT 169.075 61.200 169.740 61.370 ;
        RECT 170.920 61.360 171.670 61.880 ;
        RECT 169.060 60.270 169.390 61.030 ;
        RECT 169.570 60.440 169.740 61.200 ;
        RECT 170.000 60.270 171.670 61.360 ;
        RECT 172.305 61.410 172.475 62.080 ;
        RECT 172.730 61.910 172.900 62.080 ;
        RECT 172.645 61.580 172.900 61.910 ;
        RECT 173.125 61.580 173.320 61.910 ;
        RECT 172.305 60.440 172.640 61.410 ;
        RECT 172.810 60.270 172.980 61.410 ;
        RECT 173.150 60.610 173.320 61.580 ;
        RECT 173.490 60.950 173.660 62.080 ;
        RECT 173.830 61.290 174.000 62.090 ;
        RECT 174.205 61.490 174.480 62.310 ;
        RECT 174.650 61.290 174.840 62.650 ;
        RECT 175.020 62.285 175.530 62.820 ;
        RECT 175.750 62.010 175.995 62.615 ;
        RECT 176.445 62.080 176.700 62.650 ;
        RECT 176.870 62.420 177.200 62.820 ;
        RECT 177.625 62.285 178.155 62.650 ;
        RECT 178.345 62.480 178.620 62.650 ;
        RECT 178.340 62.310 178.620 62.480 ;
        RECT 177.625 62.250 177.800 62.285 ;
        RECT 176.870 62.080 177.800 62.250 ;
        RECT 175.040 61.840 176.270 62.010 ;
        RECT 173.830 61.120 174.840 61.290 ;
        RECT 175.010 61.275 175.760 61.465 ;
        RECT 173.490 60.780 174.615 60.950 ;
        RECT 175.010 60.610 175.180 61.275 ;
        RECT 175.930 61.030 176.270 61.840 ;
        RECT 173.150 60.440 175.180 60.610 ;
        RECT 175.350 60.270 175.520 61.030 ;
        RECT 175.755 60.620 176.270 61.030 ;
        RECT 176.445 61.410 176.615 62.080 ;
        RECT 176.870 61.910 177.040 62.080 ;
        RECT 176.785 61.580 177.040 61.910 ;
        RECT 177.265 61.580 177.460 61.910 ;
        RECT 176.445 60.440 176.780 61.410 ;
        RECT 176.950 60.270 177.120 61.410 ;
        RECT 177.290 60.610 177.460 61.580 ;
        RECT 177.630 60.950 177.800 62.080 ;
        RECT 177.970 61.290 178.140 62.090 ;
        RECT 178.345 61.490 178.620 62.310 ;
        RECT 178.790 61.290 178.980 62.650 ;
        RECT 179.160 62.285 179.670 62.820 ;
        RECT 179.890 62.010 180.135 62.615 ;
        RECT 180.580 62.275 185.925 62.820 ;
        RECT 179.180 61.840 180.410 62.010 ;
        RECT 177.970 61.120 178.980 61.290 ;
        RECT 179.150 61.275 179.900 61.465 ;
        RECT 177.630 60.780 178.755 60.950 ;
        RECT 179.150 60.610 179.320 61.275 ;
        RECT 180.070 61.030 180.410 61.840 ;
        RECT 182.165 61.445 182.505 62.275 ;
        RECT 186.100 62.050 187.770 62.820 ;
        RECT 187.940 62.095 188.230 62.820 ;
        RECT 188.400 62.050 191.910 62.820 ;
        RECT 192.080 62.145 192.340 62.650 ;
        RECT 192.520 62.440 192.850 62.820 ;
        RECT 193.030 62.270 193.200 62.650 ;
        RECT 193.460 62.275 198.805 62.820 ;
        RECT 177.290 60.440 179.320 60.610 ;
        RECT 179.490 60.270 179.660 61.030 ;
        RECT 179.895 60.620 180.410 61.030 ;
        RECT 183.985 60.705 184.335 61.955 ;
        RECT 186.100 61.530 186.850 62.050 ;
        RECT 187.020 61.360 187.770 61.880 ;
        RECT 188.400 61.530 190.050 62.050 ;
        RECT 180.580 60.270 185.925 60.705 ;
        RECT 186.100 60.270 187.770 61.360 ;
        RECT 187.940 60.270 188.230 61.435 ;
        RECT 190.220 61.360 191.910 61.880 ;
        RECT 188.400 60.270 191.910 61.360 ;
        RECT 192.080 61.345 192.250 62.145 ;
        RECT 192.535 62.100 193.200 62.270 ;
        RECT 192.535 61.845 192.705 62.100 ;
        RECT 192.420 61.515 192.705 61.845 ;
        RECT 192.940 61.550 193.270 61.920 ;
        RECT 192.535 61.370 192.705 61.515 ;
        RECT 195.045 61.445 195.385 62.275 ;
        RECT 198.980 62.050 202.490 62.820 ;
        RECT 202.670 62.480 203.860 62.650 ;
        RECT 202.670 62.310 202.980 62.480 ;
        RECT 192.080 60.440 192.350 61.345 ;
        RECT 192.535 61.200 193.200 61.370 ;
        RECT 192.520 60.270 192.850 61.030 ;
        RECT 193.030 60.440 193.200 61.200 ;
        RECT 196.865 60.705 197.215 61.955 ;
        RECT 198.980 61.530 200.630 62.050 ;
        RECT 200.800 61.360 202.490 61.880 ;
        RECT 202.665 61.505 202.980 62.140 ;
        RECT 193.460 60.270 198.805 60.705 ;
        RECT 198.980 60.270 202.490 61.360 ;
        RECT 202.670 60.270 202.980 61.335 ;
        RECT 203.150 61.120 203.360 62.310 ;
        RECT 203.530 62.190 203.860 62.480 ;
        RECT 204.100 62.360 204.270 62.820 ;
        RECT 204.500 62.190 204.830 62.650 ;
        RECT 205.010 62.360 205.180 62.820 ;
        RECT 205.360 62.190 205.690 62.650 ;
        RECT 203.530 62.020 205.690 62.190 ;
        RECT 205.880 62.050 207.550 62.820 ;
        RECT 207.740 62.335 208.530 62.600 ;
        RECT 203.700 61.460 204.195 61.830 ;
        RECT 204.375 61.630 205.175 61.830 ;
        RECT 205.345 61.460 205.675 61.850 ;
        RECT 205.880 61.530 206.630 62.050 ;
        RECT 203.640 61.290 205.675 61.460 ;
        RECT 206.800 61.360 207.550 61.880 ;
        RECT 207.720 61.660 208.105 62.140 ;
        RECT 208.275 61.480 208.530 62.335 ;
        RECT 208.700 62.155 208.930 62.600 ;
        RECT 209.110 62.325 209.440 62.820 ;
        RECT 209.615 62.190 209.865 62.650 ;
        RECT 208.700 61.660 209.110 62.155 ;
        RECT 209.695 61.980 209.865 62.190 ;
        RECT 210.035 62.160 210.310 62.820 ;
        RECT 210.480 62.320 210.780 62.650 ;
        RECT 210.950 62.340 211.225 62.820 ;
        RECT 209.295 61.480 209.525 61.910 ;
        RECT 203.150 60.940 204.800 61.120 ;
        RECT 203.150 60.440 203.385 60.940 ;
        RECT 204.500 60.780 204.800 60.940 ;
        RECT 203.555 60.270 203.885 60.730 ;
        RECT 204.080 60.610 204.270 60.770 ;
        RECT 204.970 60.610 205.190 61.120 ;
        RECT 204.080 60.440 205.190 60.610 ;
        RECT 205.360 60.270 205.690 61.120 ;
        RECT 205.880 60.270 207.550 61.360 ;
        RECT 207.735 61.310 209.525 61.480 ;
        RECT 209.695 61.460 210.310 61.980 ;
        RECT 207.735 60.945 207.990 61.310 ;
        RECT 208.160 60.950 208.490 61.140 ;
        RECT 208.715 61.015 208.965 61.310 ;
        RECT 208.160 60.775 208.350 60.950 ;
        RECT 207.720 60.270 208.350 60.775 ;
        RECT 208.530 60.440 209.005 60.780 ;
        RECT 209.190 60.270 209.405 61.115 ;
        RECT 209.710 61.110 209.880 61.460 ;
        RECT 210.480 61.410 210.650 62.320 ;
        RECT 211.405 62.170 211.700 62.560 ;
        RECT 211.870 62.340 212.125 62.820 ;
        RECT 212.300 62.170 212.560 62.560 ;
        RECT 212.730 62.340 213.010 62.820 ;
        RECT 210.820 61.580 211.170 62.150 ;
        RECT 211.405 62.000 213.055 62.170 ;
        RECT 213.700 62.095 213.990 62.820 ;
        RECT 214.360 62.190 214.690 62.550 ;
        RECT 215.320 62.360 215.570 62.820 ;
        RECT 215.740 62.360 216.290 62.650 ;
        RECT 214.360 62.000 215.750 62.190 ;
        RECT 211.340 61.660 212.480 61.830 ;
        RECT 211.340 61.410 211.510 61.660 ;
        RECT 212.650 61.490 213.055 62.000 ;
        RECT 215.580 61.910 215.750 62.000 ;
        RECT 209.605 60.440 209.880 61.110 ;
        RECT 210.050 60.270 210.310 61.280 ;
        RECT 210.480 61.240 211.510 61.410 ;
        RECT 212.300 61.320 213.055 61.490 ;
        RECT 214.160 61.580 214.850 61.830 ;
        RECT 215.080 61.580 215.410 61.830 ;
        RECT 215.580 61.580 215.870 61.910 ;
        RECT 210.480 60.440 210.790 61.240 ;
        RECT 212.300 61.070 212.560 61.320 ;
        RECT 210.960 60.270 211.270 61.070 ;
        RECT 211.440 60.900 212.560 61.070 ;
        RECT 211.440 60.440 211.700 60.900 ;
        RECT 211.870 60.270 212.125 60.730 ;
        RECT 212.300 60.440 212.560 60.900 ;
        RECT 212.730 60.270 213.015 61.140 ;
        RECT 213.700 60.270 213.990 61.435 ;
        RECT 214.160 61.140 214.475 61.580 ;
        RECT 215.580 61.330 215.750 61.580 ;
        RECT 214.810 61.160 215.750 61.330 ;
        RECT 214.360 60.270 214.640 60.940 ;
        RECT 214.810 60.610 215.110 61.160 ;
        RECT 216.040 60.990 216.290 62.360 ;
        RECT 216.460 62.020 216.750 62.820 ;
        RECT 217.120 62.190 217.450 62.550 ;
        RECT 218.080 62.360 218.330 62.820 ;
        RECT 218.500 62.360 219.050 62.650 ;
        RECT 217.120 62.000 218.510 62.190 ;
        RECT 218.340 61.910 218.510 62.000 ;
        RECT 216.920 61.580 217.610 61.830 ;
        RECT 217.840 61.580 218.170 61.830 ;
        RECT 218.340 61.580 218.630 61.910 ;
        RECT 215.320 60.270 215.650 60.990 ;
        RECT 215.840 60.440 216.290 60.990 ;
        RECT 216.460 60.270 216.750 61.410 ;
        RECT 216.920 61.140 217.235 61.580 ;
        RECT 218.340 61.330 218.510 61.580 ;
        RECT 217.570 61.160 218.510 61.330 ;
        RECT 217.120 60.270 217.400 60.940 ;
        RECT 217.570 60.610 217.870 61.160 ;
        RECT 218.800 60.990 219.050 62.360 ;
        RECT 219.220 62.020 219.510 62.820 ;
        RECT 219.880 62.190 220.210 62.550 ;
        RECT 220.840 62.360 221.090 62.820 ;
        RECT 221.260 62.360 221.810 62.650 ;
        RECT 219.880 62.000 221.270 62.190 ;
        RECT 221.100 61.910 221.270 62.000 ;
        RECT 219.680 61.580 220.370 61.830 ;
        RECT 220.600 61.580 220.930 61.830 ;
        RECT 221.100 61.580 221.390 61.910 ;
        RECT 218.080 60.270 218.410 60.990 ;
        RECT 218.600 60.440 219.050 60.990 ;
        RECT 219.220 60.270 219.510 61.410 ;
        RECT 219.680 61.140 219.995 61.580 ;
        RECT 221.100 61.330 221.270 61.580 ;
        RECT 220.330 61.160 221.270 61.330 ;
        RECT 219.880 60.270 220.160 60.940 ;
        RECT 220.330 60.610 220.630 61.160 ;
        RECT 221.560 60.990 221.810 62.360 ;
        RECT 221.980 62.020 222.270 62.820 ;
        RECT 222.440 62.275 227.785 62.820 ;
        RECT 229.045 62.310 229.285 62.820 ;
        RECT 229.465 62.310 229.745 62.640 ;
        RECT 229.975 62.310 230.190 62.820 ;
        RECT 224.025 61.445 224.365 62.275 ;
        RECT 220.840 60.270 221.170 60.990 ;
        RECT 221.360 60.440 221.810 60.990 ;
        RECT 221.980 60.270 222.270 61.410 ;
        RECT 225.845 60.705 226.195 61.955 ;
        RECT 228.940 61.580 229.295 62.140 ;
        RECT 229.465 61.410 229.635 62.310 ;
        RECT 229.805 61.580 230.070 62.140 ;
        RECT 230.360 62.080 230.975 62.650 ;
        RECT 230.320 61.410 230.490 61.910 ;
        RECT 229.065 61.240 230.490 61.410 ;
        RECT 229.065 61.065 229.455 61.240 ;
        RECT 222.440 60.270 227.785 60.705 ;
        RECT 229.940 60.270 230.270 61.070 ;
        RECT 230.660 61.060 230.975 62.080 ;
        RECT 231.385 62.040 231.885 62.650 ;
        RECT 231.180 61.580 231.530 61.830 ;
        RECT 231.715 61.410 231.885 62.040 ;
        RECT 232.515 62.170 232.845 62.650 ;
        RECT 233.015 62.360 233.240 62.820 ;
        RECT 233.410 62.170 233.740 62.650 ;
        RECT 232.515 62.000 233.740 62.170 ;
        RECT 233.930 62.020 234.180 62.820 ;
        RECT 234.350 62.020 234.690 62.650 ;
        RECT 232.055 61.630 232.385 61.830 ;
        RECT 232.555 61.630 232.885 61.830 ;
        RECT 233.055 61.630 233.475 61.830 ;
        RECT 233.650 61.660 234.345 61.830 ;
        RECT 233.650 61.410 233.820 61.660 ;
        RECT 234.515 61.410 234.690 62.020 ;
        RECT 230.440 60.440 230.975 61.060 ;
        RECT 231.385 61.240 233.820 61.410 ;
        RECT 231.385 60.440 231.715 61.240 ;
        RECT 231.885 60.270 232.215 61.070 ;
        RECT 232.515 60.440 232.845 61.240 ;
        RECT 233.490 60.270 233.740 61.070 ;
        RECT 234.010 60.270 234.180 61.410 ;
        RECT 234.350 60.440 234.690 61.410 ;
        RECT 234.870 62.095 235.200 62.605 ;
        RECT 235.370 62.420 235.700 62.820 ;
        RECT 236.750 62.250 237.080 62.590 ;
        RECT 237.250 62.420 237.580 62.820 ;
        RECT 234.870 61.330 235.060 62.095 ;
        RECT 235.370 62.080 237.735 62.250 ;
        RECT 235.370 61.910 235.540 62.080 ;
        RECT 235.230 61.580 235.540 61.910 ;
        RECT 235.710 61.580 236.015 61.910 ;
        RECT 234.870 60.480 235.200 61.330 ;
        RECT 235.370 60.270 235.620 61.410 ;
        RECT 235.800 61.250 236.015 61.580 ;
        RECT 236.190 61.250 236.475 61.910 ;
        RECT 236.670 61.250 236.935 61.910 ;
        RECT 237.150 61.250 237.395 61.910 ;
        RECT 237.565 61.080 237.735 62.080 ;
        RECT 238.080 62.070 239.290 62.820 ;
        RECT 239.460 62.095 239.750 62.820 ;
        RECT 239.920 62.275 245.265 62.820 ;
        RECT 245.440 62.275 250.785 62.820 ;
        RECT 238.080 61.530 238.600 62.070 ;
        RECT 238.770 61.360 239.290 61.900 ;
        RECT 241.505 61.445 241.845 62.275 ;
        RECT 235.810 60.910 237.100 61.080 ;
        RECT 235.810 60.490 236.060 60.910 ;
        RECT 236.290 60.270 236.620 60.740 ;
        RECT 236.850 60.490 237.100 60.910 ;
        RECT 237.280 60.910 237.735 61.080 ;
        RECT 237.280 60.480 237.610 60.910 ;
        RECT 238.080 60.270 239.290 61.360 ;
        RECT 239.460 60.270 239.750 61.435 ;
        RECT 243.325 60.705 243.675 61.955 ;
        RECT 247.025 61.445 247.365 62.275 ;
        RECT 250.960 62.070 252.170 62.820 ;
        RECT 252.340 62.190 252.680 62.650 ;
        RECT 252.850 62.360 253.020 62.820 ;
        RECT 253.650 62.385 254.010 62.650 ;
        RECT 253.655 62.380 254.010 62.385 ;
        RECT 253.660 62.370 254.010 62.380 ;
        RECT 253.665 62.365 254.010 62.370 ;
        RECT 253.670 62.355 254.010 62.365 ;
        RECT 254.250 62.360 254.420 62.820 ;
        RECT 253.675 62.350 254.010 62.355 ;
        RECT 253.685 62.340 254.010 62.350 ;
        RECT 253.695 62.330 254.010 62.340 ;
        RECT 253.190 62.190 253.520 62.270 ;
        RECT 248.845 60.705 249.195 61.955 ;
        RECT 250.960 61.530 251.480 62.070 ;
        RECT 252.340 62.000 253.520 62.190 ;
        RECT 253.710 62.190 254.010 62.330 ;
        RECT 253.710 62.000 254.420 62.190 ;
        RECT 251.650 61.360 252.170 61.900 ;
        RECT 239.920 60.270 245.265 60.705 ;
        RECT 245.440 60.270 250.785 60.705 ;
        RECT 250.960 60.270 252.170 61.360 ;
        RECT 252.340 61.630 252.670 61.830 ;
        RECT 252.980 61.810 253.310 61.830 ;
        RECT 252.860 61.630 253.310 61.810 ;
        RECT 252.340 61.290 252.570 61.630 ;
        RECT 252.350 60.270 252.680 60.990 ;
        RECT 252.860 60.515 253.075 61.630 ;
        RECT 253.480 61.600 253.950 61.830 ;
        RECT 254.135 61.430 254.420 62.000 ;
        RECT 254.590 61.875 254.930 62.650 ;
        RECT 253.270 61.215 254.420 61.430 ;
        RECT 253.270 60.440 253.600 61.215 ;
        RECT 253.770 60.270 254.480 61.045 ;
        RECT 254.650 60.440 254.930 61.875 ;
        RECT 255.100 62.050 256.770 62.820 ;
        RECT 256.950 62.090 257.250 62.820 ;
        RECT 255.100 61.530 255.850 62.050 ;
        RECT 257.430 61.910 257.660 62.530 ;
        RECT 257.860 62.260 258.085 62.640 ;
        RECT 258.255 62.430 258.585 62.820 ;
        RECT 258.780 62.275 264.125 62.820 ;
        RECT 257.860 62.080 258.190 62.260 ;
        RECT 256.020 61.360 256.770 61.880 ;
        RECT 256.955 61.580 257.250 61.910 ;
        RECT 257.430 61.580 257.845 61.910 ;
        RECT 258.015 61.410 258.190 62.080 ;
        RECT 258.360 61.580 258.600 62.230 ;
        RECT 260.365 61.445 260.705 62.275 ;
        RECT 265.220 62.095 265.510 62.820 ;
        RECT 265.680 62.050 267.350 62.820 ;
        RECT 267.520 62.080 267.905 62.650 ;
        RECT 268.075 62.360 268.400 62.820 ;
        RECT 268.920 62.190 269.200 62.650 ;
        RECT 255.100 60.270 256.770 61.360 ;
        RECT 256.950 61.050 257.845 61.380 ;
        RECT 258.015 61.220 258.600 61.410 ;
        RECT 256.950 60.880 258.155 61.050 ;
        RECT 256.950 60.450 257.280 60.880 ;
        RECT 257.460 60.270 257.655 60.710 ;
        RECT 257.825 60.450 258.155 60.880 ;
        RECT 258.325 60.450 258.600 61.220 ;
        RECT 262.185 60.705 262.535 61.955 ;
        RECT 265.680 61.530 266.430 62.050 ;
        RECT 258.780 60.270 264.125 60.705 ;
        RECT 265.220 60.270 265.510 61.435 ;
        RECT 266.600 61.360 267.350 61.880 ;
        RECT 265.680 60.270 267.350 61.360 ;
        RECT 267.520 61.410 267.800 62.080 ;
        RECT 268.075 62.020 269.200 62.190 ;
        RECT 268.075 61.910 268.525 62.020 ;
        RECT 267.970 61.580 268.525 61.910 ;
        RECT 269.390 61.850 269.790 62.650 ;
        RECT 270.190 62.360 270.460 62.820 ;
        RECT 270.630 62.190 270.915 62.650 ;
        RECT 267.520 60.440 267.905 61.410 ;
        RECT 268.075 61.120 268.525 61.580 ;
        RECT 268.695 61.290 269.790 61.850 ;
        RECT 268.075 60.900 269.200 61.120 ;
        RECT 268.075 60.270 268.400 60.730 ;
        RECT 268.920 60.440 269.200 60.900 ;
        RECT 269.390 60.440 269.790 61.290 ;
        RECT 269.960 62.020 270.915 62.190 ;
        RECT 271.200 62.070 272.410 62.820 ;
        RECT 272.585 62.080 272.840 62.650 ;
        RECT 273.010 62.420 273.340 62.820 ;
        RECT 273.765 62.285 274.295 62.650 ;
        RECT 273.765 62.250 273.940 62.285 ;
        RECT 273.010 62.080 273.940 62.250 ;
        RECT 269.960 61.120 270.170 62.020 ;
        RECT 270.340 61.290 271.030 61.850 ;
        RECT 271.200 61.530 271.720 62.070 ;
        RECT 271.890 61.360 272.410 61.900 ;
        RECT 269.960 60.900 270.915 61.120 ;
        RECT 270.190 60.270 270.460 60.730 ;
        RECT 270.630 60.440 270.915 60.900 ;
        RECT 271.200 60.270 272.410 61.360 ;
        RECT 272.585 61.410 272.755 62.080 ;
        RECT 273.010 61.910 273.180 62.080 ;
        RECT 272.925 61.580 273.180 61.910 ;
        RECT 273.405 61.580 273.600 61.910 ;
        RECT 272.585 60.440 272.920 61.410 ;
        RECT 273.090 60.270 273.260 61.410 ;
        RECT 273.430 60.610 273.600 61.580 ;
        RECT 273.770 60.950 273.940 62.080 ;
        RECT 274.110 61.290 274.280 62.090 ;
        RECT 274.485 61.800 274.760 62.650 ;
        RECT 274.480 61.630 274.760 61.800 ;
        RECT 274.485 61.490 274.760 61.630 ;
        RECT 274.930 61.290 275.120 62.650 ;
        RECT 275.300 62.285 275.810 62.820 ;
        RECT 276.030 62.010 276.275 62.615 ;
        RECT 276.720 62.050 278.390 62.820 ;
        RECT 278.560 62.190 278.900 62.650 ;
        RECT 279.070 62.360 279.240 62.820 ;
        RECT 279.870 62.385 280.230 62.650 ;
        RECT 279.875 62.380 280.230 62.385 ;
        RECT 279.880 62.370 280.230 62.380 ;
        RECT 279.885 62.365 280.230 62.370 ;
        RECT 279.890 62.355 280.230 62.365 ;
        RECT 280.470 62.360 280.640 62.820 ;
        RECT 279.895 62.350 280.230 62.355 ;
        RECT 279.905 62.340 280.230 62.350 ;
        RECT 279.915 62.330 280.230 62.340 ;
        RECT 279.410 62.190 279.740 62.270 ;
        RECT 275.320 61.840 276.550 62.010 ;
        RECT 274.110 61.120 275.120 61.290 ;
        RECT 275.290 61.275 276.040 61.465 ;
        RECT 273.770 60.780 274.895 60.950 ;
        RECT 275.290 60.610 275.460 61.275 ;
        RECT 276.210 61.030 276.550 61.840 ;
        RECT 276.720 61.530 277.470 62.050 ;
        RECT 278.560 62.000 279.740 62.190 ;
        RECT 279.930 62.190 280.230 62.330 ;
        RECT 279.930 62.000 280.640 62.190 ;
        RECT 277.640 61.360 278.390 61.880 ;
        RECT 273.430 60.440 275.460 60.610 ;
        RECT 275.630 60.270 275.800 61.030 ;
        RECT 276.035 60.620 276.550 61.030 ;
        RECT 276.720 60.270 278.390 61.360 ;
        RECT 278.560 61.630 278.890 61.830 ;
        RECT 279.200 61.810 279.530 61.830 ;
        RECT 279.080 61.630 279.530 61.810 ;
        RECT 278.560 61.290 278.790 61.630 ;
        RECT 278.570 60.270 278.900 60.990 ;
        RECT 279.080 60.515 279.295 61.630 ;
        RECT 279.700 61.600 280.170 61.830 ;
        RECT 280.355 61.430 280.640 62.000 ;
        RECT 280.810 61.875 281.150 62.650 ;
        RECT 279.490 61.215 280.640 61.430 ;
        RECT 279.490 60.440 279.820 61.215 ;
        RECT 279.990 60.270 280.700 61.045 ;
        RECT 280.870 60.440 281.150 61.875 ;
        RECT 282.245 62.080 282.500 62.650 ;
        RECT 282.670 62.420 283.000 62.820 ;
        RECT 283.425 62.285 283.955 62.650 ;
        RECT 284.145 62.480 284.420 62.650 ;
        RECT 284.140 62.310 284.420 62.480 ;
        RECT 283.425 62.250 283.600 62.285 ;
        RECT 282.670 62.080 283.600 62.250 ;
        RECT 282.245 61.410 282.415 62.080 ;
        RECT 282.670 61.910 282.840 62.080 ;
        RECT 282.585 61.580 282.840 61.910 ;
        RECT 283.065 61.580 283.260 61.910 ;
        RECT 282.245 60.440 282.580 61.410 ;
        RECT 282.750 60.270 282.920 61.410 ;
        RECT 283.090 60.610 283.260 61.580 ;
        RECT 283.430 60.950 283.600 62.080 ;
        RECT 283.770 61.290 283.940 62.090 ;
        RECT 284.145 61.490 284.420 62.310 ;
        RECT 284.590 61.290 284.780 62.650 ;
        RECT 284.960 62.285 285.470 62.820 ;
        RECT 285.690 62.010 285.935 62.615 ;
        RECT 286.655 62.010 286.900 62.615 ;
        RECT 287.120 62.285 287.630 62.820 ;
        RECT 284.980 61.840 286.210 62.010 ;
        RECT 283.770 61.120 284.780 61.290 ;
        RECT 284.950 61.275 285.700 61.465 ;
        RECT 283.430 60.780 284.555 60.950 ;
        RECT 284.950 60.610 285.120 61.275 ;
        RECT 285.870 61.030 286.210 61.840 ;
        RECT 283.090 60.440 285.120 60.610 ;
        RECT 285.290 60.270 285.460 61.030 ;
        RECT 285.695 60.620 286.210 61.030 ;
        RECT 286.380 61.840 287.610 62.010 ;
        RECT 286.380 61.030 286.720 61.840 ;
        RECT 286.890 61.275 287.640 61.465 ;
        RECT 286.380 60.620 286.895 61.030 ;
        RECT 287.130 60.270 287.300 61.030 ;
        RECT 287.470 60.610 287.640 61.275 ;
        RECT 287.810 61.290 288.000 62.650 ;
        RECT 288.170 62.480 288.445 62.650 ;
        RECT 288.170 62.310 288.450 62.480 ;
        RECT 288.170 61.490 288.445 62.310 ;
        RECT 288.635 62.285 289.165 62.650 ;
        RECT 289.590 62.420 289.920 62.820 ;
        RECT 288.990 62.250 289.165 62.285 ;
        RECT 288.650 61.290 288.820 62.090 ;
        RECT 287.810 61.120 288.820 61.290 ;
        RECT 288.990 62.080 289.920 62.250 ;
        RECT 290.090 62.080 290.345 62.650 ;
        RECT 290.980 62.095 291.270 62.820 ;
        RECT 288.990 60.950 289.160 62.080 ;
        RECT 289.750 61.910 289.920 62.080 ;
        RECT 288.035 60.780 289.160 60.950 ;
        RECT 289.330 61.580 289.525 61.910 ;
        RECT 289.750 61.580 290.005 61.910 ;
        RECT 289.330 60.610 289.500 61.580 ;
        RECT 290.175 61.410 290.345 62.080 ;
        RECT 291.440 62.070 292.650 62.820 ;
        RECT 292.910 62.270 293.080 62.650 ;
        RECT 293.260 62.440 293.590 62.820 ;
        RECT 292.910 62.100 293.575 62.270 ;
        RECT 293.770 62.145 294.030 62.650 ;
        RECT 291.440 61.530 291.960 62.070 ;
        RECT 287.470 60.440 289.500 60.610 ;
        RECT 289.670 60.270 289.840 61.410 ;
        RECT 290.010 60.440 290.345 61.410 ;
        RECT 290.980 60.270 291.270 61.435 ;
        RECT 292.130 61.360 292.650 61.900 ;
        RECT 292.840 61.550 293.170 61.920 ;
        RECT 293.405 61.845 293.575 62.100 ;
        RECT 293.405 61.515 293.690 61.845 ;
        RECT 293.405 61.370 293.575 61.515 ;
        RECT 291.440 60.270 292.650 61.360 ;
        RECT 292.910 61.200 293.575 61.370 ;
        RECT 293.860 61.345 294.030 62.145 ;
        RECT 294.205 62.270 294.460 62.560 ;
        RECT 294.630 62.440 294.960 62.820 ;
        RECT 294.205 62.100 294.955 62.270 ;
        RECT 292.910 60.440 293.080 61.200 ;
        RECT 293.260 60.270 293.590 61.030 ;
        RECT 293.760 60.440 294.030 61.345 ;
        RECT 294.205 61.280 294.555 61.930 ;
        RECT 294.725 61.110 294.955 62.100 ;
        RECT 294.205 60.940 294.955 61.110 ;
        RECT 294.205 60.440 294.460 60.940 ;
        RECT 294.630 60.270 294.960 60.770 ;
        RECT 295.130 60.440 295.300 62.560 ;
        RECT 295.660 62.460 295.990 62.820 ;
        RECT 296.160 62.430 296.655 62.600 ;
        RECT 296.860 62.430 297.715 62.600 ;
        RECT 295.530 61.240 295.990 62.290 ;
        RECT 295.470 60.455 295.795 61.240 ;
        RECT 296.160 61.070 296.330 62.430 ;
        RECT 296.500 61.520 296.850 62.140 ;
        RECT 297.020 61.920 297.375 62.140 ;
        RECT 297.020 61.330 297.190 61.920 ;
        RECT 297.545 61.720 297.715 62.430 ;
        RECT 298.590 62.360 298.920 62.820 ;
        RECT 299.130 62.460 299.480 62.630 ;
        RECT 297.920 61.890 298.710 62.140 ;
        RECT 299.130 62.070 299.390 62.460 ;
        RECT 299.700 62.370 300.650 62.650 ;
        RECT 300.820 62.380 301.010 62.820 ;
        RECT 301.180 62.440 302.250 62.610 ;
        RECT 298.880 61.720 299.050 61.900 ;
        RECT 296.160 60.900 296.555 61.070 ;
        RECT 296.725 60.940 297.190 61.330 ;
        RECT 297.360 61.550 299.050 61.720 ;
        RECT 296.385 60.770 296.555 60.900 ;
        RECT 297.360 60.770 297.530 61.550 ;
        RECT 299.220 61.380 299.390 62.070 ;
        RECT 297.890 61.210 299.390 61.380 ;
        RECT 299.580 61.410 299.790 62.200 ;
        RECT 299.960 61.580 300.310 62.200 ;
        RECT 300.480 61.590 300.650 62.370 ;
        RECT 301.180 62.210 301.350 62.440 ;
        RECT 300.820 62.040 301.350 62.210 ;
        RECT 300.820 61.760 301.040 62.040 ;
        RECT 301.520 61.870 301.760 62.270 ;
        RECT 300.480 61.420 300.885 61.590 ;
        RECT 301.220 61.500 301.760 61.870 ;
        RECT 301.930 62.085 302.250 62.440 ;
        RECT 302.495 62.360 302.800 62.820 ;
        RECT 302.970 62.110 303.220 62.640 ;
        RECT 301.930 61.910 302.255 62.085 ;
        RECT 301.930 61.610 302.845 61.910 ;
        RECT 302.105 61.580 302.845 61.610 ;
        RECT 299.580 61.250 300.255 61.410 ;
        RECT 300.715 61.330 300.885 61.420 ;
        RECT 299.580 61.240 300.545 61.250 ;
        RECT 299.220 61.070 299.390 61.210 ;
        RECT 295.965 60.270 296.215 60.730 ;
        RECT 296.385 60.440 296.635 60.770 ;
        RECT 296.850 60.440 297.530 60.770 ;
        RECT 297.700 60.870 298.775 61.040 ;
        RECT 299.220 60.900 299.780 61.070 ;
        RECT 300.085 60.950 300.545 61.240 ;
        RECT 300.715 61.160 301.935 61.330 ;
        RECT 297.700 60.530 297.870 60.870 ;
        RECT 298.105 60.270 298.435 60.700 ;
        RECT 298.605 60.530 298.775 60.870 ;
        RECT 299.070 60.270 299.440 60.730 ;
        RECT 299.610 60.440 299.780 60.900 ;
        RECT 300.715 60.780 300.885 61.160 ;
        RECT 302.105 60.990 302.275 61.580 ;
        RECT 303.015 61.460 303.220 62.110 ;
        RECT 303.390 62.065 303.640 62.820 ;
        RECT 303.860 62.275 309.205 62.820 ;
        RECT 300.015 60.440 300.885 60.780 ;
        RECT 301.475 60.820 302.275 60.990 ;
        RECT 301.055 60.270 301.305 60.730 ;
        RECT 301.475 60.530 301.645 60.820 ;
        RECT 301.825 60.270 302.155 60.650 ;
        RECT 302.495 60.270 302.800 61.410 ;
        RECT 302.970 60.580 303.220 61.460 ;
        RECT 305.445 61.445 305.785 62.275 ;
        RECT 309.840 62.070 311.050 62.820 ;
        RECT 303.390 60.270 303.640 61.410 ;
        RECT 307.265 60.705 307.615 61.955 ;
        RECT 309.840 61.360 310.360 61.900 ;
        RECT 310.530 61.530 311.050 62.070 ;
        RECT 303.860 60.270 309.205 60.705 ;
        RECT 309.840 60.270 311.050 61.360 ;
        RECT 162.095 60.100 311.135 60.270 ;
        RECT 162.180 59.010 163.390 60.100 ;
        RECT 163.560 59.010 165.230 60.100 ;
        RECT 165.405 59.430 165.660 59.930 ;
        RECT 165.830 59.600 166.160 60.100 ;
        RECT 165.405 59.260 166.155 59.430 ;
        RECT 162.180 58.300 162.700 58.840 ;
        RECT 162.870 58.470 163.390 59.010 ;
        RECT 163.560 58.320 164.310 58.840 ;
        RECT 164.480 58.490 165.230 59.010 ;
        RECT 165.405 58.440 165.755 59.090 ;
        RECT 162.180 57.550 163.390 58.300 ;
        RECT 163.560 57.550 165.230 58.320 ;
        RECT 165.925 58.270 166.155 59.260 ;
        RECT 165.405 58.100 166.155 58.270 ;
        RECT 165.405 57.810 165.660 58.100 ;
        RECT 165.830 57.550 166.160 57.930 ;
        RECT 166.330 57.810 166.500 59.930 ;
        RECT 166.670 59.130 166.995 59.915 ;
        RECT 167.165 59.640 167.415 60.100 ;
        RECT 167.585 59.600 167.835 59.930 ;
        RECT 168.050 59.600 168.730 59.930 ;
        RECT 167.585 59.470 167.755 59.600 ;
        RECT 167.360 59.300 167.755 59.470 ;
        RECT 166.730 58.080 167.190 59.130 ;
        RECT 167.360 57.940 167.530 59.300 ;
        RECT 167.925 59.040 168.390 59.430 ;
        RECT 167.700 58.230 168.050 58.850 ;
        RECT 168.220 58.450 168.390 59.040 ;
        RECT 168.560 58.820 168.730 59.600 ;
        RECT 168.900 59.500 169.070 59.840 ;
        RECT 169.305 59.670 169.635 60.100 ;
        RECT 169.805 59.500 169.975 59.840 ;
        RECT 170.270 59.640 170.640 60.100 ;
        RECT 168.900 59.330 169.975 59.500 ;
        RECT 170.810 59.470 170.980 59.930 ;
        RECT 171.215 59.590 172.085 59.930 ;
        RECT 172.255 59.640 172.505 60.100 ;
        RECT 170.420 59.300 170.980 59.470 ;
        RECT 170.420 59.160 170.590 59.300 ;
        RECT 169.090 58.990 170.590 59.160 ;
        RECT 171.285 59.130 171.745 59.420 ;
        RECT 168.560 58.650 170.250 58.820 ;
        RECT 168.220 58.230 168.575 58.450 ;
        RECT 168.745 57.940 168.915 58.650 ;
        RECT 169.120 58.230 169.910 58.480 ;
        RECT 170.080 58.470 170.250 58.650 ;
        RECT 170.420 58.300 170.590 58.990 ;
        RECT 166.860 57.550 167.190 57.910 ;
        RECT 167.360 57.770 167.855 57.940 ;
        RECT 168.060 57.770 168.915 57.940 ;
        RECT 169.790 57.550 170.120 58.010 ;
        RECT 170.330 57.910 170.590 58.300 ;
        RECT 170.780 59.120 171.745 59.130 ;
        RECT 171.915 59.210 172.085 59.590 ;
        RECT 172.675 59.550 172.845 59.840 ;
        RECT 173.025 59.720 173.355 60.100 ;
        RECT 172.675 59.380 173.475 59.550 ;
        RECT 170.780 58.960 171.455 59.120 ;
        RECT 171.915 59.040 173.135 59.210 ;
        RECT 170.780 58.170 170.990 58.960 ;
        RECT 171.915 58.950 172.085 59.040 ;
        RECT 171.160 58.170 171.510 58.790 ;
        RECT 171.680 58.780 172.085 58.950 ;
        RECT 171.680 58.000 171.850 58.780 ;
        RECT 172.020 58.330 172.240 58.610 ;
        RECT 172.420 58.500 172.960 58.870 ;
        RECT 173.305 58.790 173.475 59.380 ;
        RECT 173.695 58.960 174.000 60.100 ;
        RECT 174.170 58.910 174.420 59.790 ;
        RECT 174.590 58.960 174.840 60.100 ;
        RECT 175.060 58.935 175.350 60.100 ;
        RECT 175.985 58.960 176.320 59.930 ;
        RECT 176.490 58.960 176.660 60.100 ;
        RECT 176.830 59.760 178.860 59.930 ;
        RECT 173.305 58.760 174.045 58.790 ;
        RECT 172.020 58.160 172.550 58.330 ;
        RECT 170.330 57.740 170.680 57.910 ;
        RECT 170.900 57.720 171.850 58.000 ;
        RECT 172.020 57.550 172.210 57.990 ;
        RECT 172.380 57.930 172.550 58.160 ;
        RECT 172.720 58.100 172.960 58.500 ;
        RECT 173.130 58.460 174.045 58.760 ;
        RECT 173.130 58.285 173.455 58.460 ;
        RECT 173.130 57.930 173.450 58.285 ;
        RECT 174.215 58.260 174.420 58.910 ;
        RECT 172.380 57.760 173.450 57.930 ;
        RECT 173.695 57.550 174.000 58.010 ;
        RECT 174.170 57.730 174.420 58.260 ;
        RECT 174.590 57.550 174.840 58.305 ;
        RECT 175.985 58.290 176.155 58.960 ;
        RECT 176.830 58.790 177.000 59.760 ;
        RECT 176.325 58.460 176.580 58.790 ;
        RECT 176.805 58.460 177.000 58.790 ;
        RECT 177.170 59.420 178.295 59.590 ;
        RECT 176.410 58.290 176.580 58.460 ;
        RECT 177.170 58.290 177.340 59.420 ;
        RECT 175.060 57.550 175.350 58.275 ;
        RECT 175.985 57.720 176.240 58.290 ;
        RECT 176.410 58.120 177.340 58.290 ;
        RECT 177.510 59.080 178.520 59.250 ;
        RECT 177.510 58.280 177.680 59.080 ;
        RECT 177.885 58.400 178.160 58.880 ;
        RECT 177.880 58.230 178.160 58.400 ;
        RECT 177.165 58.085 177.340 58.120 ;
        RECT 176.410 57.550 176.740 57.950 ;
        RECT 177.165 57.720 177.695 58.085 ;
        RECT 177.885 57.720 178.160 58.230 ;
        RECT 178.330 57.720 178.520 59.080 ;
        RECT 178.690 59.095 178.860 59.760 ;
        RECT 179.030 59.340 179.200 60.100 ;
        RECT 179.435 59.340 179.950 59.750 ;
        RECT 178.690 58.905 179.440 59.095 ;
        RECT 179.610 58.530 179.950 59.340 ;
        RECT 178.720 58.360 179.950 58.530 ;
        RECT 180.125 58.960 180.460 59.930 ;
        RECT 180.630 58.960 180.800 60.100 ;
        RECT 180.970 59.760 183.000 59.930 ;
        RECT 178.700 57.550 179.210 58.085 ;
        RECT 179.430 57.755 179.675 58.360 ;
        RECT 180.125 58.290 180.295 58.960 ;
        RECT 180.970 58.790 181.140 59.760 ;
        RECT 180.465 58.460 180.720 58.790 ;
        RECT 180.945 58.460 181.140 58.790 ;
        RECT 181.310 59.420 182.435 59.590 ;
        RECT 180.550 58.290 180.720 58.460 ;
        RECT 181.310 58.290 181.480 59.420 ;
        RECT 180.125 57.720 180.380 58.290 ;
        RECT 180.550 58.120 181.480 58.290 ;
        RECT 181.650 59.080 182.660 59.250 ;
        RECT 181.650 58.280 181.820 59.080 ;
        RECT 181.305 58.085 181.480 58.120 ;
        RECT 180.550 57.550 180.880 57.950 ;
        RECT 181.305 57.720 181.835 58.085 ;
        RECT 182.025 58.060 182.300 58.880 ;
        RECT 182.020 57.890 182.300 58.060 ;
        RECT 182.025 57.720 182.300 57.890 ;
        RECT 182.470 57.720 182.660 59.080 ;
        RECT 182.830 59.095 183.000 59.760 ;
        RECT 183.170 59.340 183.340 60.100 ;
        RECT 183.575 59.340 184.090 59.750 ;
        RECT 182.830 58.905 183.580 59.095 ;
        RECT 183.750 58.530 184.090 59.340 ;
        RECT 184.260 59.010 187.770 60.100 ;
        RECT 187.945 59.430 188.200 59.930 ;
        RECT 188.370 59.600 188.700 60.100 ;
        RECT 187.945 59.260 188.695 59.430 ;
        RECT 182.860 58.360 184.090 58.530 ;
        RECT 182.840 57.550 183.350 58.085 ;
        RECT 183.570 57.755 183.815 58.360 ;
        RECT 184.260 58.320 185.910 58.840 ;
        RECT 186.080 58.490 187.770 59.010 ;
        RECT 187.945 58.440 188.295 59.090 ;
        RECT 184.260 57.550 187.770 58.320 ;
        RECT 188.465 58.270 188.695 59.260 ;
        RECT 187.945 58.100 188.695 58.270 ;
        RECT 187.945 57.810 188.200 58.100 ;
        RECT 188.370 57.550 188.700 57.930 ;
        RECT 188.870 57.810 189.040 59.930 ;
        RECT 189.210 59.130 189.535 59.915 ;
        RECT 189.705 59.640 189.955 60.100 ;
        RECT 190.125 59.600 190.375 59.930 ;
        RECT 190.590 59.600 191.270 59.930 ;
        RECT 190.125 59.470 190.295 59.600 ;
        RECT 189.900 59.300 190.295 59.470 ;
        RECT 189.270 58.080 189.730 59.130 ;
        RECT 189.900 57.940 190.070 59.300 ;
        RECT 190.465 59.040 190.930 59.430 ;
        RECT 190.240 58.230 190.590 58.850 ;
        RECT 190.760 58.450 190.930 59.040 ;
        RECT 191.100 58.820 191.270 59.600 ;
        RECT 191.440 59.500 191.610 59.840 ;
        RECT 191.845 59.670 192.175 60.100 ;
        RECT 192.345 59.500 192.515 59.840 ;
        RECT 192.810 59.640 193.180 60.100 ;
        RECT 191.440 59.330 192.515 59.500 ;
        RECT 193.350 59.470 193.520 59.930 ;
        RECT 193.755 59.590 194.625 59.930 ;
        RECT 194.795 59.640 195.045 60.100 ;
        RECT 192.960 59.300 193.520 59.470 ;
        RECT 192.960 59.160 193.130 59.300 ;
        RECT 191.630 58.990 193.130 59.160 ;
        RECT 193.825 59.130 194.285 59.420 ;
        RECT 191.100 58.650 192.790 58.820 ;
        RECT 190.760 58.230 191.115 58.450 ;
        RECT 191.285 57.940 191.455 58.650 ;
        RECT 191.660 58.230 192.450 58.480 ;
        RECT 192.620 58.470 192.790 58.650 ;
        RECT 192.960 58.300 193.130 58.990 ;
        RECT 189.400 57.550 189.730 57.910 ;
        RECT 189.900 57.770 190.395 57.940 ;
        RECT 190.600 57.770 191.455 57.940 ;
        RECT 192.330 57.550 192.660 58.010 ;
        RECT 192.870 57.910 193.130 58.300 ;
        RECT 193.320 59.120 194.285 59.130 ;
        RECT 194.455 59.210 194.625 59.590 ;
        RECT 195.215 59.550 195.385 59.840 ;
        RECT 195.565 59.720 195.895 60.100 ;
        RECT 195.215 59.380 196.015 59.550 ;
        RECT 193.320 58.960 193.995 59.120 ;
        RECT 194.455 59.040 195.675 59.210 ;
        RECT 193.320 58.170 193.530 58.960 ;
        RECT 194.455 58.950 194.625 59.040 ;
        RECT 193.700 58.170 194.050 58.790 ;
        RECT 194.220 58.780 194.625 58.950 ;
        RECT 194.220 58.000 194.390 58.780 ;
        RECT 194.560 58.330 194.780 58.610 ;
        RECT 194.960 58.500 195.500 58.870 ;
        RECT 195.845 58.760 196.015 59.380 ;
        RECT 196.190 59.040 196.360 60.100 ;
        RECT 196.570 59.090 196.860 59.930 ;
        RECT 197.030 59.260 197.200 60.100 ;
        RECT 197.410 59.090 197.660 59.930 ;
        RECT 197.870 59.260 198.040 60.100 ;
        RECT 196.570 58.920 198.295 59.090 ;
        RECT 194.560 58.160 195.090 58.330 ;
        RECT 192.870 57.740 193.220 57.910 ;
        RECT 193.440 57.720 194.390 58.000 ;
        RECT 194.560 57.550 194.750 57.990 ;
        RECT 194.920 57.930 195.090 58.160 ;
        RECT 195.260 58.100 195.500 58.500 ;
        RECT 195.670 58.750 196.015 58.760 ;
        RECT 195.670 58.540 197.700 58.750 ;
        RECT 195.670 58.285 195.995 58.540 ;
        RECT 197.885 58.370 198.295 58.920 ;
        RECT 195.670 57.930 195.990 58.285 ;
        RECT 194.920 57.760 195.990 57.930 ;
        RECT 196.190 57.550 196.360 58.360 ;
        RECT 196.530 58.200 198.295 58.370 ;
        RECT 198.520 59.025 198.790 59.930 ;
        RECT 198.960 59.340 199.290 60.100 ;
        RECT 199.470 59.170 199.640 59.930 ;
        RECT 198.520 58.225 198.690 59.025 ;
        RECT 198.975 59.000 199.640 59.170 ;
        RECT 198.975 58.855 199.145 59.000 ;
        RECT 200.820 58.935 201.110 60.100 ;
        RECT 201.280 59.010 202.950 60.100 ;
        RECT 198.860 58.525 199.145 58.855 ;
        RECT 198.975 58.270 199.145 58.525 ;
        RECT 199.380 58.450 199.710 58.820 ;
        RECT 201.280 58.320 202.030 58.840 ;
        RECT 202.200 58.490 202.950 59.010 ;
        RECT 203.125 58.960 203.460 59.930 ;
        RECT 203.630 58.960 203.800 60.100 ;
        RECT 203.970 59.760 206.000 59.930 ;
        RECT 196.530 57.720 196.860 58.200 ;
        RECT 197.030 57.550 197.200 58.020 ;
        RECT 197.370 57.720 197.700 58.200 ;
        RECT 197.870 57.550 198.040 58.020 ;
        RECT 198.520 57.720 198.780 58.225 ;
        RECT 198.975 58.100 199.640 58.270 ;
        RECT 198.960 57.550 199.290 57.930 ;
        RECT 199.470 57.720 199.640 58.100 ;
        RECT 200.820 57.550 201.110 58.275 ;
        RECT 201.280 57.550 202.950 58.320 ;
        RECT 203.125 58.290 203.295 58.960 ;
        RECT 203.970 58.790 204.140 59.760 ;
        RECT 203.465 58.460 203.720 58.790 ;
        RECT 203.945 58.460 204.140 58.790 ;
        RECT 204.310 59.420 205.435 59.590 ;
        RECT 203.550 58.290 203.720 58.460 ;
        RECT 204.310 58.290 204.480 59.420 ;
        RECT 203.125 57.720 203.380 58.290 ;
        RECT 203.550 58.120 204.480 58.290 ;
        RECT 204.650 59.080 205.660 59.250 ;
        RECT 204.650 58.280 204.820 59.080 ;
        RECT 205.025 58.740 205.300 58.880 ;
        RECT 205.020 58.570 205.300 58.740 ;
        RECT 204.305 58.085 204.480 58.120 ;
        RECT 203.550 57.550 203.880 57.950 ;
        RECT 204.305 57.720 204.835 58.085 ;
        RECT 205.025 57.720 205.300 58.570 ;
        RECT 205.470 57.720 205.660 59.080 ;
        RECT 205.830 59.095 206.000 59.760 ;
        RECT 206.170 59.340 206.340 60.100 ;
        RECT 206.575 59.340 207.090 59.750 ;
        RECT 205.830 58.905 206.580 59.095 ;
        RECT 206.750 58.530 207.090 59.340 ;
        RECT 205.860 58.360 207.090 58.530 ;
        RECT 207.260 59.130 207.570 59.930 ;
        RECT 207.740 59.300 208.050 60.100 ;
        RECT 208.220 59.470 208.480 59.930 ;
        RECT 208.650 59.640 208.905 60.100 ;
        RECT 209.080 59.470 209.340 59.930 ;
        RECT 208.220 59.300 209.340 59.470 ;
        RECT 207.260 58.960 208.290 59.130 ;
        RECT 205.840 57.550 206.350 58.085 ;
        RECT 206.570 57.755 206.815 58.360 ;
        RECT 207.260 58.050 207.430 58.960 ;
        RECT 207.600 58.220 207.950 58.790 ;
        RECT 208.120 58.710 208.290 58.960 ;
        RECT 209.080 59.050 209.340 59.300 ;
        RECT 209.510 59.230 209.795 60.100 ;
        RECT 210.020 59.665 215.365 60.100 ;
        RECT 209.080 58.880 209.835 59.050 ;
        RECT 208.120 58.540 209.260 58.710 ;
        RECT 209.430 58.370 209.835 58.880 ;
        RECT 208.185 58.200 209.835 58.370 ;
        RECT 207.260 57.720 207.560 58.050 ;
        RECT 207.730 57.550 208.005 58.030 ;
        RECT 208.185 57.810 208.480 58.200 ;
        RECT 208.650 57.550 208.905 58.030 ;
        RECT 209.080 57.810 209.340 58.200 ;
        RECT 211.605 58.095 211.945 58.925 ;
        RECT 213.425 58.415 213.775 59.665 ;
        RECT 215.540 59.010 217.210 60.100 ;
        RECT 215.540 58.320 216.290 58.840 ;
        RECT 216.460 58.490 217.210 59.010 ;
        RECT 217.380 58.960 217.670 60.100 ;
        RECT 217.840 59.380 218.290 59.930 ;
        RECT 218.480 59.380 218.810 60.100 ;
        RECT 209.510 57.550 209.790 58.030 ;
        RECT 210.020 57.550 215.365 58.095 ;
        RECT 215.540 57.550 217.210 58.320 ;
        RECT 217.380 57.550 217.670 58.350 ;
        RECT 217.840 58.010 218.090 59.380 ;
        RECT 219.020 59.210 219.320 59.760 ;
        RECT 219.490 59.430 219.770 60.100 ;
        RECT 218.380 59.040 219.320 59.210 ;
        RECT 218.380 58.790 218.550 59.040 ;
        RECT 219.655 58.790 219.970 59.230 ;
        RECT 220.140 59.010 223.650 60.100 ;
        RECT 218.260 58.460 218.550 58.790 ;
        RECT 218.720 58.540 219.050 58.790 ;
        RECT 219.280 58.540 219.970 58.790 ;
        RECT 218.380 58.370 218.550 58.460 ;
        RECT 218.380 58.180 219.770 58.370 ;
        RECT 217.840 57.720 218.390 58.010 ;
        RECT 218.560 57.550 218.810 58.010 ;
        RECT 219.440 57.820 219.770 58.180 ;
        RECT 220.140 58.320 221.790 58.840 ;
        RECT 221.960 58.490 223.650 59.010 ;
        RECT 224.315 59.310 224.850 59.930 ;
        RECT 220.140 57.550 223.650 58.320 ;
        RECT 224.315 58.290 224.630 59.310 ;
        RECT 225.020 59.300 225.350 60.100 ;
        RECT 225.835 59.130 226.225 59.305 ;
        RECT 224.800 58.960 226.225 59.130 ;
        RECT 224.800 58.460 224.970 58.960 ;
        RECT 224.315 57.720 224.930 58.290 ;
        RECT 225.220 58.230 225.485 58.790 ;
        RECT 225.655 58.060 225.825 58.960 ;
        RECT 226.580 58.935 226.870 60.100 ;
        RECT 227.245 59.130 227.575 59.930 ;
        RECT 227.745 59.300 228.075 60.100 ;
        RECT 228.375 59.130 228.705 59.930 ;
        RECT 229.350 59.300 229.600 60.100 ;
        RECT 227.245 58.960 229.680 59.130 ;
        RECT 229.870 58.960 230.040 60.100 ;
        RECT 230.210 58.960 230.550 59.930 ;
        RECT 230.720 59.760 231.900 59.930 ;
        RECT 230.720 58.960 231.060 59.760 ;
        RECT 225.995 58.230 226.350 58.790 ;
        RECT 227.040 58.540 227.390 58.790 ;
        RECT 227.575 58.330 227.745 58.960 ;
        RECT 227.915 58.540 228.245 58.740 ;
        RECT 228.415 58.540 228.745 58.740 ;
        RECT 228.915 58.540 229.335 58.740 ;
        RECT 229.510 58.710 229.680 58.960 ;
        RECT 229.510 58.540 230.205 58.710 ;
        RECT 225.100 57.550 225.315 58.060 ;
        RECT 225.545 57.730 225.825 58.060 ;
        RECT 226.005 57.550 226.245 58.060 ;
        RECT 226.580 57.550 226.870 58.275 ;
        RECT 227.245 57.720 227.745 58.330 ;
        RECT 228.375 58.200 229.600 58.370 ;
        RECT 230.375 58.350 230.550 58.960 ;
        RECT 231.230 58.790 231.465 59.515 ;
        RECT 231.635 59.130 231.900 59.760 ;
        RECT 232.070 59.300 232.770 60.100 ;
        RECT 231.635 58.960 232.725 59.130 ;
        RECT 230.720 58.540 231.060 58.790 ;
        RECT 231.230 58.540 231.690 58.790 ;
        RECT 231.860 58.540 232.335 58.790 ;
        RECT 232.505 58.710 232.725 58.960 ;
        RECT 232.980 59.090 233.230 59.930 ;
        RECT 233.400 59.260 233.650 60.100 ;
        RECT 233.820 59.090 234.070 59.930 ;
        RECT 234.240 59.260 234.490 60.100 ;
        RECT 232.980 58.920 234.690 59.090 ;
        RECT 232.505 58.540 234.230 58.710 ;
        RECT 232.505 58.370 232.725 58.540 ;
        RECT 234.400 58.370 234.690 58.920 ;
        RECT 228.375 57.720 228.705 58.200 ;
        RECT 228.875 57.550 229.100 58.010 ;
        RECT 229.270 57.720 229.600 58.200 ;
        RECT 229.790 57.550 230.040 58.350 ;
        RECT 230.210 57.720 230.550 58.350 ;
        RECT 230.720 58.190 232.725 58.370 ;
        RECT 232.940 58.200 234.690 58.370 ;
        RECT 234.870 59.040 235.200 59.890 ;
        RECT 234.870 58.910 235.090 59.040 ;
        RECT 235.370 58.960 235.620 60.100 ;
        RECT 235.810 59.460 236.060 59.880 ;
        RECT 236.290 59.630 236.620 60.100 ;
        RECT 236.850 59.460 237.100 59.880 ;
        RECT 235.810 59.290 237.100 59.460 ;
        RECT 237.280 59.460 237.610 59.890 ;
        RECT 237.280 59.290 237.735 59.460 ;
        RECT 234.870 58.275 235.060 58.910 ;
        RECT 235.800 58.790 236.015 59.120 ;
        RECT 235.230 58.460 235.540 58.790 ;
        RECT 235.710 58.460 236.015 58.790 ;
        RECT 236.190 58.460 236.475 59.120 ;
        RECT 236.670 58.460 236.935 59.120 ;
        RECT 237.150 58.460 237.395 59.120 ;
        RECT 235.370 58.290 235.540 58.460 ;
        RECT 237.565 58.290 237.735 59.290 ;
        RECT 239.185 59.130 239.575 59.305 ;
        RECT 240.060 59.300 240.390 60.100 ;
        RECT 240.560 59.310 241.095 59.930 ;
        RECT 239.185 58.960 240.610 59.130 ;
        RECT 230.720 57.720 231.060 58.190 ;
        RECT 231.230 57.550 231.400 58.020 ;
        RECT 231.570 57.720 231.900 58.190 ;
        RECT 232.070 57.550 232.770 58.020 ;
        RECT 232.940 57.730 233.270 58.200 ;
        RECT 233.440 57.550 233.610 58.020 ;
        RECT 233.780 57.730 234.110 58.200 ;
        RECT 234.280 57.550 234.450 58.020 ;
        RECT 234.870 57.765 235.200 58.275 ;
        RECT 235.370 58.120 237.735 58.290 ;
        RECT 239.060 58.230 239.415 58.790 ;
        RECT 235.370 57.550 235.700 57.950 ;
        RECT 236.750 57.780 237.080 58.120 ;
        RECT 239.585 58.060 239.755 58.960 ;
        RECT 239.925 58.230 240.190 58.790 ;
        RECT 240.440 58.460 240.610 58.960 ;
        RECT 240.780 58.290 241.095 59.310 ;
        RECT 237.250 57.550 237.580 57.950 ;
        RECT 239.165 57.550 239.405 58.060 ;
        RECT 239.585 57.730 239.865 58.060 ;
        RECT 240.095 57.550 240.310 58.060 ;
        RECT 240.480 57.720 241.095 58.290 ;
        RECT 241.310 59.040 241.640 59.890 ;
        RECT 241.310 58.275 241.500 59.040 ;
        RECT 241.810 58.960 242.060 60.100 ;
        RECT 242.250 59.460 242.500 59.880 ;
        RECT 242.730 59.630 243.060 60.100 ;
        RECT 243.290 59.460 243.540 59.880 ;
        RECT 242.250 59.290 243.540 59.460 ;
        RECT 243.720 59.460 244.050 59.890 ;
        RECT 243.720 59.290 244.175 59.460 ;
        RECT 242.240 58.790 242.455 59.120 ;
        RECT 241.670 58.460 241.980 58.790 ;
        RECT 242.150 58.460 242.455 58.790 ;
        RECT 242.630 58.460 242.915 59.120 ;
        RECT 243.110 58.460 243.375 59.120 ;
        RECT 243.590 58.460 243.835 59.120 ;
        RECT 241.810 58.290 241.980 58.460 ;
        RECT 244.005 58.290 244.175 59.290 ;
        RECT 241.310 57.765 241.640 58.275 ;
        RECT 241.810 58.120 244.175 58.290 ;
        RECT 241.810 57.550 242.140 57.950 ;
        RECT 243.190 57.780 243.520 58.120 ;
        RECT 243.690 57.550 244.020 57.950 ;
        RECT 245.440 57.720 246.190 59.930 ;
        RECT 247.465 59.130 247.855 59.305 ;
        RECT 248.340 59.300 248.670 60.100 ;
        RECT 248.840 59.310 249.375 59.930 ;
        RECT 247.465 58.960 248.890 59.130 ;
        RECT 247.340 58.230 247.695 58.790 ;
        RECT 247.865 58.060 248.035 58.960 ;
        RECT 248.205 58.230 248.470 58.790 ;
        RECT 248.720 58.460 248.890 58.960 ;
        RECT 249.060 58.290 249.375 59.310 ;
        RECT 249.670 59.170 249.840 59.930 ;
        RECT 250.055 59.340 250.385 60.100 ;
        RECT 249.670 59.000 250.385 59.170 ;
        RECT 250.555 59.025 250.810 59.930 ;
        RECT 249.580 58.450 249.935 58.820 ;
        RECT 250.215 58.790 250.385 59.000 ;
        RECT 250.215 58.460 250.470 58.790 ;
        RECT 247.445 57.550 247.685 58.060 ;
        RECT 247.865 57.730 248.145 58.060 ;
        RECT 248.375 57.550 248.590 58.060 ;
        RECT 248.760 57.720 249.375 58.290 ;
        RECT 250.215 58.270 250.385 58.460 ;
        RECT 250.640 58.295 250.810 59.025 ;
        RECT 250.985 58.950 251.245 60.100 ;
        RECT 252.340 58.935 252.630 60.100 ;
        RECT 252.800 59.010 254.010 60.100 ;
        RECT 249.670 58.100 250.385 58.270 ;
        RECT 249.670 57.720 249.840 58.100 ;
        RECT 250.055 57.550 250.385 57.930 ;
        RECT 250.555 57.720 250.810 58.295 ;
        RECT 250.985 57.550 251.245 58.390 ;
        RECT 252.800 58.300 253.320 58.840 ;
        RECT 253.490 58.470 254.010 59.010 ;
        RECT 254.385 59.130 254.715 59.930 ;
        RECT 254.885 59.300 255.215 60.100 ;
        RECT 255.515 59.130 255.845 59.930 ;
        RECT 256.490 59.300 256.740 60.100 ;
        RECT 254.385 58.960 256.820 59.130 ;
        RECT 257.010 58.960 257.180 60.100 ;
        RECT 257.350 58.960 257.690 59.930 ;
        RECT 258.045 59.130 258.435 59.305 ;
        RECT 258.920 59.300 259.250 60.100 ;
        RECT 259.420 59.310 259.955 59.930 ;
        RECT 260.920 59.460 261.250 59.890 ;
        RECT 258.045 58.960 259.470 59.130 ;
        RECT 254.180 58.540 254.530 58.790 ;
        RECT 254.715 58.330 254.885 58.960 ;
        RECT 255.055 58.540 255.385 58.740 ;
        RECT 255.555 58.540 255.885 58.740 ;
        RECT 256.055 58.540 256.475 58.740 ;
        RECT 256.650 58.710 256.820 58.960 ;
        RECT 256.650 58.540 257.345 58.710 ;
        RECT 252.340 57.550 252.630 58.275 ;
        RECT 252.800 57.550 254.010 58.300 ;
        RECT 254.385 57.720 254.885 58.330 ;
        RECT 255.515 58.200 256.740 58.370 ;
        RECT 257.515 58.350 257.690 58.960 ;
        RECT 255.515 57.720 255.845 58.200 ;
        RECT 256.015 57.550 256.240 58.010 ;
        RECT 256.410 57.720 256.740 58.200 ;
        RECT 256.930 57.550 257.180 58.350 ;
        RECT 257.350 57.720 257.690 58.350 ;
        RECT 257.920 58.230 258.275 58.790 ;
        RECT 258.445 58.060 258.615 58.960 ;
        RECT 258.785 58.230 259.050 58.790 ;
        RECT 259.300 58.460 259.470 58.960 ;
        RECT 259.640 58.290 259.955 59.310 ;
        RECT 258.025 57.550 258.265 58.060 ;
        RECT 258.445 57.730 258.725 58.060 ;
        RECT 258.955 57.550 259.170 58.060 ;
        RECT 259.340 57.720 259.955 58.290 ;
        RECT 260.795 59.290 261.250 59.460 ;
        RECT 261.430 59.460 261.680 59.880 ;
        RECT 261.910 59.630 262.240 60.100 ;
        RECT 262.470 59.460 262.720 59.880 ;
        RECT 261.430 59.290 262.720 59.460 ;
        RECT 260.795 58.290 260.965 59.290 ;
        RECT 261.135 58.460 261.380 59.120 ;
        RECT 261.595 58.460 261.860 59.120 ;
        RECT 262.055 58.460 262.340 59.120 ;
        RECT 262.515 58.790 262.730 59.120 ;
        RECT 262.910 58.960 263.160 60.100 ;
        RECT 263.330 59.040 263.660 59.890 ;
        RECT 262.515 58.460 262.820 58.790 ;
        RECT 262.990 58.460 263.300 58.790 ;
        RECT 262.990 58.290 263.160 58.460 ;
        RECT 260.795 58.120 263.160 58.290 ;
        RECT 263.470 58.275 263.660 59.040 ;
        RECT 263.840 58.920 264.160 60.100 ;
        RECT 264.330 59.080 264.530 59.870 ;
        RECT 264.855 59.270 265.240 59.930 ;
        RECT 265.635 59.340 266.420 60.100 ;
        RECT 264.830 59.170 265.240 59.270 ;
        RECT 264.330 58.910 264.660 59.080 ;
        RECT 264.830 58.960 266.440 59.170 ;
        RECT 264.480 58.790 264.660 58.910 ;
        RECT 263.840 58.540 264.305 58.740 ;
        RECT 264.480 58.540 264.810 58.790 ;
        RECT 264.980 58.740 265.445 58.790 ;
        RECT 264.980 58.570 265.450 58.740 ;
        RECT 264.980 58.540 265.445 58.570 ;
        RECT 265.640 58.540 265.995 58.790 ;
        RECT 266.165 58.360 266.440 58.960 ;
        RECT 260.950 57.550 261.280 57.950 ;
        RECT 261.450 57.780 261.780 58.120 ;
        RECT 262.830 57.550 263.160 57.950 ;
        RECT 263.330 57.765 263.660 58.275 ;
        RECT 263.840 58.160 265.020 58.330 ;
        RECT 263.840 57.745 264.180 58.160 ;
        RECT 264.350 57.550 264.520 57.990 ;
        RECT 264.690 57.940 265.020 58.160 ;
        RECT 265.190 58.180 266.440 58.360 ;
        RECT 265.190 58.110 265.555 58.180 ;
        RECT 264.690 57.760 265.940 57.940 ;
        RECT 266.210 57.550 266.380 58.010 ;
        RECT 266.610 57.830 266.890 59.930 ;
        RECT 267.060 59.010 268.270 60.100 ;
        RECT 267.060 58.300 267.580 58.840 ;
        RECT 267.750 58.470 268.270 59.010 ;
        RECT 268.440 58.960 268.825 59.930 ;
        RECT 268.995 59.640 269.320 60.100 ;
        RECT 269.840 59.470 270.120 59.930 ;
        RECT 268.995 59.250 270.120 59.470 ;
        RECT 267.060 57.550 268.270 58.300 ;
        RECT 268.440 58.290 268.720 58.960 ;
        RECT 268.995 58.790 269.445 59.250 ;
        RECT 270.310 59.080 270.710 59.930 ;
        RECT 271.110 59.640 271.380 60.100 ;
        RECT 271.550 59.470 271.835 59.930 ;
        RECT 272.120 59.665 277.465 60.100 ;
        RECT 268.890 58.460 269.445 58.790 ;
        RECT 269.615 58.520 270.710 59.080 ;
        RECT 268.995 58.350 269.445 58.460 ;
        RECT 268.440 57.720 268.825 58.290 ;
        RECT 268.995 58.180 270.120 58.350 ;
        RECT 268.995 57.550 269.320 58.010 ;
        RECT 269.840 57.720 270.120 58.180 ;
        RECT 270.310 57.720 270.710 58.520 ;
        RECT 270.880 59.250 271.835 59.470 ;
        RECT 270.880 58.350 271.090 59.250 ;
        RECT 271.260 58.520 271.950 59.080 ;
        RECT 270.880 58.180 271.835 58.350 ;
        RECT 271.110 57.550 271.380 58.010 ;
        RECT 271.550 57.720 271.835 58.180 ;
        RECT 273.705 58.095 274.045 58.925 ;
        RECT 275.525 58.415 275.875 59.665 ;
        RECT 278.100 58.935 278.390 60.100 ;
        RECT 279.110 59.170 279.280 59.930 ;
        RECT 279.460 59.340 279.790 60.100 ;
        RECT 279.110 59.000 279.775 59.170 ;
        RECT 279.960 59.025 280.230 59.930 ;
        RECT 280.405 59.430 280.660 59.930 ;
        RECT 280.830 59.600 281.160 60.100 ;
        RECT 280.405 59.260 281.155 59.430 ;
        RECT 279.605 58.855 279.775 59.000 ;
        RECT 279.040 58.450 279.370 58.820 ;
        RECT 279.605 58.525 279.890 58.855 ;
        RECT 272.120 57.550 277.465 58.095 ;
        RECT 278.100 57.550 278.390 58.275 ;
        RECT 279.605 58.270 279.775 58.525 ;
        RECT 279.110 58.100 279.775 58.270 ;
        RECT 280.060 58.225 280.230 59.025 ;
        RECT 280.405 58.440 280.755 59.090 ;
        RECT 280.925 58.270 281.155 59.260 ;
        RECT 279.110 57.720 279.280 58.100 ;
        RECT 279.460 57.550 279.790 57.930 ;
        RECT 279.970 57.720 280.230 58.225 ;
        RECT 280.405 58.100 281.155 58.270 ;
        RECT 280.405 57.810 280.660 58.100 ;
        RECT 280.830 57.550 281.160 57.930 ;
        RECT 281.330 57.810 281.500 59.930 ;
        RECT 281.670 59.130 281.995 59.915 ;
        RECT 282.165 59.640 282.415 60.100 ;
        RECT 282.585 59.600 282.835 59.930 ;
        RECT 283.050 59.600 283.730 59.930 ;
        RECT 282.585 59.470 282.755 59.600 ;
        RECT 282.360 59.300 282.755 59.470 ;
        RECT 281.730 58.080 282.190 59.130 ;
        RECT 282.360 57.940 282.530 59.300 ;
        RECT 282.925 59.040 283.390 59.430 ;
        RECT 282.700 58.230 283.050 58.850 ;
        RECT 283.220 58.450 283.390 59.040 ;
        RECT 283.560 58.820 283.730 59.600 ;
        RECT 283.900 59.500 284.070 59.840 ;
        RECT 284.305 59.670 284.635 60.100 ;
        RECT 284.805 59.500 284.975 59.840 ;
        RECT 285.270 59.640 285.640 60.100 ;
        RECT 283.900 59.330 284.975 59.500 ;
        RECT 285.810 59.470 285.980 59.930 ;
        RECT 286.215 59.590 287.085 59.930 ;
        RECT 287.255 59.640 287.505 60.100 ;
        RECT 285.420 59.300 285.980 59.470 ;
        RECT 285.420 59.160 285.590 59.300 ;
        RECT 284.090 58.990 285.590 59.160 ;
        RECT 286.285 59.130 286.745 59.420 ;
        RECT 283.560 58.650 285.250 58.820 ;
        RECT 283.220 58.230 283.575 58.450 ;
        RECT 283.745 57.940 283.915 58.650 ;
        RECT 284.120 58.230 284.910 58.480 ;
        RECT 285.080 58.470 285.250 58.650 ;
        RECT 285.420 58.300 285.590 58.990 ;
        RECT 281.860 57.550 282.190 57.910 ;
        RECT 282.360 57.770 282.855 57.940 ;
        RECT 283.060 57.770 283.915 57.940 ;
        RECT 284.790 57.550 285.120 58.010 ;
        RECT 285.330 57.910 285.590 58.300 ;
        RECT 285.780 59.120 286.745 59.130 ;
        RECT 286.915 59.210 287.085 59.590 ;
        RECT 287.675 59.550 287.845 59.840 ;
        RECT 288.025 59.720 288.355 60.100 ;
        RECT 287.675 59.380 288.475 59.550 ;
        RECT 285.780 58.960 286.455 59.120 ;
        RECT 286.915 59.040 288.135 59.210 ;
        RECT 285.780 58.170 285.990 58.960 ;
        RECT 286.915 58.950 287.085 59.040 ;
        RECT 286.160 58.170 286.510 58.790 ;
        RECT 286.680 58.780 287.085 58.950 ;
        RECT 286.680 58.000 286.850 58.780 ;
        RECT 287.020 58.330 287.240 58.610 ;
        RECT 287.420 58.500 287.960 58.870 ;
        RECT 288.305 58.790 288.475 59.380 ;
        RECT 288.695 58.960 289.000 60.100 ;
        RECT 289.170 58.910 289.425 59.790 ;
        RECT 288.305 58.760 289.045 58.790 ;
        RECT 287.020 58.160 287.550 58.330 ;
        RECT 285.330 57.740 285.680 57.910 ;
        RECT 285.900 57.720 286.850 58.000 ;
        RECT 287.020 57.550 287.210 57.990 ;
        RECT 287.380 57.930 287.550 58.160 ;
        RECT 287.720 58.100 287.960 58.500 ;
        RECT 288.130 58.460 289.045 58.760 ;
        RECT 288.130 58.285 288.455 58.460 ;
        RECT 288.130 57.930 288.450 58.285 ;
        RECT 289.215 58.260 289.425 58.910 ;
        RECT 287.380 57.760 288.450 57.930 ;
        RECT 288.695 57.550 289.000 58.010 ;
        RECT 289.170 57.730 289.425 58.260 ;
        RECT 289.600 59.025 289.870 59.930 ;
        RECT 290.040 59.340 290.370 60.100 ;
        RECT 290.550 59.170 290.720 59.930 ;
        RECT 289.600 58.225 289.770 59.025 ;
        RECT 290.055 59.000 290.720 59.170 ;
        RECT 290.980 59.010 294.490 60.100 ;
        RECT 290.055 58.855 290.225 59.000 ;
        RECT 289.940 58.525 290.225 58.855 ;
        RECT 290.055 58.270 290.225 58.525 ;
        RECT 290.460 58.450 290.790 58.820 ;
        RECT 290.980 58.320 292.630 58.840 ;
        RECT 292.800 58.490 294.490 59.010 ;
        RECT 294.665 58.960 295.000 59.930 ;
        RECT 295.170 58.960 295.340 60.100 ;
        RECT 295.510 59.760 297.540 59.930 ;
        RECT 289.600 57.720 289.860 58.225 ;
        RECT 290.055 58.100 290.720 58.270 ;
        RECT 290.040 57.550 290.370 57.930 ;
        RECT 290.550 57.720 290.720 58.100 ;
        RECT 290.980 57.550 294.490 58.320 ;
        RECT 294.665 58.290 294.835 58.960 ;
        RECT 295.510 58.790 295.680 59.760 ;
        RECT 295.005 58.460 295.260 58.790 ;
        RECT 295.485 58.460 295.680 58.790 ;
        RECT 295.850 59.420 296.975 59.590 ;
        RECT 295.090 58.290 295.260 58.460 ;
        RECT 295.850 58.290 296.020 59.420 ;
        RECT 294.665 57.720 294.920 58.290 ;
        RECT 295.090 58.120 296.020 58.290 ;
        RECT 296.190 59.080 297.200 59.250 ;
        RECT 296.190 58.280 296.360 59.080 ;
        RECT 296.565 58.400 296.840 58.880 ;
        RECT 296.560 58.230 296.840 58.400 ;
        RECT 295.845 58.085 296.020 58.120 ;
        RECT 295.090 57.550 295.420 57.950 ;
        RECT 295.845 57.720 296.375 58.085 ;
        RECT 296.565 57.720 296.840 58.230 ;
        RECT 297.010 57.720 297.200 59.080 ;
        RECT 297.370 59.095 297.540 59.760 ;
        RECT 297.710 59.340 297.880 60.100 ;
        RECT 298.115 59.340 298.630 59.750 ;
        RECT 297.370 58.905 298.120 59.095 ;
        RECT 298.290 58.530 298.630 59.340 ;
        RECT 297.400 58.360 298.630 58.530 ;
        RECT 298.800 59.025 299.070 59.930 ;
        RECT 299.240 59.340 299.570 60.100 ;
        RECT 299.750 59.170 299.920 59.930 ;
        RECT 297.380 57.550 297.890 58.085 ;
        RECT 298.110 57.755 298.355 58.360 ;
        RECT 298.800 58.225 298.970 59.025 ;
        RECT 299.255 59.000 299.920 59.170 ;
        RECT 300.180 59.010 303.690 60.100 ;
        RECT 299.255 58.855 299.425 59.000 ;
        RECT 299.140 58.525 299.425 58.855 ;
        RECT 299.255 58.270 299.425 58.525 ;
        RECT 299.660 58.450 299.990 58.820 ;
        RECT 300.180 58.320 301.830 58.840 ;
        RECT 302.000 58.490 303.690 59.010 ;
        RECT 303.860 58.935 304.150 60.100 ;
        RECT 304.320 59.665 309.665 60.100 ;
        RECT 298.800 57.720 299.060 58.225 ;
        RECT 299.255 58.100 299.920 58.270 ;
        RECT 299.240 57.550 299.570 57.930 ;
        RECT 299.750 57.720 299.920 58.100 ;
        RECT 300.180 57.550 303.690 58.320 ;
        RECT 303.860 57.550 304.150 58.275 ;
        RECT 305.905 58.095 306.245 58.925 ;
        RECT 307.725 58.415 308.075 59.665 ;
        RECT 309.840 59.010 311.050 60.100 ;
        RECT 309.840 58.470 310.360 59.010 ;
        RECT 310.530 58.300 311.050 58.840 ;
        RECT 304.320 57.550 309.665 58.095 ;
        RECT 309.840 57.550 311.050 58.300 ;
        RECT 162.095 57.380 311.135 57.550 ;
        RECT 162.180 56.630 163.390 57.380 ;
        RECT 162.180 56.090 162.700 56.630 ;
        RECT 163.560 56.610 166.150 57.380 ;
        RECT 166.320 56.705 166.580 57.210 ;
        RECT 166.760 57.000 167.090 57.380 ;
        RECT 167.270 56.830 167.440 57.210 ;
        RECT 162.870 55.920 163.390 56.460 ;
        RECT 163.560 56.090 164.770 56.610 ;
        RECT 164.940 55.920 166.150 56.440 ;
        RECT 162.180 54.830 163.390 55.920 ;
        RECT 163.560 54.830 166.150 55.920 ;
        RECT 166.320 55.905 166.490 56.705 ;
        RECT 166.775 56.660 167.440 56.830 ;
        RECT 167.705 56.830 167.960 57.120 ;
        RECT 168.130 57.000 168.460 57.380 ;
        RECT 167.705 56.660 168.455 56.830 ;
        RECT 166.775 56.405 166.945 56.660 ;
        RECT 166.660 56.075 166.945 56.405 ;
        RECT 167.180 56.110 167.510 56.480 ;
        RECT 166.775 55.930 166.945 56.075 ;
        RECT 166.320 55.000 166.590 55.905 ;
        RECT 166.775 55.760 167.440 55.930 ;
        RECT 167.705 55.840 168.055 56.490 ;
        RECT 166.760 54.830 167.090 55.590 ;
        RECT 167.270 55.000 167.440 55.760 ;
        RECT 168.225 55.670 168.455 56.660 ;
        RECT 167.705 55.500 168.455 55.670 ;
        RECT 167.705 55.000 167.960 55.500 ;
        RECT 168.130 54.830 168.460 55.330 ;
        RECT 168.630 55.000 168.800 57.120 ;
        RECT 169.160 57.020 169.490 57.380 ;
        RECT 169.660 56.990 170.155 57.160 ;
        RECT 170.360 56.990 171.215 57.160 ;
        RECT 169.030 55.800 169.490 56.850 ;
        RECT 168.970 55.015 169.295 55.800 ;
        RECT 169.660 55.630 169.830 56.990 ;
        RECT 170.000 56.080 170.350 56.700 ;
        RECT 170.520 56.480 170.875 56.700 ;
        RECT 170.520 55.890 170.690 56.480 ;
        RECT 171.045 56.280 171.215 56.990 ;
        RECT 172.090 56.920 172.420 57.380 ;
        RECT 172.630 57.020 172.980 57.190 ;
        RECT 171.420 56.450 172.210 56.700 ;
        RECT 172.630 56.630 172.890 57.020 ;
        RECT 173.200 56.930 174.150 57.210 ;
        RECT 174.320 56.940 174.510 57.380 ;
        RECT 174.680 57.000 175.750 57.170 ;
        RECT 172.380 56.280 172.550 56.460 ;
        RECT 169.660 55.460 170.055 55.630 ;
        RECT 170.225 55.500 170.690 55.890 ;
        RECT 170.860 56.110 172.550 56.280 ;
        RECT 169.885 55.330 170.055 55.460 ;
        RECT 170.860 55.330 171.030 56.110 ;
        RECT 172.720 55.940 172.890 56.630 ;
        RECT 171.390 55.770 172.890 55.940 ;
        RECT 173.080 55.970 173.290 56.760 ;
        RECT 173.460 56.140 173.810 56.760 ;
        RECT 173.980 56.150 174.150 56.930 ;
        RECT 174.680 56.770 174.850 57.000 ;
        RECT 174.320 56.600 174.850 56.770 ;
        RECT 174.320 56.320 174.540 56.600 ;
        RECT 175.020 56.430 175.260 56.830 ;
        RECT 173.980 55.980 174.385 56.150 ;
        RECT 174.720 56.060 175.260 56.430 ;
        RECT 175.430 56.645 175.750 57.000 ;
        RECT 175.995 56.920 176.300 57.380 ;
        RECT 176.470 56.670 176.720 57.200 ;
        RECT 175.430 56.470 175.755 56.645 ;
        RECT 175.430 56.170 176.345 56.470 ;
        RECT 175.605 56.140 176.345 56.170 ;
        RECT 173.080 55.810 173.755 55.970 ;
        RECT 174.215 55.890 174.385 55.980 ;
        RECT 173.080 55.800 174.045 55.810 ;
        RECT 172.720 55.630 172.890 55.770 ;
        RECT 169.465 54.830 169.715 55.290 ;
        RECT 169.885 55.000 170.135 55.330 ;
        RECT 170.350 55.000 171.030 55.330 ;
        RECT 171.200 55.430 172.275 55.600 ;
        RECT 172.720 55.460 173.280 55.630 ;
        RECT 173.585 55.510 174.045 55.800 ;
        RECT 174.215 55.720 175.435 55.890 ;
        RECT 171.200 55.090 171.370 55.430 ;
        RECT 171.605 54.830 171.935 55.260 ;
        RECT 172.105 55.090 172.275 55.430 ;
        RECT 172.570 54.830 172.940 55.290 ;
        RECT 173.110 55.000 173.280 55.460 ;
        RECT 174.215 55.340 174.385 55.720 ;
        RECT 175.605 55.550 175.775 56.140 ;
        RECT 176.515 56.020 176.720 56.670 ;
        RECT 176.890 56.625 177.140 57.380 ;
        RECT 177.365 56.830 177.620 57.120 ;
        RECT 177.790 57.000 178.120 57.380 ;
        RECT 177.365 56.660 178.115 56.830 ;
        RECT 173.515 55.000 174.385 55.340 ;
        RECT 174.975 55.380 175.775 55.550 ;
        RECT 174.555 54.830 174.805 55.290 ;
        RECT 174.975 55.090 175.145 55.380 ;
        RECT 175.325 54.830 175.655 55.210 ;
        RECT 175.995 54.830 176.300 55.970 ;
        RECT 176.470 55.140 176.720 56.020 ;
        RECT 176.890 54.830 177.140 55.970 ;
        RECT 177.365 55.840 177.715 56.490 ;
        RECT 177.885 55.670 178.115 56.660 ;
        RECT 177.365 55.500 178.115 55.670 ;
        RECT 177.365 55.000 177.620 55.500 ;
        RECT 177.790 54.830 178.120 55.330 ;
        RECT 178.290 55.000 178.460 57.120 ;
        RECT 178.820 57.020 179.150 57.380 ;
        RECT 179.320 56.990 179.815 57.160 ;
        RECT 180.020 56.990 180.875 57.160 ;
        RECT 178.690 55.800 179.150 56.850 ;
        RECT 178.630 55.015 178.955 55.800 ;
        RECT 179.320 55.630 179.490 56.990 ;
        RECT 179.660 56.080 180.010 56.700 ;
        RECT 180.180 56.480 180.535 56.700 ;
        RECT 180.180 55.890 180.350 56.480 ;
        RECT 180.705 56.280 180.875 56.990 ;
        RECT 181.750 56.920 182.080 57.380 ;
        RECT 182.290 57.020 182.640 57.190 ;
        RECT 181.080 56.450 181.870 56.700 ;
        RECT 182.290 56.630 182.550 57.020 ;
        RECT 182.860 56.930 183.810 57.210 ;
        RECT 183.980 56.940 184.170 57.380 ;
        RECT 184.340 57.000 185.410 57.170 ;
        RECT 182.040 56.280 182.210 56.460 ;
        RECT 179.320 55.460 179.715 55.630 ;
        RECT 179.885 55.500 180.350 55.890 ;
        RECT 180.520 56.110 182.210 56.280 ;
        RECT 179.545 55.330 179.715 55.460 ;
        RECT 180.520 55.330 180.690 56.110 ;
        RECT 182.380 55.940 182.550 56.630 ;
        RECT 181.050 55.770 182.550 55.940 ;
        RECT 182.740 55.970 182.950 56.760 ;
        RECT 183.120 56.140 183.470 56.760 ;
        RECT 183.640 56.150 183.810 56.930 ;
        RECT 184.340 56.770 184.510 57.000 ;
        RECT 183.980 56.600 184.510 56.770 ;
        RECT 183.980 56.320 184.200 56.600 ;
        RECT 184.680 56.430 184.920 56.830 ;
        RECT 183.640 55.980 184.045 56.150 ;
        RECT 184.380 56.060 184.920 56.430 ;
        RECT 185.090 56.645 185.410 57.000 ;
        RECT 185.090 56.390 185.415 56.645 ;
        RECT 185.610 56.570 185.780 57.380 ;
        RECT 185.950 56.730 186.280 57.210 ;
        RECT 186.450 56.910 186.620 57.380 ;
        RECT 186.790 56.730 187.120 57.210 ;
        RECT 187.290 56.910 187.460 57.380 ;
        RECT 185.950 56.560 187.715 56.730 ;
        RECT 187.940 56.655 188.230 57.380 ;
        RECT 185.090 56.180 187.120 56.390 ;
        RECT 185.090 56.170 185.435 56.180 ;
        RECT 182.740 55.810 183.415 55.970 ;
        RECT 183.875 55.890 184.045 55.980 ;
        RECT 182.740 55.800 183.705 55.810 ;
        RECT 182.380 55.630 182.550 55.770 ;
        RECT 179.125 54.830 179.375 55.290 ;
        RECT 179.545 55.000 179.795 55.330 ;
        RECT 180.010 55.000 180.690 55.330 ;
        RECT 180.860 55.430 181.935 55.600 ;
        RECT 182.380 55.460 182.940 55.630 ;
        RECT 183.245 55.510 183.705 55.800 ;
        RECT 183.875 55.720 185.095 55.890 ;
        RECT 180.860 55.090 181.030 55.430 ;
        RECT 181.265 54.830 181.595 55.260 ;
        RECT 181.765 55.090 181.935 55.430 ;
        RECT 182.230 54.830 182.600 55.290 ;
        RECT 182.770 55.000 182.940 55.460 ;
        RECT 183.875 55.340 184.045 55.720 ;
        RECT 185.265 55.550 185.435 56.170 ;
        RECT 187.305 56.010 187.715 56.560 ;
        RECT 188.400 56.610 190.990 57.380 ;
        RECT 191.165 56.830 191.420 57.120 ;
        RECT 191.590 57.000 191.920 57.380 ;
        RECT 191.165 56.660 191.915 56.830 ;
        RECT 188.400 56.090 189.610 56.610 ;
        RECT 183.175 55.000 184.045 55.340 ;
        RECT 184.635 55.380 185.435 55.550 ;
        RECT 184.215 54.830 184.465 55.290 ;
        RECT 184.635 55.090 184.805 55.380 ;
        RECT 184.985 54.830 185.315 55.210 ;
        RECT 185.610 54.830 185.780 55.890 ;
        RECT 185.990 55.840 187.715 56.010 ;
        RECT 185.990 55.000 186.280 55.840 ;
        RECT 186.450 54.830 186.620 55.670 ;
        RECT 186.830 55.000 187.080 55.840 ;
        RECT 187.290 54.830 187.460 55.670 ;
        RECT 187.940 54.830 188.230 55.995 ;
        RECT 189.780 55.920 190.990 56.440 ;
        RECT 188.400 54.830 190.990 55.920 ;
        RECT 191.165 55.840 191.515 56.490 ;
        RECT 191.685 55.670 191.915 56.660 ;
        RECT 191.165 55.500 191.915 55.670 ;
        RECT 191.165 55.000 191.420 55.500 ;
        RECT 191.590 54.830 191.920 55.330 ;
        RECT 192.090 55.000 192.260 57.120 ;
        RECT 192.620 57.020 192.950 57.380 ;
        RECT 193.120 56.990 193.615 57.160 ;
        RECT 193.820 56.990 194.675 57.160 ;
        RECT 192.490 55.800 192.950 56.850 ;
        RECT 192.430 55.015 192.755 55.800 ;
        RECT 193.120 55.630 193.290 56.990 ;
        RECT 193.460 56.080 193.810 56.700 ;
        RECT 193.980 56.480 194.335 56.700 ;
        RECT 193.980 55.890 194.150 56.480 ;
        RECT 194.505 56.280 194.675 56.990 ;
        RECT 195.550 56.920 195.880 57.380 ;
        RECT 196.090 57.020 196.440 57.190 ;
        RECT 194.880 56.450 195.670 56.700 ;
        RECT 196.090 56.630 196.350 57.020 ;
        RECT 196.660 56.930 197.610 57.210 ;
        RECT 197.780 56.940 197.970 57.380 ;
        RECT 198.140 57.000 199.210 57.170 ;
        RECT 195.840 56.280 196.010 56.460 ;
        RECT 193.120 55.460 193.515 55.630 ;
        RECT 193.685 55.500 194.150 55.890 ;
        RECT 194.320 56.110 196.010 56.280 ;
        RECT 193.345 55.330 193.515 55.460 ;
        RECT 194.320 55.330 194.490 56.110 ;
        RECT 196.180 55.940 196.350 56.630 ;
        RECT 194.850 55.770 196.350 55.940 ;
        RECT 196.540 55.970 196.750 56.760 ;
        RECT 196.920 56.140 197.270 56.760 ;
        RECT 197.440 56.150 197.610 56.930 ;
        RECT 198.140 56.770 198.310 57.000 ;
        RECT 197.780 56.600 198.310 56.770 ;
        RECT 197.780 56.320 198.000 56.600 ;
        RECT 198.480 56.430 198.720 56.830 ;
        RECT 197.440 55.980 197.845 56.150 ;
        RECT 198.180 56.060 198.720 56.430 ;
        RECT 198.890 56.645 199.210 57.000 ;
        RECT 199.455 56.920 199.760 57.380 ;
        RECT 199.930 56.670 200.180 57.200 ;
        RECT 198.890 56.470 199.215 56.645 ;
        RECT 198.890 56.170 199.805 56.470 ;
        RECT 199.065 56.140 199.805 56.170 ;
        RECT 196.540 55.810 197.215 55.970 ;
        RECT 197.675 55.890 197.845 55.980 ;
        RECT 196.540 55.800 197.505 55.810 ;
        RECT 196.180 55.630 196.350 55.770 ;
        RECT 192.925 54.830 193.175 55.290 ;
        RECT 193.345 55.000 193.595 55.330 ;
        RECT 193.810 55.000 194.490 55.330 ;
        RECT 194.660 55.430 195.735 55.600 ;
        RECT 196.180 55.460 196.740 55.630 ;
        RECT 197.045 55.510 197.505 55.800 ;
        RECT 197.675 55.720 198.895 55.890 ;
        RECT 194.660 55.090 194.830 55.430 ;
        RECT 195.065 54.830 195.395 55.260 ;
        RECT 195.565 55.090 195.735 55.430 ;
        RECT 196.030 54.830 196.400 55.290 ;
        RECT 196.570 55.000 196.740 55.460 ;
        RECT 197.675 55.340 197.845 55.720 ;
        RECT 199.065 55.550 199.235 56.140 ;
        RECT 199.975 56.020 200.180 56.670 ;
        RECT 200.350 56.625 200.600 57.380 ;
        RECT 200.820 56.610 202.490 57.380 ;
        RECT 202.665 56.640 202.920 57.210 ;
        RECT 203.090 56.980 203.420 57.380 ;
        RECT 203.845 56.845 204.375 57.210 ;
        RECT 204.565 57.040 204.840 57.210 ;
        RECT 204.560 56.870 204.840 57.040 ;
        RECT 203.845 56.810 204.020 56.845 ;
        RECT 203.090 56.640 204.020 56.810 ;
        RECT 200.820 56.090 201.570 56.610 ;
        RECT 196.975 55.000 197.845 55.340 ;
        RECT 198.435 55.380 199.235 55.550 ;
        RECT 198.015 54.830 198.265 55.290 ;
        RECT 198.435 55.090 198.605 55.380 ;
        RECT 198.785 54.830 199.115 55.210 ;
        RECT 199.455 54.830 199.760 55.970 ;
        RECT 199.930 55.140 200.180 56.020 ;
        RECT 200.350 54.830 200.600 55.970 ;
        RECT 201.740 55.920 202.490 56.440 ;
        RECT 200.820 54.830 202.490 55.920 ;
        RECT 202.665 55.970 202.835 56.640 ;
        RECT 203.090 56.470 203.260 56.640 ;
        RECT 203.005 56.140 203.260 56.470 ;
        RECT 203.485 56.140 203.680 56.470 ;
        RECT 202.665 55.000 203.000 55.970 ;
        RECT 203.170 54.830 203.340 55.970 ;
        RECT 203.510 55.170 203.680 56.140 ;
        RECT 203.850 55.510 204.020 56.640 ;
        RECT 204.190 55.850 204.360 56.650 ;
        RECT 204.565 56.050 204.840 56.870 ;
        RECT 205.010 55.850 205.200 57.210 ;
        RECT 205.380 56.845 205.890 57.380 ;
        RECT 206.110 56.570 206.355 57.175 ;
        RECT 206.805 57.125 207.140 57.170 ;
        RECT 206.800 56.660 207.140 57.125 ;
        RECT 207.310 57.000 207.640 57.380 ;
        RECT 205.400 56.400 206.630 56.570 ;
        RECT 204.190 55.680 205.200 55.850 ;
        RECT 205.370 55.835 206.120 56.025 ;
        RECT 203.850 55.340 204.975 55.510 ;
        RECT 205.370 55.170 205.540 55.835 ;
        RECT 206.290 55.590 206.630 56.400 ;
        RECT 203.510 55.000 205.540 55.170 ;
        RECT 205.710 54.830 205.880 55.590 ;
        RECT 206.115 55.180 206.630 55.590 ;
        RECT 206.800 55.970 206.970 56.660 ;
        RECT 207.140 56.140 207.400 56.470 ;
        RECT 206.800 55.000 207.060 55.970 ;
        RECT 207.230 55.590 207.400 56.140 ;
        RECT 207.570 55.770 207.910 56.800 ;
        RECT 208.100 56.360 208.370 57.045 ;
        RECT 208.100 56.190 208.410 56.360 ;
        RECT 208.100 55.770 208.370 56.190 ;
        RECT 208.595 55.770 208.875 57.045 ;
        RECT 209.075 56.880 209.305 57.210 ;
        RECT 209.550 57.000 209.880 57.380 ;
        RECT 209.075 55.590 209.245 56.880 ;
        RECT 210.050 56.810 210.225 57.210 ;
        RECT 209.595 56.640 210.225 56.810 ;
        RECT 209.595 56.470 209.765 56.640 ;
        RECT 210.500 56.580 210.740 57.380 ;
        RECT 209.415 56.140 209.765 56.470 ;
        RECT 207.230 55.420 209.245 55.590 ;
        RECT 209.595 55.620 209.765 56.140 ;
        RECT 209.945 55.790 210.310 56.470 ;
        RECT 209.595 55.450 210.225 55.620 ;
        RECT 207.255 54.830 207.585 55.240 ;
        RECT 207.785 55.000 207.955 55.420 ;
        RECT 208.170 54.830 208.840 55.240 ;
        RECT 209.075 55.000 209.245 55.420 ;
        RECT 209.550 54.830 209.880 55.270 ;
        RECT 210.050 55.000 210.225 55.450 ;
        RECT 210.485 54.830 210.740 55.830 ;
        RECT 210.925 55.000 211.170 57.210 ;
        RECT 211.340 57.000 211.670 57.380 ;
        RECT 211.860 56.830 212.190 57.210 ;
        RECT 212.740 57.000 213.070 57.380 ;
        RECT 211.340 56.625 212.190 56.830 ;
        RECT 212.360 56.830 212.570 57.000 ;
        RECT 213.240 56.830 213.515 56.970 ;
        RECT 212.360 56.640 213.515 56.830 ;
        RECT 213.700 56.655 213.990 57.380 ;
        RECT 214.620 57.000 214.950 57.380 ;
        RECT 214.175 56.830 214.450 56.970 ;
        RECT 215.120 56.830 215.330 57.000 ;
        RECT 214.175 56.640 215.330 56.830 ;
        RECT 215.500 56.830 215.830 57.210 ;
        RECT 216.020 57.000 216.350 57.380 ;
        RECT 215.500 56.625 216.350 56.830 ;
        RECT 211.340 56.135 211.670 56.625 ;
        RECT 211.500 55.680 211.670 56.135 ;
        RECT 211.840 55.850 212.250 56.455 ;
        RECT 212.420 56.065 213.005 56.440 ;
        RECT 212.800 55.680 213.005 56.065 ;
        RECT 213.260 56.015 213.520 56.470 ;
        RECT 214.170 56.015 214.430 56.470 ;
        RECT 214.685 56.065 215.270 56.440 ;
        RECT 214.685 56.020 214.890 56.065 ;
        RECT 211.500 55.460 212.620 55.680 ;
        RECT 212.800 55.510 213.010 55.680 ;
        RECT 212.800 55.480 213.005 55.510 ;
        RECT 211.340 54.830 212.190 55.280 ;
        RECT 212.360 55.000 212.620 55.460 ;
        RECT 213.190 54.830 213.515 55.815 ;
        RECT 213.700 54.830 213.990 55.995 ;
        RECT 214.680 55.850 214.890 56.020 ;
        RECT 215.440 55.850 215.850 56.455 ;
        RECT 216.020 56.135 216.350 56.625 ;
        RECT 214.175 54.830 214.500 55.815 ;
        RECT 214.685 55.480 214.890 55.850 ;
        RECT 216.020 55.680 216.190 56.135 ;
        RECT 215.070 55.460 216.190 55.680 ;
        RECT 215.070 55.000 215.330 55.460 ;
        RECT 215.500 54.830 216.350 55.280 ;
        RECT 216.520 55.000 216.765 57.210 ;
        RECT 216.950 56.580 217.190 57.380 ;
        RECT 217.380 56.835 222.725 57.380 ;
        RECT 218.965 56.005 219.305 56.835 ;
        RECT 223.910 56.830 224.080 57.210 ;
        RECT 224.295 57.000 224.625 57.380 ;
        RECT 223.910 56.660 224.625 56.830 ;
        RECT 216.950 54.830 217.205 55.830 ;
        RECT 220.785 55.265 221.135 56.515 ;
        RECT 223.820 56.110 224.175 56.480 ;
        RECT 224.455 56.470 224.625 56.660 ;
        RECT 224.795 56.635 225.050 57.210 ;
        RECT 224.455 56.140 224.710 56.470 ;
        RECT 224.455 55.930 224.625 56.140 ;
        RECT 223.910 55.760 224.625 55.930 ;
        RECT 224.880 55.905 225.050 56.635 ;
        RECT 225.225 56.540 225.485 57.380 ;
        RECT 217.380 54.830 222.725 55.265 ;
        RECT 223.910 55.000 224.080 55.760 ;
        RECT 224.295 54.830 224.625 55.590 ;
        RECT 224.795 55.000 225.050 55.905 ;
        RECT 225.225 54.830 225.485 55.980 ;
        RECT 225.670 55.000 225.930 57.210 ;
        RECT 226.110 56.900 226.420 57.380 ;
        RECT 226.600 56.730 226.940 57.210 ;
        RECT 226.270 56.560 226.940 56.730 ;
        RECT 226.270 56.470 226.440 56.560 ;
        RECT 226.100 56.140 226.440 56.470 ;
        RECT 227.110 56.390 227.320 57.075 ;
        RECT 226.840 56.140 227.320 56.390 ;
        RECT 227.500 56.140 227.770 57.075 ;
        RECT 228.020 56.470 228.265 57.075 ;
        RECT 228.445 56.760 228.735 57.210 ;
        RECT 228.905 56.930 229.195 57.380 ;
        RECT 229.365 56.760 229.630 57.210 ;
        RECT 228.445 56.590 229.630 56.760 ;
        RECT 229.960 56.560 230.250 57.380 ;
        RECT 230.420 56.650 230.750 57.210 ;
        RECT 228.020 56.140 228.280 56.470 ;
        RECT 230.500 56.390 230.750 56.650 ;
        RECT 230.930 56.560 231.220 57.380 ;
        RECT 231.390 56.740 231.720 57.210 ;
        RECT 231.890 56.910 232.060 57.380 ;
        RECT 232.230 56.740 232.560 57.210 ;
        RECT 232.730 56.910 232.900 57.380 ;
        RECT 233.070 56.740 233.400 57.210 ;
        RECT 233.570 56.910 233.740 57.380 ;
        RECT 233.910 56.740 234.240 57.210 ;
        RECT 231.390 56.560 234.240 56.740 ;
        RECT 234.410 56.560 234.690 57.380 ;
        RECT 234.860 56.610 238.370 57.380 ;
        RECT 239.460 56.655 239.750 57.380 ;
        RECT 228.625 56.140 229.110 56.390 ;
        RECT 226.270 55.970 226.440 56.140 ;
        RECT 226.270 55.800 228.755 55.970 ;
        RECT 226.100 54.830 226.910 55.630 ;
        RECT 227.080 55.000 227.410 55.800 ;
        RECT 227.595 54.830 228.335 55.630 ;
        RECT 228.505 55.000 228.755 55.800 ;
        RECT 228.925 55.050 229.110 56.140 ;
        RECT 229.280 55.805 229.610 56.390 ;
        RECT 229.800 56.145 230.330 56.390 ;
        RECT 230.500 56.190 231.980 56.390 ;
        RECT 229.305 54.830 229.630 55.630 ;
        RECT 229.845 54.830 230.250 55.970 ;
        RECT 230.500 55.890 230.750 56.190 ;
        RECT 232.150 56.020 232.480 56.560 ;
        RECT 232.975 56.190 234.415 56.390 ;
        RECT 234.860 56.090 236.510 56.610 ;
        RECT 239.920 56.580 240.260 57.210 ;
        RECT 240.430 56.580 240.680 57.380 ;
        RECT 240.870 56.730 241.200 57.210 ;
        RECT 241.370 56.920 241.595 57.380 ;
        RECT 241.765 56.730 242.095 57.210 ;
        RECT 230.420 55.000 230.750 55.890 ;
        RECT 230.920 55.170 231.300 55.890 ;
        RECT 231.470 55.720 232.480 56.020 ;
        RECT 231.470 55.340 231.640 55.720 ;
        RECT 231.810 55.170 232.140 55.530 ;
        RECT 232.310 55.340 232.480 55.720 ;
        RECT 232.650 55.800 234.690 56.010 ;
        RECT 236.680 55.920 238.370 56.440 ;
        RECT 232.650 55.170 232.980 55.800 ;
        RECT 230.920 55.000 232.980 55.170 ;
        RECT 233.150 54.830 233.400 55.630 ;
        RECT 233.570 55.000 233.740 55.800 ;
        RECT 233.910 54.830 234.240 55.630 ;
        RECT 234.410 55.000 234.690 55.800 ;
        RECT 234.860 54.830 238.370 55.920 ;
        RECT 239.460 54.830 239.750 55.995 ;
        RECT 239.920 55.970 240.095 56.580 ;
        RECT 240.870 56.560 242.095 56.730 ;
        RECT 242.725 56.600 243.225 57.210 ;
        RECT 243.600 56.630 244.810 57.380 ;
        RECT 244.995 56.810 245.250 57.160 ;
        RECT 245.420 56.980 245.750 57.380 ;
        RECT 245.920 56.810 246.090 57.160 ;
        RECT 246.260 56.980 246.640 57.380 ;
        RECT 244.995 56.640 246.660 56.810 ;
        RECT 246.830 56.705 247.105 57.050 ;
        RECT 240.265 56.220 240.960 56.390 ;
        RECT 240.790 55.970 240.960 56.220 ;
        RECT 241.135 56.190 241.555 56.390 ;
        RECT 241.725 56.190 242.055 56.390 ;
        RECT 242.225 56.190 242.555 56.390 ;
        RECT 242.725 55.970 242.895 56.600 ;
        RECT 243.080 56.140 243.430 56.390 ;
        RECT 243.600 56.090 244.120 56.630 ;
        RECT 246.490 56.470 246.660 56.640 ;
        RECT 239.920 55.000 240.260 55.970 ;
        RECT 240.430 54.830 240.600 55.970 ;
        RECT 240.790 55.800 243.225 55.970 ;
        RECT 244.290 55.920 244.810 56.460 ;
        RECT 244.980 56.140 245.325 56.470 ;
        RECT 245.495 56.140 246.320 56.470 ;
        RECT 246.490 56.140 246.765 56.470 ;
        RECT 240.870 54.830 241.120 55.630 ;
        RECT 241.765 55.000 242.095 55.800 ;
        RECT 242.395 54.830 242.725 55.630 ;
        RECT 242.895 55.000 243.225 55.800 ;
        RECT 243.600 54.830 244.810 55.920 ;
        RECT 245.000 55.680 245.325 55.970 ;
        RECT 245.495 55.850 245.690 56.140 ;
        RECT 246.490 55.970 246.660 56.140 ;
        RECT 246.935 55.970 247.105 56.705 ;
        RECT 247.760 56.750 248.090 57.210 ;
        RECT 248.270 56.920 248.440 57.380 ;
        RECT 248.620 56.750 248.950 57.210 ;
        RECT 249.180 56.920 249.350 57.380 ;
        RECT 249.590 57.040 250.780 57.210 ;
        RECT 249.590 56.750 249.920 57.040 ;
        RECT 250.470 56.870 250.780 57.040 ;
        RECT 247.760 56.580 249.920 56.750 ;
        RECT 246.000 55.800 246.660 55.970 ;
        RECT 246.000 55.680 246.170 55.800 ;
        RECT 245.000 55.510 246.170 55.680 ;
        RECT 244.980 55.050 246.170 55.340 ;
        RECT 246.340 54.830 246.620 55.630 ;
        RECT 246.830 55.000 247.105 55.970 ;
        RECT 247.775 56.020 248.105 56.410 ;
        RECT 248.275 56.190 249.075 56.390 ;
        RECT 249.255 56.020 249.750 56.390 ;
        RECT 247.775 55.850 249.750 56.020 ;
        RECT 250.090 55.680 250.300 56.870 ;
        RECT 250.960 56.760 251.225 57.210 ;
        RECT 251.395 56.930 251.685 57.380 ;
        RECT 251.855 56.760 252.145 57.210 ;
        RECT 250.470 56.065 250.785 56.700 ;
        RECT 250.960 56.590 252.145 56.760 ;
        RECT 252.325 56.470 252.570 57.075 ;
        RECT 247.760 54.830 248.090 55.680 ;
        RECT 248.260 55.170 248.480 55.680 ;
        RECT 248.650 55.500 250.300 55.680 ;
        RECT 248.650 55.340 248.950 55.500 ;
        RECT 249.180 55.170 249.370 55.330 ;
        RECT 248.260 55.000 249.370 55.170 ;
        RECT 249.565 54.830 249.895 55.290 ;
        RECT 250.065 55.000 250.300 55.500 ;
        RECT 250.470 54.830 250.780 55.895 ;
        RECT 250.980 55.805 251.310 56.390 ;
        RECT 251.480 56.140 251.965 56.390 ;
        RECT 252.310 56.140 252.570 56.470 ;
        RECT 252.820 56.140 253.090 57.075 ;
        RECT 253.270 56.390 253.480 57.075 ;
        RECT 253.650 56.730 253.990 57.210 ;
        RECT 254.170 56.900 254.480 57.380 ;
        RECT 253.650 56.560 254.320 56.730 ;
        RECT 254.150 56.470 254.320 56.560 ;
        RECT 253.270 56.140 253.750 56.390 ;
        RECT 254.150 56.140 254.490 56.470 ;
        RECT 250.960 54.830 251.285 55.630 ;
        RECT 251.480 55.050 251.665 56.140 ;
        RECT 254.150 55.970 254.320 56.140 ;
        RECT 251.835 55.800 254.320 55.970 ;
        RECT 251.835 55.000 252.085 55.800 ;
        RECT 252.255 54.830 252.995 55.630 ;
        RECT 253.180 55.000 253.510 55.800 ;
        RECT 253.680 54.830 254.490 55.630 ;
        RECT 254.660 55.000 254.920 57.210 ;
        RECT 255.100 56.560 255.360 57.380 ;
        RECT 255.530 56.560 255.860 56.980 ;
        RECT 256.040 56.810 256.300 57.210 ;
        RECT 256.470 56.980 256.800 57.380 ;
        RECT 256.970 56.810 257.140 57.160 ;
        RECT 257.310 56.980 257.685 57.380 ;
        RECT 256.040 56.640 257.705 56.810 ;
        RECT 257.875 56.705 258.150 57.050 ;
        RECT 255.610 56.470 255.860 56.560 ;
        RECT 257.535 56.470 257.705 56.640 ;
        RECT 255.105 56.140 255.440 56.390 ;
        RECT 255.610 56.140 256.325 56.470 ;
        RECT 256.540 56.140 257.365 56.470 ;
        RECT 257.535 56.140 257.810 56.470 ;
        RECT 255.100 54.830 255.360 55.970 ;
        RECT 255.610 55.580 255.780 56.140 ;
        RECT 256.040 55.680 256.370 55.970 ;
        RECT 256.540 55.850 256.785 56.140 ;
        RECT 257.535 55.970 257.705 56.140 ;
        RECT 257.980 55.970 258.150 56.705 ;
        RECT 258.320 56.610 260.910 57.380 ;
        RECT 261.540 56.640 262.050 57.210 ;
        RECT 262.220 56.820 262.390 57.380 ;
        RECT 262.595 56.810 262.925 57.210 ;
        RECT 263.100 56.980 263.430 57.380 ;
        RECT 263.665 57.000 265.050 57.210 ;
        RECT 263.665 56.810 263.995 57.000 ;
        RECT 262.595 56.640 263.995 56.810 ;
        RECT 264.165 56.640 264.590 56.830 ;
        RECT 264.760 56.730 265.050 57.000 ;
        RECT 265.220 56.655 265.510 57.380 ;
        RECT 265.780 56.730 266.110 57.210 ;
        RECT 266.280 56.920 266.610 57.380 ;
        RECT 266.825 56.730 267.155 57.210 ;
        RECT 267.355 56.920 267.685 57.380 ;
        RECT 267.910 56.730 268.080 57.050 ;
        RECT 258.320 56.090 259.530 56.610 ;
        RECT 257.045 55.800 257.705 55.970 ;
        RECT 257.045 55.680 257.215 55.800 ;
        RECT 256.040 55.510 257.215 55.680 ;
        RECT 255.600 55.010 257.215 55.340 ;
        RECT 257.385 54.830 257.665 55.630 ;
        RECT 257.875 55.000 258.150 55.970 ;
        RECT 259.700 55.920 260.910 56.440 ;
        RECT 258.320 54.830 260.910 55.920 ;
        RECT 261.540 55.970 261.715 56.640 ;
        RECT 261.900 56.390 262.090 56.470 ;
        RECT 262.460 56.390 262.630 56.470 ;
        RECT 261.900 56.140 262.265 56.390 ;
        RECT 262.460 56.140 262.710 56.390 ;
        RECT 262.920 56.140 263.265 56.470 ;
        RECT 262.095 55.970 262.265 56.140 ;
        RECT 261.540 55.010 261.925 55.970 ;
        RECT 262.095 55.800 262.770 55.970 ;
        RECT 262.140 54.830 262.430 55.630 ;
        RECT 262.600 55.170 262.770 55.800 ;
        RECT 262.940 55.340 263.265 56.140 ;
        RECT 263.435 55.805 263.710 56.470 ;
        RECT 263.895 55.805 264.250 56.470 ;
        RECT 264.420 55.630 264.590 56.640 ;
        RECT 265.780 56.560 268.080 56.730 ;
        RECT 268.250 56.750 268.580 57.195 ;
        RECT 268.850 56.920 269.020 57.380 ;
        RECT 268.250 56.560 269.000 56.750 ;
        RECT 269.310 56.580 269.650 57.210 ;
        RECT 264.775 56.140 265.050 56.470 ;
        RECT 268.630 56.390 269.000 56.560 ;
        RECT 265.740 56.140 266.250 56.390 ;
        RECT 263.635 55.380 264.590 55.630 ;
        RECT 263.635 55.170 263.965 55.380 ;
        RECT 262.600 55.000 263.965 55.170 ;
        RECT 264.760 54.830 265.050 55.970 ;
        RECT 265.220 54.830 265.510 55.995 ;
        RECT 265.800 54.830 266.130 55.950 ;
        RECT 266.460 55.075 266.830 56.390 ;
        RECT 267.000 55.075 267.330 56.390 ;
        RECT 267.540 55.075 267.870 56.390 ;
        RECT 268.040 56.180 268.460 56.390 ;
        RECT 268.630 56.180 269.210 56.390 ;
        RECT 268.630 56.010 268.890 56.180 ;
        RECT 269.380 56.010 269.650 56.580 ;
        RECT 269.820 56.610 271.490 57.380 ;
        RECT 272.125 56.670 272.380 57.200 ;
        RECT 272.550 56.920 272.855 57.380 ;
        RECT 273.100 57.000 274.170 57.170 ;
        RECT 269.820 56.090 270.570 56.610 ;
        RECT 268.140 55.720 268.890 56.010 ;
        RECT 268.140 55.000 268.390 55.720 ;
        RECT 268.560 54.830 268.890 55.550 ;
        RECT 269.125 55.000 269.650 56.010 ;
        RECT 270.740 55.920 271.490 56.440 ;
        RECT 269.820 54.830 271.490 55.920 ;
        RECT 272.125 56.020 272.335 56.670 ;
        RECT 273.100 56.645 273.420 57.000 ;
        RECT 273.095 56.470 273.420 56.645 ;
        RECT 272.505 56.170 273.420 56.470 ;
        RECT 273.590 56.430 273.830 56.830 ;
        RECT 274.000 56.770 274.170 57.000 ;
        RECT 274.340 56.940 274.530 57.380 ;
        RECT 274.700 56.930 275.650 57.210 ;
        RECT 275.870 57.020 276.220 57.190 ;
        RECT 274.000 56.600 274.530 56.770 ;
        RECT 272.505 56.140 273.245 56.170 ;
        RECT 272.125 55.140 272.380 56.020 ;
        RECT 272.550 54.830 272.855 55.970 ;
        RECT 273.075 55.550 273.245 56.140 ;
        RECT 273.590 56.060 274.130 56.430 ;
        RECT 274.310 56.320 274.530 56.600 ;
        RECT 274.700 56.150 274.870 56.930 ;
        RECT 274.465 55.980 274.870 56.150 ;
        RECT 275.040 56.140 275.390 56.760 ;
        RECT 274.465 55.890 274.635 55.980 ;
        RECT 275.560 55.970 275.770 56.760 ;
        RECT 273.415 55.720 274.635 55.890 ;
        RECT 275.095 55.810 275.770 55.970 ;
        RECT 273.075 55.380 273.875 55.550 ;
        RECT 273.195 54.830 273.525 55.210 ;
        RECT 273.705 55.090 273.875 55.380 ;
        RECT 274.465 55.340 274.635 55.720 ;
        RECT 274.805 55.800 275.770 55.810 ;
        RECT 275.960 56.630 276.220 57.020 ;
        RECT 276.430 56.920 276.760 57.380 ;
        RECT 277.635 56.990 278.490 57.160 ;
        RECT 278.695 56.990 279.190 57.160 ;
        RECT 279.360 57.020 279.690 57.380 ;
        RECT 275.960 55.940 276.130 56.630 ;
        RECT 276.300 56.280 276.470 56.460 ;
        RECT 276.640 56.450 277.430 56.700 ;
        RECT 277.635 56.280 277.805 56.990 ;
        RECT 277.975 56.480 278.330 56.700 ;
        RECT 276.300 56.110 277.990 56.280 ;
        RECT 274.805 55.510 275.265 55.800 ;
        RECT 275.960 55.770 277.460 55.940 ;
        RECT 275.960 55.630 276.130 55.770 ;
        RECT 275.570 55.460 276.130 55.630 ;
        RECT 274.045 54.830 274.295 55.290 ;
        RECT 274.465 55.000 275.335 55.340 ;
        RECT 275.570 55.000 275.740 55.460 ;
        RECT 276.575 55.430 277.650 55.600 ;
        RECT 275.910 54.830 276.280 55.290 ;
        RECT 276.575 55.090 276.745 55.430 ;
        RECT 276.915 54.830 277.245 55.260 ;
        RECT 277.480 55.090 277.650 55.430 ;
        RECT 277.820 55.330 277.990 56.110 ;
        RECT 278.160 55.890 278.330 56.480 ;
        RECT 278.500 56.080 278.850 56.700 ;
        RECT 278.160 55.500 278.625 55.890 ;
        RECT 279.020 55.630 279.190 56.990 ;
        RECT 279.360 55.800 279.820 56.850 ;
        RECT 278.795 55.460 279.190 55.630 ;
        RECT 278.795 55.330 278.965 55.460 ;
        RECT 277.820 55.000 278.500 55.330 ;
        RECT 278.715 55.000 278.965 55.330 ;
        RECT 279.135 54.830 279.385 55.290 ;
        RECT 279.555 55.015 279.880 55.800 ;
        RECT 280.050 55.000 280.220 57.120 ;
        RECT 280.390 57.000 280.720 57.380 ;
        RECT 280.890 56.830 281.145 57.120 ;
        RECT 280.395 56.660 281.145 56.830 ;
        RECT 280.395 55.670 280.625 56.660 ;
        RECT 281.370 56.625 281.620 57.380 ;
        RECT 281.790 56.670 282.040 57.200 ;
        RECT 282.210 56.920 282.515 57.380 ;
        RECT 282.760 57.000 283.830 57.170 ;
        RECT 280.795 55.840 281.145 56.490 ;
        RECT 281.790 56.020 281.995 56.670 ;
        RECT 282.760 56.645 283.080 57.000 ;
        RECT 282.755 56.470 283.080 56.645 ;
        RECT 282.165 56.170 283.080 56.470 ;
        RECT 283.250 56.430 283.490 56.830 ;
        RECT 283.660 56.770 283.830 57.000 ;
        RECT 284.000 56.940 284.190 57.380 ;
        RECT 284.360 56.930 285.310 57.210 ;
        RECT 285.530 57.020 285.880 57.190 ;
        RECT 283.660 56.600 284.190 56.770 ;
        RECT 282.165 56.140 282.905 56.170 ;
        RECT 280.395 55.500 281.145 55.670 ;
        RECT 280.390 54.830 280.720 55.330 ;
        RECT 280.890 55.000 281.145 55.500 ;
        RECT 281.370 54.830 281.620 55.970 ;
        RECT 281.790 55.140 282.040 56.020 ;
        RECT 282.210 54.830 282.515 55.970 ;
        RECT 282.735 55.550 282.905 56.140 ;
        RECT 283.250 56.060 283.790 56.430 ;
        RECT 283.970 56.320 284.190 56.600 ;
        RECT 284.360 56.150 284.530 56.930 ;
        RECT 284.125 55.980 284.530 56.150 ;
        RECT 284.700 56.140 285.050 56.760 ;
        RECT 284.125 55.890 284.295 55.980 ;
        RECT 285.220 55.970 285.430 56.760 ;
        RECT 283.075 55.720 284.295 55.890 ;
        RECT 284.755 55.810 285.430 55.970 ;
        RECT 282.735 55.380 283.535 55.550 ;
        RECT 282.855 54.830 283.185 55.210 ;
        RECT 283.365 55.090 283.535 55.380 ;
        RECT 284.125 55.340 284.295 55.720 ;
        RECT 284.465 55.800 285.430 55.810 ;
        RECT 285.620 56.630 285.880 57.020 ;
        RECT 286.090 56.920 286.420 57.380 ;
        RECT 287.295 56.990 288.150 57.160 ;
        RECT 288.355 56.990 288.850 57.160 ;
        RECT 289.020 57.020 289.350 57.380 ;
        RECT 285.620 55.940 285.790 56.630 ;
        RECT 285.960 56.280 286.130 56.460 ;
        RECT 286.300 56.450 287.090 56.700 ;
        RECT 287.295 56.280 287.465 56.990 ;
        RECT 287.635 56.480 287.990 56.700 ;
        RECT 285.960 56.110 287.650 56.280 ;
        RECT 284.465 55.510 284.925 55.800 ;
        RECT 285.620 55.770 287.120 55.940 ;
        RECT 285.620 55.630 285.790 55.770 ;
        RECT 285.230 55.460 285.790 55.630 ;
        RECT 283.705 54.830 283.955 55.290 ;
        RECT 284.125 55.000 284.995 55.340 ;
        RECT 285.230 55.000 285.400 55.460 ;
        RECT 286.235 55.430 287.310 55.600 ;
        RECT 285.570 54.830 285.940 55.290 ;
        RECT 286.235 55.090 286.405 55.430 ;
        RECT 286.575 54.830 286.905 55.260 ;
        RECT 287.140 55.090 287.310 55.430 ;
        RECT 287.480 55.330 287.650 56.110 ;
        RECT 287.820 55.890 287.990 56.480 ;
        RECT 288.160 56.080 288.510 56.700 ;
        RECT 287.820 55.500 288.285 55.890 ;
        RECT 288.680 55.630 288.850 56.990 ;
        RECT 289.020 55.800 289.480 56.850 ;
        RECT 288.455 55.460 288.850 55.630 ;
        RECT 288.455 55.330 288.625 55.460 ;
        RECT 287.480 55.000 288.160 55.330 ;
        RECT 288.375 55.000 288.625 55.330 ;
        RECT 288.795 54.830 289.045 55.290 ;
        RECT 289.215 55.015 289.540 55.800 ;
        RECT 289.710 55.000 289.880 57.120 ;
        RECT 290.050 57.000 290.380 57.380 ;
        RECT 290.550 56.830 290.805 57.120 ;
        RECT 290.055 56.660 290.805 56.830 ;
        RECT 290.055 55.670 290.285 56.660 ;
        RECT 290.980 56.655 291.270 57.380 ;
        RECT 291.440 56.610 293.110 57.380 ;
        RECT 293.370 56.830 293.540 57.210 ;
        RECT 293.720 57.000 294.050 57.380 ;
        RECT 293.370 56.660 294.035 56.830 ;
        RECT 294.230 56.705 294.490 57.210 ;
        RECT 290.455 55.840 290.805 56.490 ;
        RECT 291.440 56.090 292.190 56.610 ;
        RECT 290.055 55.500 290.805 55.670 ;
        RECT 290.050 54.830 290.380 55.330 ;
        RECT 290.550 55.000 290.805 55.500 ;
        RECT 290.980 54.830 291.270 55.995 ;
        RECT 292.360 55.920 293.110 56.440 ;
        RECT 293.300 56.110 293.630 56.480 ;
        RECT 293.865 56.405 294.035 56.660 ;
        RECT 293.865 56.075 294.150 56.405 ;
        RECT 293.865 55.930 294.035 56.075 ;
        RECT 291.440 54.830 293.110 55.920 ;
        RECT 293.370 55.760 294.035 55.930 ;
        RECT 294.320 55.905 294.490 56.705 ;
        RECT 294.660 56.610 297.250 57.380 ;
        RECT 297.425 56.830 297.680 57.120 ;
        RECT 297.850 57.000 298.180 57.380 ;
        RECT 297.425 56.660 298.175 56.830 ;
        RECT 294.660 56.090 295.870 56.610 ;
        RECT 296.040 55.920 297.250 56.440 ;
        RECT 293.370 55.000 293.540 55.760 ;
        RECT 293.720 54.830 294.050 55.590 ;
        RECT 294.220 55.000 294.490 55.905 ;
        RECT 294.660 54.830 297.250 55.920 ;
        RECT 297.425 55.840 297.775 56.490 ;
        RECT 297.945 55.670 298.175 56.660 ;
        RECT 297.425 55.500 298.175 55.670 ;
        RECT 297.425 55.000 297.680 55.500 ;
        RECT 297.850 54.830 298.180 55.330 ;
        RECT 298.350 55.000 298.520 57.120 ;
        RECT 298.880 57.020 299.210 57.380 ;
        RECT 299.380 56.990 299.875 57.160 ;
        RECT 300.080 56.990 300.935 57.160 ;
        RECT 298.750 55.800 299.210 56.850 ;
        RECT 298.690 55.015 299.015 55.800 ;
        RECT 299.380 55.630 299.550 56.990 ;
        RECT 299.720 56.080 300.070 56.700 ;
        RECT 300.240 56.480 300.595 56.700 ;
        RECT 300.240 55.890 300.410 56.480 ;
        RECT 300.765 56.280 300.935 56.990 ;
        RECT 301.810 56.920 302.140 57.380 ;
        RECT 302.350 57.020 302.700 57.190 ;
        RECT 301.140 56.450 301.930 56.700 ;
        RECT 302.350 56.630 302.610 57.020 ;
        RECT 302.920 56.930 303.870 57.210 ;
        RECT 304.040 56.940 304.230 57.380 ;
        RECT 304.400 57.000 305.470 57.170 ;
        RECT 302.100 56.280 302.270 56.460 ;
        RECT 299.380 55.460 299.775 55.630 ;
        RECT 299.945 55.500 300.410 55.890 ;
        RECT 300.580 56.110 302.270 56.280 ;
        RECT 299.605 55.330 299.775 55.460 ;
        RECT 300.580 55.330 300.750 56.110 ;
        RECT 302.440 55.940 302.610 56.630 ;
        RECT 301.110 55.770 302.610 55.940 ;
        RECT 302.800 55.970 303.010 56.760 ;
        RECT 303.180 56.140 303.530 56.760 ;
        RECT 303.700 56.150 303.870 56.930 ;
        RECT 304.400 56.770 304.570 57.000 ;
        RECT 304.040 56.600 304.570 56.770 ;
        RECT 304.040 56.320 304.260 56.600 ;
        RECT 304.740 56.430 304.980 56.830 ;
        RECT 303.700 55.980 304.105 56.150 ;
        RECT 304.440 56.060 304.980 56.430 ;
        RECT 305.150 56.645 305.470 57.000 ;
        RECT 305.715 56.920 306.020 57.380 ;
        RECT 306.190 56.670 306.440 57.200 ;
        RECT 305.150 56.470 305.475 56.645 ;
        RECT 305.150 56.170 306.065 56.470 ;
        RECT 305.325 56.140 306.065 56.170 ;
        RECT 302.800 55.810 303.475 55.970 ;
        RECT 303.935 55.890 304.105 55.980 ;
        RECT 302.800 55.800 303.765 55.810 ;
        RECT 302.440 55.630 302.610 55.770 ;
        RECT 299.185 54.830 299.435 55.290 ;
        RECT 299.605 55.000 299.855 55.330 ;
        RECT 300.070 55.000 300.750 55.330 ;
        RECT 300.920 55.430 301.995 55.600 ;
        RECT 302.440 55.460 303.000 55.630 ;
        RECT 303.305 55.510 303.765 55.800 ;
        RECT 303.935 55.720 305.155 55.890 ;
        RECT 300.920 55.090 301.090 55.430 ;
        RECT 301.325 54.830 301.655 55.260 ;
        RECT 301.825 55.090 301.995 55.430 ;
        RECT 302.290 54.830 302.660 55.290 ;
        RECT 302.830 55.000 303.000 55.460 ;
        RECT 303.935 55.340 304.105 55.720 ;
        RECT 305.325 55.550 305.495 56.140 ;
        RECT 306.235 56.020 306.440 56.670 ;
        RECT 306.610 56.625 306.860 57.380 ;
        RECT 307.080 56.630 308.290 57.380 ;
        RECT 308.460 56.705 308.720 57.210 ;
        RECT 308.900 57.000 309.230 57.380 ;
        RECT 309.410 56.830 309.580 57.210 ;
        RECT 307.080 56.090 307.600 56.630 ;
        RECT 303.235 55.000 304.105 55.340 ;
        RECT 304.695 55.380 305.495 55.550 ;
        RECT 304.275 54.830 304.525 55.290 ;
        RECT 304.695 55.090 304.865 55.380 ;
        RECT 305.045 54.830 305.375 55.210 ;
        RECT 305.715 54.830 306.020 55.970 ;
        RECT 306.190 55.140 306.440 56.020 ;
        RECT 306.610 54.830 306.860 55.970 ;
        RECT 307.770 55.920 308.290 56.460 ;
        RECT 307.080 54.830 308.290 55.920 ;
        RECT 308.460 55.905 308.630 56.705 ;
        RECT 308.915 56.660 309.580 56.830 ;
        RECT 308.915 56.405 309.085 56.660 ;
        RECT 309.840 56.630 311.050 57.380 ;
        RECT 308.800 56.075 309.085 56.405 ;
        RECT 309.320 56.110 309.650 56.480 ;
        RECT 308.915 55.930 309.085 56.075 ;
        RECT 308.460 55.000 308.730 55.905 ;
        RECT 308.915 55.760 309.580 55.930 ;
        RECT 308.900 54.830 309.230 55.590 ;
        RECT 309.410 55.000 309.580 55.760 ;
        RECT 309.840 55.920 310.360 56.460 ;
        RECT 310.530 56.090 311.050 56.630 ;
        RECT 309.840 54.830 311.050 55.920 ;
        RECT 162.095 54.660 311.135 54.830 ;
        RECT 162.180 53.570 163.390 54.660 ;
        RECT 163.560 53.570 165.230 54.660 ;
        RECT 165.405 53.990 165.660 54.490 ;
        RECT 165.830 54.160 166.160 54.660 ;
        RECT 165.405 53.820 166.155 53.990 ;
        RECT 162.180 52.860 162.700 53.400 ;
        RECT 162.870 53.030 163.390 53.570 ;
        RECT 163.560 52.880 164.310 53.400 ;
        RECT 164.480 53.050 165.230 53.570 ;
        RECT 165.405 53.000 165.755 53.650 ;
        RECT 162.180 52.110 163.390 52.860 ;
        RECT 163.560 52.110 165.230 52.880 ;
        RECT 165.925 52.830 166.155 53.820 ;
        RECT 165.405 52.660 166.155 52.830 ;
        RECT 165.405 52.370 165.660 52.660 ;
        RECT 165.830 52.110 166.160 52.490 ;
        RECT 166.330 52.370 166.500 54.490 ;
        RECT 166.670 53.690 166.995 54.475 ;
        RECT 167.165 54.200 167.415 54.660 ;
        RECT 167.585 54.160 167.835 54.490 ;
        RECT 168.050 54.160 168.730 54.490 ;
        RECT 167.585 54.030 167.755 54.160 ;
        RECT 167.360 53.860 167.755 54.030 ;
        RECT 166.730 52.640 167.190 53.690 ;
        RECT 167.360 52.500 167.530 53.860 ;
        RECT 167.925 53.600 168.390 53.990 ;
        RECT 167.700 52.790 168.050 53.410 ;
        RECT 168.220 53.010 168.390 53.600 ;
        RECT 168.560 53.380 168.730 54.160 ;
        RECT 168.900 54.060 169.070 54.400 ;
        RECT 169.305 54.230 169.635 54.660 ;
        RECT 169.805 54.060 169.975 54.400 ;
        RECT 170.270 54.200 170.640 54.660 ;
        RECT 168.900 53.890 169.975 54.060 ;
        RECT 170.810 54.030 170.980 54.490 ;
        RECT 171.215 54.150 172.085 54.490 ;
        RECT 172.255 54.200 172.505 54.660 ;
        RECT 170.420 53.860 170.980 54.030 ;
        RECT 170.420 53.720 170.590 53.860 ;
        RECT 169.090 53.550 170.590 53.720 ;
        RECT 171.285 53.690 171.745 53.980 ;
        RECT 168.560 53.210 170.250 53.380 ;
        RECT 168.220 52.790 168.575 53.010 ;
        RECT 168.745 52.500 168.915 53.210 ;
        RECT 169.120 52.790 169.910 53.040 ;
        RECT 170.080 53.030 170.250 53.210 ;
        RECT 170.420 52.860 170.590 53.550 ;
        RECT 166.860 52.110 167.190 52.470 ;
        RECT 167.360 52.330 167.855 52.500 ;
        RECT 168.060 52.330 168.915 52.500 ;
        RECT 169.790 52.110 170.120 52.570 ;
        RECT 170.330 52.470 170.590 52.860 ;
        RECT 170.780 53.680 171.745 53.690 ;
        RECT 171.915 53.770 172.085 54.150 ;
        RECT 172.675 54.110 172.845 54.400 ;
        RECT 173.025 54.280 173.355 54.660 ;
        RECT 172.675 53.940 173.475 54.110 ;
        RECT 170.780 53.520 171.455 53.680 ;
        RECT 171.915 53.600 173.135 53.770 ;
        RECT 170.780 52.730 170.990 53.520 ;
        RECT 171.915 53.510 172.085 53.600 ;
        RECT 171.160 52.730 171.510 53.350 ;
        RECT 171.680 53.340 172.085 53.510 ;
        RECT 171.680 52.560 171.850 53.340 ;
        RECT 172.020 52.890 172.240 53.170 ;
        RECT 172.420 53.060 172.960 53.430 ;
        RECT 173.305 53.350 173.475 53.940 ;
        RECT 173.695 53.520 174.000 54.660 ;
        RECT 174.170 53.470 174.420 54.350 ;
        RECT 174.590 53.520 174.840 54.660 ;
        RECT 175.060 53.495 175.350 54.660 ;
        RECT 175.520 53.585 175.790 54.490 ;
        RECT 175.960 53.900 176.290 54.660 ;
        RECT 176.470 53.730 176.640 54.490 ;
        RECT 173.305 53.320 174.045 53.350 ;
        RECT 172.020 52.720 172.550 52.890 ;
        RECT 170.330 52.300 170.680 52.470 ;
        RECT 170.900 52.280 171.850 52.560 ;
        RECT 172.020 52.110 172.210 52.550 ;
        RECT 172.380 52.490 172.550 52.720 ;
        RECT 172.720 52.660 172.960 53.060 ;
        RECT 173.130 53.020 174.045 53.320 ;
        RECT 173.130 52.845 173.455 53.020 ;
        RECT 173.130 52.490 173.450 52.845 ;
        RECT 174.215 52.820 174.420 53.470 ;
        RECT 172.380 52.320 173.450 52.490 ;
        RECT 173.695 52.110 174.000 52.570 ;
        RECT 174.170 52.290 174.420 52.820 ;
        RECT 174.590 52.110 174.840 52.865 ;
        RECT 175.060 52.110 175.350 52.835 ;
        RECT 175.520 52.785 175.690 53.585 ;
        RECT 175.975 53.560 176.640 53.730 ;
        RECT 176.900 53.570 180.410 54.660 ;
        RECT 175.975 53.415 176.145 53.560 ;
        RECT 175.860 53.085 176.145 53.415 ;
        RECT 175.975 52.830 176.145 53.085 ;
        RECT 176.380 53.010 176.710 53.380 ;
        RECT 176.900 52.880 178.550 53.400 ;
        RECT 178.720 53.050 180.410 53.570 ;
        RECT 180.580 53.585 180.850 54.490 ;
        RECT 181.020 53.900 181.350 54.660 ;
        RECT 181.530 53.730 181.700 54.490 ;
        RECT 181.960 54.225 187.305 54.660 ;
        RECT 175.520 52.280 175.780 52.785 ;
        RECT 175.975 52.660 176.640 52.830 ;
        RECT 175.960 52.110 176.290 52.490 ;
        RECT 176.470 52.280 176.640 52.660 ;
        RECT 176.900 52.110 180.410 52.880 ;
        RECT 180.580 52.785 180.750 53.585 ;
        RECT 181.035 53.560 181.700 53.730 ;
        RECT 181.035 53.415 181.205 53.560 ;
        RECT 180.920 53.085 181.205 53.415 ;
        RECT 181.035 52.830 181.205 53.085 ;
        RECT 181.440 53.010 181.770 53.380 ;
        RECT 180.580 52.280 180.840 52.785 ;
        RECT 181.035 52.660 181.700 52.830 ;
        RECT 181.020 52.110 181.350 52.490 ;
        RECT 181.530 52.280 181.700 52.660 ;
        RECT 183.545 52.655 183.885 53.485 ;
        RECT 185.365 52.975 185.715 54.225 ;
        RECT 187.480 53.570 190.070 54.660 ;
        RECT 190.490 53.930 190.785 54.660 ;
        RECT 190.955 53.760 191.215 54.485 ;
        RECT 191.385 53.930 191.645 54.660 ;
        RECT 191.815 53.760 192.075 54.485 ;
        RECT 192.245 53.930 192.505 54.660 ;
        RECT 192.675 53.760 192.935 54.485 ;
        RECT 193.105 53.930 193.365 54.660 ;
        RECT 193.535 53.760 193.795 54.485 ;
        RECT 187.480 52.880 188.690 53.400 ;
        RECT 188.860 53.050 190.070 53.570 ;
        RECT 190.485 53.520 193.795 53.760 ;
        RECT 193.965 53.550 194.225 54.660 ;
        RECT 190.485 52.930 191.455 53.520 ;
        RECT 194.395 53.350 194.645 54.485 ;
        RECT 194.825 53.550 195.120 54.660 ;
        RECT 195.300 54.225 200.645 54.660 ;
        RECT 191.625 53.100 194.645 53.350 ;
        RECT 181.960 52.110 187.305 52.655 ;
        RECT 187.480 52.110 190.070 52.880 ;
        RECT 190.485 52.760 193.795 52.930 ;
        RECT 190.485 52.110 190.785 52.590 ;
        RECT 190.955 52.305 191.215 52.760 ;
        RECT 191.385 52.110 191.645 52.590 ;
        RECT 191.815 52.305 192.075 52.760 ;
        RECT 192.245 52.110 192.505 52.590 ;
        RECT 192.675 52.305 192.935 52.760 ;
        RECT 193.105 52.110 193.365 52.590 ;
        RECT 193.535 52.305 193.795 52.760 ;
        RECT 193.965 52.110 194.225 52.635 ;
        RECT 194.395 52.290 194.645 53.100 ;
        RECT 194.815 52.740 195.130 53.350 ;
        RECT 196.885 52.655 197.225 53.485 ;
        RECT 198.705 52.975 199.055 54.225 ;
        RECT 200.820 53.495 201.110 54.660 ;
        RECT 201.280 54.060 201.540 54.480 ;
        RECT 201.710 54.230 202.040 54.660 ;
        RECT 202.320 54.320 203.640 54.490 ;
        RECT 202.320 54.060 202.490 54.320 ;
        RECT 201.280 53.890 202.490 54.060 ;
        RECT 202.705 53.980 203.300 54.150 ;
        RECT 201.280 52.850 201.450 53.890 ;
        RECT 201.620 53.020 201.970 53.720 ;
        RECT 202.185 53.550 202.790 53.720 ;
        RECT 202.600 53.350 202.790 53.550 ;
        RECT 202.140 53.020 202.430 53.350 ;
        RECT 202.600 53.020 202.890 53.350 ;
        RECT 202.600 52.850 202.790 53.020 ;
        RECT 194.825 52.110 195.070 52.570 ;
        RECT 195.300 52.110 200.645 52.655 ;
        RECT 200.820 52.110 201.110 52.835 ;
        RECT 201.280 52.475 201.595 52.850 ;
        RECT 201.850 52.110 202.020 52.850 ;
        RECT 202.270 52.680 202.790 52.850 ;
        RECT 203.130 52.850 203.300 53.980 ;
        RECT 203.470 53.020 203.640 54.320 ;
        RECT 203.990 53.810 204.310 54.400 ;
        RECT 204.595 53.820 204.845 54.660 ;
        RECT 203.990 53.475 204.200 53.810 ;
        RECT 205.070 53.650 205.320 54.490 ;
        RECT 205.490 53.820 205.740 54.660 ;
        RECT 205.910 53.650 206.160 54.490 ;
        RECT 206.330 53.820 206.580 54.660 ;
        RECT 203.870 53.020 204.200 53.475 ;
        RECT 204.430 53.470 204.865 53.640 ;
        RECT 205.070 53.480 206.630 53.650 ;
        RECT 206.800 53.570 209.390 54.660 ;
        RECT 209.650 54.080 209.820 54.490 ;
        RECT 209.990 54.280 210.320 54.660 ;
        RECT 210.965 54.280 211.635 54.660 ;
        RECT 211.870 54.110 212.040 54.490 ;
        RECT 212.210 54.280 212.550 54.660 ;
        RECT 212.720 54.110 212.890 54.490 ;
        RECT 213.230 54.280 213.560 54.660 ;
        RECT 213.730 54.110 213.990 54.490 ;
        RECT 214.170 54.280 214.500 54.660 ;
        RECT 209.650 53.910 211.400 54.080 ;
        RECT 205.480 53.470 205.650 53.480 ;
        RECT 204.430 53.020 204.600 53.470 ;
        RECT 204.770 53.100 206.230 53.270 ;
        RECT 204.770 52.850 204.940 53.100 ;
        RECT 206.400 52.930 206.630 53.480 ;
        RECT 203.130 52.680 204.940 52.850 ;
        RECT 205.110 52.750 206.630 52.930 ;
        RECT 206.800 52.880 208.010 53.400 ;
        RECT 208.180 53.050 209.390 53.570 ;
        RECT 209.625 53.300 209.805 53.660 ;
        RECT 209.620 53.130 209.805 53.300 ;
        RECT 209.625 53.020 209.805 53.130 ;
        RECT 202.270 52.475 202.440 52.680 ;
        RECT 202.710 52.110 203.040 52.505 ;
        RECT 203.290 52.330 203.460 52.680 ;
        RECT 203.660 52.110 203.990 52.510 ;
        RECT 204.160 52.330 204.330 52.680 ;
        RECT 204.550 52.110 204.930 52.510 ;
        RECT 205.110 52.280 205.360 52.750 ;
        RECT 205.530 52.110 205.700 52.580 ;
        RECT 205.870 52.280 206.200 52.750 ;
        RECT 206.370 52.110 206.540 52.580 ;
        RECT 206.800 52.110 209.390 52.880 ;
        RECT 209.975 52.830 210.145 53.910 ;
        RECT 210.465 53.570 210.795 53.740 ;
        RECT 209.650 52.660 210.145 52.830 ;
        RECT 209.650 52.280 209.820 52.660 ;
        RECT 209.990 52.110 210.320 52.490 ;
        RECT 210.490 52.280 210.715 53.570 ;
        RECT 211.230 53.350 211.400 53.910 ;
        RECT 211.710 53.940 212.890 54.110 ;
        RECT 213.060 53.940 213.990 54.110 ;
        RECT 210.890 52.830 211.060 53.350 ;
        RECT 211.230 53.020 211.540 53.350 ;
        RECT 211.710 52.830 211.880 53.940 ;
        RECT 213.060 53.770 213.230 53.940 ;
        RECT 212.050 53.600 213.230 53.770 ;
        RECT 212.050 53.425 212.220 53.600 ;
        RECT 212.380 53.130 212.650 53.300 ;
        RECT 210.890 52.660 211.880 52.830 ;
        RECT 210.885 52.110 211.215 52.490 ;
        RECT 211.485 52.280 211.655 52.660 ;
        RECT 212.385 52.445 212.650 53.130 ;
        RECT 212.825 52.450 213.130 53.430 ;
        RECT 213.300 52.790 213.650 53.330 ;
        RECT 213.820 52.610 213.990 53.940 ;
        RECT 214.200 52.780 214.405 54.100 ;
        RECT 214.675 53.690 214.925 54.490 ;
        RECT 215.145 53.940 215.475 54.660 ;
        RECT 215.660 53.690 215.910 54.490 ;
        RECT 216.310 53.860 216.640 54.660 ;
        RECT 216.810 54.320 217.145 54.490 ;
        RECT 216.810 54.150 217.150 54.320 ;
        RECT 214.575 53.520 216.630 53.690 ;
        RECT 216.810 53.520 217.145 54.150 ;
        RECT 217.320 53.860 217.650 54.660 ;
        RECT 218.140 54.020 218.470 54.450 ;
        RECT 214.575 52.610 214.745 53.520 ;
        RECT 213.310 52.110 213.560 52.610 ;
        RECT 213.730 52.280 213.990 52.610 ;
        RECT 214.250 52.280 214.745 52.610 ;
        RECT 214.965 52.445 215.320 53.350 ;
        RECT 215.495 53.330 215.665 53.350 ;
        RECT 215.495 52.440 215.795 53.330 ;
        RECT 215.975 52.440 216.235 53.350 ;
        RECT 216.405 53.340 216.630 53.520 ;
        RECT 216.405 53.100 216.800 53.340 ;
        RECT 216.405 52.110 216.640 52.915 ;
        RECT 216.970 52.830 217.145 53.520 ;
        RECT 218.015 53.850 218.470 54.020 ;
        RECT 218.650 54.020 218.900 54.440 ;
        RECT 219.130 54.190 219.460 54.660 ;
        RECT 219.690 54.020 219.940 54.440 ;
        RECT 218.650 53.850 219.940 54.020 ;
        RECT 218.015 52.850 218.185 53.850 ;
        RECT 218.355 53.020 218.600 53.680 ;
        RECT 218.815 53.020 219.080 53.680 ;
        RECT 219.275 53.020 219.560 53.680 ;
        RECT 219.735 53.350 219.950 53.680 ;
        RECT 220.130 53.520 220.380 54.660 ;
        RECT 220.550 53.600 220.880 54.450 ;
        RECT 221.330 53.860 221.580 54.660 ;
        RECT 219.735 53.020 220.040 53.350 ;
        RECT 220.210 53.020 220.520 53.350 ;
        RECT 220.210 52.850 220.380 53.020 ;
        RECT 216.810 52.365 217.145 52.830 ;
        RECT 216.810 52.320 217.140 52.365 ;
        RECT 217.330 52.110 217.660 52.835 ;
        RECT 218.015 52.680 220.380 52.850 ;
        RECT 220.690 52.835 220.880 53.600 ;
        RECT 221.750 53.690 222.080 54.490 ;
        RECT 222.250 53.860 222.420 54.660 ;
        RECT 222.590 53.690 222.920 54.490 ;
        RECT 223.090 53.860 223.260 54.660 ;
        RECT 223.430 53.690 223.760 54.490 ;
        RECT 223.930 53.860 224.100 54.660 ;
        RECT 224.270 53.690 224.600 54.490 ;
        RECT 221.750 53.520 224.600 53.690 ;
        RECT 224.770 53.520 225.025 54.660 ;
        RECT 225.200 53.570 226.410 54.660 ;
        RECT 221.060 53.100 222.500 53.350 ;
        RECT 222.670 53.100 223.205 53.520 ;
        RECT 223.385 53.100 225.005 53.350 ;
        RECT 218.170 52.110 218.500 52.510 ;
        RECT 218.670 52.340 219.000 52.680 ;
        RECT 220.050 52.110 220.380 52.510 ;
        RECT 220.550 52.325 220.880 52.835 ;
        RECT 221.330 52.490 221.580 52.910 ;
        RECT 222.670 52.830 222.920 53.100 ;
        RECT 221.750 52.660 222.920 52.830 ;
        RECT 223.090 52.740 225.025 52.930 ;
        RECT 223.090 52.490 223.340 52.740 ;
        RECT 221.330 52.280 223.340 52.490 ;
        RECT 223.510 52.110 223.680 52.570 ;
        RECT 223.850 52.280 224.180 52.740 ;
        RECT 224.350 52.110 224.520 52.570 ;
        RECT 224.690 52.280 225.025 52.740 ;
        RECT 225.200 52.860 225.720 53.400 ;
        RECT 225.890 53.030 226.410 53.570 ;
        RECT 226.580 53.495 226.870 54.660 ;
        RECT 225.200 52.110 226.410 52.860 ;
        RECT 226.580 52.110 226.870 52.835 ;
        RECT 227.040 52.390 227.320 54.490 ;
        RECT 227.510 53.900 228.295 54.660 ;
        RECT 228.690 53.830 229.075 54.490 ;
        RECT 228.690 53.730 229.100 53.830 ;
        RECT 227.490 53.520 229.100 53.730 ;
        RECT 229.400 53.640 229.600 54.430 ;
        RECT 227.490 52.920 227.765 53.520 ;
        RECT 229.270 53.470 229.600 53.640 ;
        RECT 229.770 53.480 230.090 54.660 ;
        RECT 230.720 53.520 231.105 54.490 ;
        RECT 231.275 54.200 231.600 54.660 ;
        RECT 232.120 54.030 232.400 54.490 ;
        RECT 231.275 53.810 232.400 54.030 ;
        RECT 229.270 53.350 229.450 53.470 ;
        RECT 227.935 53.100 228.290 53.350 ;
        RECT 228.485 53.300 228.950 53.350 ;
        RECT 228.480 53.130 228.950 53.300 ;
        RECT 228.485 53.100 228.950 53.130 ;
        RECT 229.120 53.100 229.450 53.350 ;
        RECT 229.625 53.100 230.090 53.300 ;
        RECT 227.490 52.740 228.740 52.920 ;
        RECT 228.375 52.670 228.740 52.740 ;
        RECT 228.910 52.720 230.090 52.890 ;
        RECT 227.550 52.110 227.720 52.570 ;
        RECT 228.910 52.500 229.240 52.720 ;
        RECT 227.990 52.320 229.240 52.500 ;
        RECT 229.410 52.110 229.580 52.550 ;
        RECT 229.750 52.305 230.090 52.720 ;
        RECT 230.720 52.850 231.000 53.520 ;
        RECT 231.275 53.350 231.725 53.810 ;
        RECT 232.590 53.640 232.990 54.490 ;
        RECT 233.390 54.200 233.660 54.660 ;
        RECT 233.830 54.030 234.115 54.490 ;
        RECT 231.170 53.020 231.725 53.350 ;
        RECT 231.895 53.080 232.990 53.640 ;
        RECT 231.275 52.910 231.725 53.020 ;
        RECT 230.720 52.280 231.105 52.850 ;
        RECT 231.275 52.740 232.400 52.910 ;
        RECT 231.275 52.110 231.600 52.570 ;
        RECT 232.120 52.280 232.400 52.740 ;
        RECT 232.590 52.280 232.990 53.080 ;
        RECT 233.160 53.810 234.115 54.030 ;
        RECT 233.160 52.910 233.370 53.810 ;
        RECT 233.540 53.080 234.230 53.640 ;
        RECT 234.400 53.520 234.785 54.480 ;
        RECT 235.000 53.860 235.290 54.660 ;
        RECT 235.460 54.320 236.825 54.490 ;
        RECT 235.460 53.690 235.630 54.320 ;
        RECT 234.955 53.520 235.630 53.690 ;
        RECT 233.160 52.740 234.115 52.910 ;
        RECT 233.390 52.110 233.660 52.570 ;
        RECT 233.830 52.280 234.115 52.740 ;
        RECT 234.400 52.850 234.575 53.520 ;
        RECT 234.955 53.350 235.125 53.520 ;
        RECT 235.800 53.350 236.125 54.150 ;
        RECT 236.495 54.110 236.825 54.320 ;
        RECT 236.495 53.860 237.450 54.110 ;
        RECT 234.760 53.100 235.125 53.350 ;
        RECT 235.320 53.100 235.570 53.350 ;
        RECT 234.760 53.020 234.950 53.100 ;
        RECT 235.320 53.020 235.490 53.100 ;
        RECT 235.780 53.020 236.125 53.350 ;
        RECT 236.295 53.020 236.570 53.685 ;
        RECT 236.755 53.020 237.110 53.685 ;
        RECT 237.280 52.850 237.450 53.860 ;
        RECT 237.620 53.520 237.910 54.660 ;
        RECT 237.635 53.020 237.910 53.350 ;
        RECT 234.400 52.280 234.910 52.850 ;
        RECT 235.455 52.680 236.855 52.850 ;
        RECT 235.080 52.110 235.250 52.670 ;
        RECT 235.455 52.280 235.785 52.680 ;
        RECT 235.960 52.110 236.290 52.510 ;
        RECT 236.525 52.490 236.855 52.680 ;
        RECT 237.025 52.660 237.450 52.850 ;
        RECT 237.620 52.490 237.910 52.760 ;
        RECT 236.525 52.280 237.910 52.490 ;
        RECT 238.090 52.280 238.350 54.490 ;
        RECT 238.520 53.860 239.330 54.660 ;
        RECT 239.500 53.690 239.830 54.490 ;
        RECT 240.015 53.860 240.755 54.660 ;
        RECT 240.925 53.690 241.175 54.490 ;
        RECT 238.690 53.520 241.175 53.690 ;
        RECT 238.690 53.350 238.860 53.520 ;
        RECT 241.345 53.350 241.530 54.440 ;
        RECT 241.725 53.860 242.050 54.660 ;
        RECT 238.520 53.020 238.860 53.350 ;
        RECT 239.260 53.100 239.740 53.350 ;
        RECT 238.690 52.930 238.860 53.020 ;
        RECT 238.690 52.760 239.360 52.930 ;
        RECT 238.530 52.110 238.840 52.590 ;
        RECT 239.020 52.280 239.360 52.760 ;
        RECT 239.530 52.415 239.740 53.100 ;
        RECT 239.920 52.415 240.190 53.350 ;
        RECT 240.440 53.020 240.700 53.350 ;
        RECT 241.045 53.100 241.530 53.350 ;
        RECT 241.700 53.100 242.030 53.685 ;
        RECT 242.220 53.570 244.810 54.660 ;
        RECT 240.440 52.415 240.685 53.020 ;
        RECT 240.865 52.730 242.050 52.900 ;
        RECT 240.865 52.280 241.155 52.730 ;
        RECT 241.325 52.110 241.615 52.560 ;
        RECT 241.785 52.280 242.050 52.730 ;
        RECT 242.220 52.880 243.430 53.400 ;
        RECT 243.600 53.050 244.810 53.570 ;
        RECT 244.980 53.520 245.365 54.480 ;
        RECT 245.580 53.860 245.870 54.660 ;
        RECT 246.040 54.320 247.405 54.490 ;
        RECT 246.040 53.690 246.210 54.320 ;
        RECT 245.535 53.520 246.210 53.690 ;
        RECT 244.980 53.470 245.210 53.520 ;
        RECT 242.220 52.110 244.810 52.880 ;
        RECT 244.980 52.850 245.155 53.470 ;
        RECT 245.535 53.350 245.705 53.520 ;
        RECT 246.380 53.350 246.705 54.150 ;
        RECT 247.075 54.110 247.405 54.320 ;
        RECT 247.075 53.860 248.030 54.110 ;
        RECT 245.340 53.100 245.705 53.350 ;
        RECT 245.900 53.100 246.150 53.350 ;
        RECT 245.340 53.020 245.530 53.100 ;
        RECT 245.900 53.020 246.070 53.100 ;
        RECT 246.360 53.020 246.705 53.350 ;
        RECT 246.875 53.020 247.150 53.685 ;
        RECT 247.335 53.020 247.690 53.685 ;
        RECT 247.860 52.850 248.030 53.860 ;
        RECT 248.200 53.520 248.490 54.660 ;
        RECT 248.660 53.790 248.935 54.490 ;
        RECT 249.145 54.115 249.360 54.660 ;
        RECT 249.530 54.150 250.005 54.490 ;
        RECT 250.175 54.155 250.790 54.660 ;
        RECT 250.175 53.980 250.370 54.155 ;
        RECT 248.215 53.020 248.490 53.350 ;
        RECT 244.980 52.280 245.490 52.850 ;
        RECT 246.035 52.680 247.435 52.850 ;
        RECT 245.660 52.110 245.830 52.670 ;
        RECT 246.035 52.280 246.365 52.680 ;
        RECT 246.540 52.110 246.870 52.510 ;
        RECT 247.105 52.490 247.435 52.680 ;
        RECT 247.605 52.660 248.030 52.850 ;
        RECT 248.660 52.760 248.830 53.790 ;
        RECT 249.105 53.620 249.820 53.915 ;
        RECT 250.040 53.790 250.370 53.980 ;
        RECT 250.540 53.620 250.790 53.985 ;
        RECT 249.000 53.450 250.790 53.620 ;
        RECT 249.000 53.020 249.230 53.450 ;
        RECT 248.200 52.490 248.490 52.760 ;
        RECT 247.105 52.280 248.490 52.490 ;
        RECT 248.660 52.280 248.920 52.760 ;
        RECT 249.400 52.750 249.810 53.270 ;
        RECT 249.090 52.110 249.420 52.570 ;
        RECT 249.610 52.330 249.810 52.750 ;
        RECT 249.980 52.595 250.235 53.450 ;
        RECT 251.030 53.270 251.200 54.490 ;
        RECT 251.450 54.150 251.710 54.660 ;
        RECT 250.405 53.020 251.200 53.270 ;
        RECT 251.370 53.100 251.710 53.980 ;
        RECT 252.340 53.495 252.630 54.660 ;
        RECT 252.800 53.520 253.080 54.660 ;
        RECT 253.250 53.510 253.580 54.490 ;
        RECT 253.750 53.520 254.010 54.660 ;
        RECT 254.180 54.225 259.525 54.660 ;
        RECT 252.810 53.080 253.145 53.350 ;
        RECT 250.950 52.930 251.200 53.020 ;
        RECT 249.980 52.330 250.770 52.595 ;
        RECT 250.950 52.510 251.280 52.930 ;
        RECT 251.450 52.110 251.710 52.930 ;
        RECT 253.315 52.910 253.485 53.510 ;
        RECT 253.655 53.100 253.990 53.350 ;
        RECT 252.340 52.110 252.630 52.835 ;
        RECT 252.800 52.110 253.110 52.910 ;
        RECT 253.315 52.280 254.010 52.910 ;
        RECT 255.765 52.655 256.105 53.485 ;
        RECT 257.585 52.975 257.935 54.225 ;
        RECT 259.885 53.690 260.275 53.865 ;
        RECT 260.760 53.860 261.090 54.660 ;
        RECT 261.260 53.870 261.795 54.490 ;
        RECT 259.885 53.520 261.310 53.690 ;
        RECT 259.760 52.790 260.115 53.350 ;
        RECT 254.180 52.110 259.525 52.655 ;
        RECT 260.285 52.620 260.455 53.520 ;
        RECT 260.625 52.790 260.890 53.350 ;
        RECT 261.140 53.020 261.310 53.520 ;
        RECT 261.480 52.850 261.795 53.870 ;
        RECT 262.005 53.990 262.260 54.490 ;
        RECT 262.430 54.160 262.760 54.660 ;
        RECT 262.005 53.820 262.755 53.990 ;
        RECT 262.005 53.000 262.355 53.650 ;
        RECT 259.865 52.110 260.105 52.620 ;
        RECT 260.285 52.290 260.565 52.620 ;
        RECT 260.795 52.110 261.010 52.620 ;
        RECT 261.180 52.280 261.795 52.850 ;
        RECT 262.525 52.830 262.755 53.820 ;
        RECT 262.005 52.660 262.755 52.830 ;
        RECT 262.005 52.370 262.260 52.660 ;
        RECT 262.430 52.110 262.760 52.490 ;
        RECT 262.930 52.370 263.100 54.490 ;
        RECT 263.270 53.690 263.595 54.475 ;
        RECT 263.765 54.200 264.015 54.660 ;
        RECT 264.185 54.160 264.435 54.490 ;
        RECT 264.650 54.160 265.330 54.490 ;
        RECT 264.185 54.030 264.355 54.160 ;
        RECT 263.960 53.860 264.355 54.030 ;
        RECT 263.330 52.640 263.790 53.690 ;
        RECT 263.960 52.500 264.130 53.860 ;
        RECT 264.525 53.600 264.990 53.990 ;
        RECT 264.300 52.790 264.650 53.410 ;
        RECT 264.820 53.010 264.990 53.600 ;
        RECT 265.160 53.380 265.330 54.160 ;
        RECT 265.500 54.060 265.670 54.400 ;
        RECT 265.905 54.230 266.235 54.660 ;
        RECT 266.405 54.060 266.575 54.400 ;
        RECT 266.870 54.200 267.240 54.660 ;
        RECT 265.500 53.890 266.575 54.060 ;
        RECT 267.410 54.030 267.580 54.490 ;
        RECT 267.815 54.150 268.685 54.490 ;
        RECT 268.855 54.200 269.105 54.660 ;
        RECT 267.020 53.860 267.580 54.030 ;
        RECT 267.020 53.720 267.190 53.860 ;
        RECT 265.690 53.550 267.190 53.720 ;
        RECT 267.885 53.690 268.345 53.980 ;
        RECT 265.160 53.210 266.850 53.380 ;
        RECT 264.820 52.790 265.175 53.010 ;
        RECT 265.345 52.500 265.515 53.210 ;
        RECT 265.720 52.790 266.510 53.040 ;
        RECT 266.680 53.030 266.850 53.210 ;
        RECT 267.020 52.860 267.190 53.550 ;
        RECT 263.460 52.110 263.790 52.470 ;
        RECT 263.960 52.330 264.455 52.500 ;
        RECT 264.660 52.330 265.515 52.500 ;
        RECT 266.390 52.110 266.720 52.570 ;
        RECT 266.930 52.470 267.190 52.860 ;
        RECT 267.380 53.680 268.345 53.690 ;
        RECT 268.515 53.770 268.685 54.150 ;
        RECT 269.275 54.110 269.445 54.400 ;
        RECT 269.625 54.280 269.955 54.660 ;
        RECT 269.275 53.940 270.075 54.110 ;
        RECT 267.380 53.520 268.055 53.680 ;
        RECT 268.515 53.600 269.735 53.770 ;
        RECT 267.380 52.730 267.590 53.520 ;
        RECT 268.515 53.510 268.685 53.600 ;
        RECT 267.760 52.730 268.110 53.350 ;
        RECT 268.280 53.340 268.685 53.510 ;
        RECT 268.280 52.560 268.450 53.340 ;
        RECT 268.620 52.890 268.840 53.170 ;
        RECT 269.020 53.060 269.560 53.430 ;
        RECT 269.905 53.350 270.075 53.940 ;
        RECT 270.295 53.520 270.600 54.660 ;
        RECT 270.770 53.470 271.025 54.350 ;
        RECT 269.905 53.320 270.645 53.350 ;
        RECT 268.620 52.720 269.150 52.890 ;
        RECT 266.930 52.300 267.280 52.470 ;
        RECT 267.500 52.280 268.450 52.560 ;
        RECT 268.620 52.110 268.810 52.550 ;
        RECT 268.980 52.490 269.150 52.720 ;
        RECT 269.320 52.660 269.560 53.060 ;
        RECT 269.730 53.020 270.645 53.320 ;
        RECT 269.730 52.845 270.055 53.020 ;
        RECT 269.730 52.490 270.050 52.845 ;
        RECT 270.815 52.820 271.025 53.470 ;
        RECT 268.980 52.320 270.050 52.490 ;
        RECT 270.295 52.110 270.600 52.570 ;
        RECT 270.770 52.290 271.025 52.820 ;
        RECT 271.200 53.520 271.585 54.490 ;
        RECT 271.755 54.200 272.080 54.660 ;
        RECT 272.600 54.030 272.880 54.490 ;
        RECT 271.755 53.810 272.880 54.030 ;
        RECT 271.200 52.850 271.480 53.520 ;
        RECT 271.755 53.350 272.205 53.810 ;
        RECT 273.070 53.640 273.470 54.490 ;
        RECT 273.870 54.200 274.140 54.660 ;
        RECT 274.310 54.030 274.595 54.490 ;
        RECT 271.650 53.020 272.205 53.350 ;
        RECT 272.375 53.080 273.470 53.640 ;
        RECT 271.755 52.910 272.205 53.020 ;
        RECT 271.200 52.280 271.585 52.850 ;
        RECT 271.755 52.740 272.880 52.910 ;
        RECT 271.755 52.110 272.080 52.570 ;
        RECT 272.600 52.280 272.880 52.740 ;
        RECT 273.070 52.280 273.470 53.080 ;
        RECT 273.640 53.810 274.595 54.030 ;
        RECT 273.640 52.910 273.850 53.810 ;
        RECT 274.020 53.080 274.710 53.640 ;
        RECT 274.880 53.570 277.470 54.660 ;
        RECT 273.640 52.740 274.595 52.910 ;
        RECT 273.870 52.110 274.140 52.570 ;
        RECT 274.310 52.280 274.595 52.740 ;
        RECT 274.880 52.880 276.090 53.400 ;
        RECT 276.260 53.050 277.470 53.570 ;
        RECT 278.100 53.495 278.390 54.660 ;
        RECT 278.560 53.570 280.230 54.660 ;
        RECT 278.560 52.880 279.310 53.400 ;
        RECT 279.480 53.050 280.230 53.570 ;
        RECT 280.400 53.940 280.860 54.490 ;
        RECT 281.050 53.940 281.380 54.660 ;
        RECT 274.880 52.110 277.470 52.880 ;
        RECT 278.100 52.110 278.390 52.835 ;
        RECT 278.560 52.110 280.230 52.880 ;
        RECT 280.400 52.570 280.650 53.940 ;
        RECT 281.580 53.770 281.880 54.320 ;
        RECT 282.050 53.990 282.330 54.660 ;
        RECT 280.940 53.600 281.880 53.770 ;
        RECT 280.940 53.350 281.110 53.600 ;
        RECT 282.250 53.350 282.515 53.710 ;
        RECT 282.700 53.570 284.370 54.660 ;
        RECT 280.820 53.020 281.110 53.350 ;
        RECT 281.280 53.100 281.620 53.350 ;
        RECT 281.840 53.100 282.515 53.350 ;
        RECT 280.940 52.930 281.110 53.020 ;
        RECT 280.940 52.740 282.330 52.930 ;
        RECT 280.400 52.280 280.960 52.570 ;
        RECT 281.130 52.110 281.380 52.570 ;
        RECT 282.000 52.380 282.330 52.740 ;
        RECT 282.700 52.880 283.450 53.400 ;
        RECT 283.620 53.050 284.370 53.570 ;
        RECT 284.550 53.550 284.845 54.660 ;
        RECT 285.025 53.350 285.275 54.485 ;
        RECT 285.445 53.550 285.705 54.660 ;
        RECT 285.875 53.760 286.135 54.485 ;
        RECT 286.305 53.930 286.565 54.660 ;
        RECT 286.735 53.760 286.995 54.485 ;
        RECT 287.165 53.930 287.425 54.660 ;
        RECT 287.595 53.760 287.855 54.485 ;
        RECT 288.025 53.930 288.285 54.660 ;
        RECT 288.455 53.760 288.715 54.485 ;
        RECT 288.885 53.930 289.180 54.660 ;
        RECT 285.875 53.520 289.185 53.760 ;
        RECT 289.600 53.570 291.270 54.660 ;
        RECT 282.700 52.110 284.370 52.880 ;
        RECT 284.540 52.740 284.855 53.350 ;
        RECT 285.025 53.100 288.045 53.350 ;
        RECT 284.600 52.110 284.845 52.570 ;
        RECT 285.025 52.290 285.275 53.100 ;
        RECT 288.215 52.930 289.185 53.520 ;
        RECT 285.875 52.760 289.185 52.930 ;
        RECT 289.600 52.880 290.350 53.400 ;
        RECT 290.520 53.050 291.270 53.570 ;
        RECT 291.440 53.940 291.900 54.490 ;
        RECT 292.090 53.940 292.420 54.660 ;
        RECT 285.445 52.110 285.705 52.635 ;
        RECT 285.875 52.305 286.135 52.760 ;
        RECT 286.305 52.110 286.565 52.590 ;
        RECT 286.735 52.305 286.995 52.760 ;
        RECT 287.165 52.110 287.425 52.590 ;
        RECT 287.595 52.305 287.855 52.760 ;
        RECT 288.025 52.110 288.285 52.590 ;
        RECT 288.455 52.305 288.715 52.760 ;
        RECT 288.885 52.110 289.185 52.590 ;
        RECT 289.600 52.110 291.270 52.880 ;
        RECT 291.440 52.570 291.690 53.940 ;
        RECT 292.620 53.770 292.920 54.320 ;
        RECT 293.090 53.990 293.370 54.660 ;
        RECT 294.665 53.990 294.920 54.490 ;
        RECT 295.090 54.160 295.420 54.660 ;
        RECT 294.665 53.820 295.415 53.990 ;
        RECT 291.980 53.600 292.920 53.770 ;
        RECT 291.980 53.350 292.150 53.600 ;
        RECT 293.290 53.350 293.555 53.710 ;
        RECT 291.860 53.020 292.150 53.350 ;
        RECT 292.320 53.100 292.660 53.350 ;
        RECT 292.880 53.100 293.555 53.350 ;
        RECT 291.980 52.930 292.150 53.020 ;
        RECT 294.665 53.000 295.015 53.650 ;
        RECT 291.980 52.740 293.370 52.930 ;
        RECT 295.185 52.830 295.415 53.820 ;
        RECT 291.440 52.280 292.000 52.570 ;
        RECT 292.170 52.110 292.420 52.570 ;
        RECT 293.040 52.380 293.370 52.740 ;
        RECT 294.665 52.660 295.415 52.830 ;
        RECT 294.665 52.370 294.920 52.660 ;
        RECT 295.090 52.110 295.420 52.490 ;
        RECT 295.590 52.370 295.760 54.490 ;
        RECT 295.930 53.690 296.255 54.475 ;
        RECT 296.425 54.200 296.675 54.660 ;
        RECT 296.845 54.160 297.095 54.490 ;
        RECT 297.310 54.160 297.990 54.490 ;
        RECT 296.845 54.030 297.015 54.160 ;
        RECT 296.620 53.860 297.015 54.030 ;
        RECT 295.990 52.640 296.450 53.690 ;
        RECT 296.620 52.500 296.790 53.860 ;
        RECT 297.185 53.600 297.650 53.990 ;
        RECT 296.960 52.790 297.310 53.410 ;
        RECT 297.480 53.010 297.650 53.600 ;
        RECT 297.820 53.380 297.990 54.160 ;
        RECT 298.160 54.060 298.330 54.400 ;
        RECT 298.565 54.230 298.895 54.660 ;
        RECT 299.065 54.060 299.235 54.400 ;
        RECT 299.530 54.200 299.900 54.660 ;
        RECT 298.160 53.890 299.235 54.060 ;
        RECT 300.070 54.030 300.240 54.490 ;
        RECT 300.475 54.150 301.345 54.490 ;
        RECT 301.515 54.200 301.765 54.660 ;
        RECT 299.680 53.860 300.240 54.030 ;
        RECT 299.680 53.720 299.850 53.860 ;
        RECT 298.350 53.550 299.850 53.720 ;
        RECT 300.545 53.690 301.005 53.980 ;
        RECT 297.820 53.210 299.510 53.380 ;
        RECT 297.480 52.790 297.835 53.010 ;
        RECT 298.005 52.500 298.175 53.210 ;
        RECT 298.380 52.790 299.170 53.040 ;
        RECT 299.340 53.030 299.510 53.210 ;
        RECT 299.680 52.860 299.850 53.550 ;
        RECT 296.120 52.110 296.450 52.470 ;
        RECT 296.620 52.330 297.115 52.500 ;
        RECT 297.320 52.330 298.175 52.500 ;
        RECT 299.050 52.110 299.380 52.570 ;
        RECT 299.590 52.470 299.850 52.860 ;
        RECT 300.040 53.680 301.005 53.690 ;
        RECT 301.175 53.770 301.345 54.150 ;
        RECT 301.935 54.110 302.105 54.400 ;
        RECT 302.285 54.280 302.615 54.660 ;
        RECT 301.935 53.940 302.735 54.110 ;
        RECT 300.040 53.520 300.715 53.680 ;
        RECT 301.175 53.600 302.395 53.770 ;
        RECT 300.040 52.730 300.250 53.520 ;
        RECT 301.175 53.510 301.345 53.600 ;
        RECT 300.420 52.730 300.770 53.350 ;
        RECT 300.940 53.340 301.345 53.510 ;
        RECT 300.940 52.560 301.110 53.340 ;
        RECT 301.280 52.890 301.500 53.170 ;
        RECT 301.680 53.060 302.220 53.430 ;
        RECT 302.565 53.350 302.735 53.940 ;
        RECT 302.955 53.520 303.260 54.660 ;
        RECT 303.430 53.470 303.685 54.350 ;
        RECT 303.860 53.495 304.150 54.660 ;
        RECT 304.320 53.570 305.990 54.660 ;
        RECT 302.565 53.320 303.305 53.350 ;
        RECT 301.280 52.720 301.810 52.890 ;
        RECT 299.590 52.300 299.940 52.470 ;
        RECT 300.160 52.280 301.110 52.560 ;
        RECT 301.280 52.110 301.470 52.550 ;
        RECT 301.640 52.490 301.810 52.720 ;
        RECT 301.980 52.660 302.220 53.060 ;
        RECT 302.390 53.020 303.305 53.320 ;
        RECT 302.390 52.845 302.715 53.020 ;
        RECT 302.390 52.490 302.710 52.845 ;
        RECT 303.475 52.820 303.685 53.470 ;
        RECT 304.320 52.880 305.070 53.400 ;
        RECT 305.240 53.050 305.990 53.570 ;
        RECT 306.160 53.520 306.545 54.490 ;
        RECT 306.715 54.200 307.040 54.660 ;
        RECT 307.560 54.030 307.840 54.490 ;
        RECT 306.715 53.810 307.840 54.030 ;
        RECT 301.640 52.320 302.710 52.490 ;
        RECT 302.955 52.110 303.260 52.570 ;
        RECT 303.430 52.290 303.685 52.820 ;
        RECT 303.860 52.110 304.150 52.835 ;
        RECT 304.320 52.110 305.990 52.880 ;
        RECT 306.160 52.850 306.440 53.520 ;
        RECT 306.715 53.350 307.165 53.810 ;
        RECT 308.030 53.640 308.430 54.490 ;
        RECT 308.830 54.200 309.100 54.660 ;
        RECT 309.270 54.030 309.555 54.490 ;
        RECT 306.610 53.020 307.165 53.350 ;
        RECT 307.335 53.080 308.430 53.640 ;
        RECT 306.715 52.910 307.165 53.020 ;
        RECT 306.160 52.280 306.545 52.850 ;
        RECT 306.715 52.740 307.840 52.910 ;
        RECT 306.715 52.110 307.040 52.570 ;
        RECT 307.560 52.280 307.840 52.740 ;
        RECT 308.030 52.280 308.430 53.080 ;
        RECT 308.600 53.810 309.555 54.030 ;
        RECT 308.600 52.910 308.810 53.810 ;
        RECT 308.980 53.080 309.670 53.640 ;
        RECT 309.840 53.570 311.050 54.660 ;
        RECT 309.840 53.030 310.360 53.570 ;
        RECT 308.600 52.740 309.555 52.910 ;
        RECT 310.530 52.860 311.050 53.400 ;
        RECT 308.830 52.110 309.100 52.570 ;
        RECT 309.270 52.280 309.555 52.740 ;
        RECT 309.840 52.110 311.050 52.860 ;
        RECT 162.095 51.940 311.135 52.110 ;
        RECT 162.180 51.190 163.390 51.940 ;
        RECT 163.560 51.395 168.905 51.940 ;
        RECT 169.080 51.395 174.425 51.940 ;
        RECT 174.600 51.395 179.945 51.940 ;
        RECT 180.120 51.395 185.465 51.940 ;
        RECT 162.180 50.650 162.700 51.190 ;
        RECT 162.870 50.480 163.390 51.020 ;
        RECT 165.145 50.565 165.485 51.395 ;
        RECT 162.180 49.390 163.390 50.480 ;
        RECT 166.965 49.825 167.315 51.075 ;
        RECT 170.665 50.565 171.005 51.395 ;
        RECT 172.485 49.825 172.835 51.075 ;
        RECT 176.185 50.565 176.525 51.395 ;
        RECT 178.005 49.825 178.355 51.075 ;
        RECT 181.705 50.565 182.045 51.395 ;
        RECT 185.640 51.170 187.310 51.940 ;
        RECT 187.940 51.215 188.230 51.940 ;
        RECT 188.400 51.190 189.610 51.940 ;
        RECT 190.025 51.460 190.325 51.940 ;
        RECT 190.495 51.290 190.755 51.745 ;
        RECT 190.925 51.460 191.185 51.940 ;
        RECT 191.355 51.290 191.615 51.745 ;
        RECT 191.785 51.460 192.045 51.940 ;
        RECT 192.215 51.290 192.475 51.745 ;
        RECT 192.645 51.460 192.905 51.940 ;
        RECT 193.075 51.290 193.335 51.745 ;
        RECT 193.505 51.415 193.765 51.940 ;
        RECT 183.525 49.825 183.875 51.075 ;
        RECT 185.640 50.650 186.390 51.170 ;
        RECT 186.560 50.480 187.310 51.000 ;
        RECT 188.400 50.650 188.920 51.190 ;
        RECT 190.025 51.120 193.335 51.290 ;
        RECT 163.560 49.390 168.905 49.825 ;
        RECT 169.080 49.390 174.425 49.825 ;
        RECT 174.600 49.390 179.945 49.825 ;
        RECT 180.120 49.390 185.465 49.825 ;
        RECT 185.640 49.390 187.310 50.480 ;
        RECT 187.940 49.390 188.230 50.555 ;
        RECT 189.090 50.480 189.610 51.020 ;
        RECT 188.400 49.390 189.610 50.480 ;
        RECT 190.025 50.530 190.995 51.120 ;
        RECT 193.935 50.950 194.185 51.760 ;
        RECT 194.365 51.480 194.610 51.940 ;
        RECT 191.165 50.700 194.185 50.950 ;
        RECT 194.355 50.700 194.670 51.310 ;
        RECT 194.840 51.170 198.350 51.940 ;
        RECT 199.070 51.390 199.240 51.770 ;
        RECT 199.420 51.560 199.750 51.940 ;
        RECT 199.070 51.220 199.735 51.390 ;
        RECT 199.930 51.265 200.190 51.770 ;
        RECT 190.025 50.290 193.335 50.530 ;
        RECT 190.030 49.390 190.325 50.120 ;
        RECT 190.495 49.565 190.755 50.290 ;
        RECT 190.925 49.390 191.185 50.120 ;
        RECT 191.355 49.565 191.615 50.290 ;
        RECT 191.785 49.390 192.045 50.120 ;
        RECT 192.215 49.565 192.475 50.290 ;
        RECT 192.645 49.390 192.905 50.120 ;
        RECT 193.075 49.565 193.335 50.290 ;
        RECT 193.505 49.390 193.765 50.500 ;
        RECT 193.935 49.565 194.185 50.700 ;
        RECT 194.840 50.650 196.490 51.170 ;
        RECT 194.365 49.390 194.660 50.500 ;
        RECT 196.660 50.480 198.350 51.000 ;
        RECT 199.000 50.670 199.330 51.040 ;
        RECT 199.565 50.965 199.735 51.220 ;
        RECT 199.565 50.635 199.850 50.965 ;
        RECT 199.565 50.490 199.735 50.635 ;
        RECT 194.840 49.390 198.350 50.480 ;
        RECT 199.070 50.320 199.735 50.490 ;
        RECT 200.020 50.465 200.190 51.265 ;
        RECT 200.360 51.200 200.620 51.940 ;
        RECT 200.870 51.120 201.060 51.590 ;
        RECT 201.310 51.440 201.560 51.940 ;
        RECT 201.890 51.370 202.060 51.720 ;
        RECT 202.260 51.540 202.590 51.940 ;
        RECT 202.760 51.370 202.930 51.720 ;
        RECT 203.150 51.540 203.530 51.940 ;
        RECT 200.890 51.030 201.060 51.120 ;
        RECT 201.730 51.200 203.540 51.370 ;
        RECT 199.070 49.560 199.240 50.320 ;
        RECT 199.420 49.390 199.750 50.150 ;
        RECT 199.920 49.560 200.190 50.465 ;
        RECT 200.380 50.070 200.720 51.030 ;
        RECT 200.890 50.700 201.490 51.030 ;
        RECT 200.890 49.960 201.060 50.700 ;
        RECT 201.730 50.450 201.900 51.200 ;
        RECT 200.360 49.390 200.640 49.890 ;
        RECT 200.870 49.570 201.060 49.960 ;
        RECT 201.310 50.280 201.900 50.450 ;
        RECT 202.070 50.405 202.240 51.030 ;
        RECT 202.470 50.575 202.800 51.030 ;
        RECT 201.310 49.575 201.640 50.280 ;
        RECT 202.070 49.650 202.430 50.405 ;
        RECT 202.610 50.240 202.800 50.575 ;
        RECT 203.030 50.580 203.200 51.030 ;
        RECT 203.370 50.950 203.540 51.200 ;
        RECT 203.710 51.300 203.960 51.770 ;
        RECT 204.130 51.470 204.300 51.940 ;
        RECT 204.470 51.300 204.800 51.770 ;
        RECT 204.970 51.470 205.140 51.940 ;
        RECT 203.710 51.120 205.240 51.300 ;
        RECT 203.370 50.780 204.830 50.950 ;
        RECT 203.030 50.410 203.465 50.580 ;
        RECT 205.000 50.570 205.240 51.120 ;
        RECT 203.670 50.400 205.240 50.570 ;
        RECT 205.425 51.200 205.680 51.770 ;
        RECT 205.850 51.540 206.180 51.940 ;
        RECT 206.605 51.405 207.135 51.770 ;
        RECT 207.325 51.600 207.600 51.770 ;
        RECT 207.320 51.430 207.600 51.600 ;
        RECT 206.605 51.370 206.780 51.405 ;
        RECT 205.850 51.200 206.780 51.370 ;
        RECT 205.425 50.530 205.595 51.200 ;
        RECT 205.850 51.030 206.020 51.200 ;
        RECT 205.765 50.700 206.020 51.030 ;
        RECT 206.245 50.700 206.440 51.030 ;
        RECT 202.610 49.650 202.910 50.240 ;
        RECT 203.195 49.390 203.445 50.230 ;
        RECT 203.670 49.560 203.920 50.400 ;
        RECT 204.090 49.390 204.340 50.230 ;
        RECT 204.510 49.560 204.760 50.400 ;
        RECT 204.930 49.390 205.180 50.230 ;
        RECT 205.425 49.560 205.760 50.530 ;
        RECT 205.930 49.390 206.100 50.530 ;
        RECT 206.270 49.730 206.440 50.700 ;
        RECT 206.610 50.070 206.780 51.200 ;
        RECT 206.950 50.410 207.120 51.210 ;
        RECT 207.325 50.610 207.600 51.430 ;
        RECT 207.770 50.410 207.960 51.770 ;
        RECT 208.140 51.405 208.650 51.940 ;
        RECT 208.870 51.130 209.115 51.735 ;
        RECT 209.645 51.440 210.140 51.770 ;
        RECT 208.160 50.960 209.390 51.130 ;
        RECT 206.950 50.240 207.960 50.410 ;
        RECT 208.130 50.395 208.880 50.585 ;
        RECT 206.610 49.900 207.735 50.070 ;
        RECT 208.130 49.730 208.300 50.395 ;
        RECT 209.050 50.150 209.390 50.960 ;
        RECT 206.270 49.560 208.300 49.730 ;
        RECT 208.470 49.390 208.640 50.150 ;
        RECT 208.875 49.740 209.390 50.150 ;
        RECT 209.560 49.950 209.800 51.260 ;
        RECT 209.970 50.530 210.140 51.440 ;
        RECT 210.360 50.700 210.710 51.665 ;
        RECT 210.890 50.700 211.190 51.670 ;
        RECT 211.370 50.700 211.650 51.670 ;
        RECT 211.830 51.140 212.100 51.940 ;
        RECT 212.270 51.220 212.610 51.730 ;
        RECT 211.845 50.700 212.175 50.950 ;
        RECT 211.845 50.530 212.160 50.700 ;
        RECT 209.970 50.360 212.160 50.530 ;
        RECT 209.565 49.390 209.900 49.770 ;
        RECT 210.070 49.560 210.320 50.360 ;
        RECT 210.540 49.390 210.870 50.110 ;
        RECT 211.055 49.560 211.305 50.360 ;
        RECT 211.770 49.390 212.100 50.190 ;
        RECT 212.350 49.820 212.610 51.220 ;
        RECT 213.700 51.215 213.990 51.940 ;
        RECT 214.245 51.370 214.420 51.770 ;
        RECT 214.590 51.560 214.920 51.940 ;
        RECT 215.165 51.440 215.395 51.770 ;
        RECT 214.245 51.200 214.875 51.370 ;
        RECT 214.705 51.030 214.875 51.200 ;
        RECT 212.270 49.560 212.610 49.820 ;
        RECT 213.700 49.390 213.990 50.555 ;
        RECT 214.160 50.350 214.525 51.030 ;
        RECT 214.705 50.700 215.055 51.030 ;
        RECT 214.705 50.180 214.875 50.700 ;
        RECT 214.245 50.010 214.875 50.180 ;
        RECT 215.225 50.150 215.395 51.440 ;
        RECT 215.595 50.330 215.875 51.605 ;
        RECT 216.100 50.580 216.370 51.605 ;
        RECT 216.830 51.560 217.160 51.940 ;
        RECT 217.330 51.685 217.665 51.730 ;
        RECT 216.060 50.410 216.370 50.580 ;
        RECT 216.100 50.330 216.370 50.410 ;
        RECT 216.560 50.330 216.900 51.360 ;
        RECT 217.330 51.220 217.670 51.685 ;
        RECT 218.085 51.460 218.385 51.940 ;
        RECT 218.555 51.290 218.815 51.745 ;
        RECT 218.985 51.460 219.245 51.940 ;
        RECT 219.415 51.290 219.675 51.745 ;
        RECT 219.845 51.460 220.105 51.940 ;
        RECT 220.275 51.290 220.535 51.745 ;
        RECT 220.705 51.460 220.965 51.940 ;
        RECT 221.135 51.290 221.395 51.745 ;
        RECT 221.565 51.415 221.825 51.940 ;
        RECT 217.070 50.700 217.330 51.030 ;
        RECT 217.070 50.150 217.240 50.700 ;
        RECT 217.500 50.530 217.670 51.220 ;
        RECT 214.245 49.560 214.420 50.010 ;
        RECT 215.225 49.980 217.240 50.150 ;
        RECT 214.590 49.390 214.920 49.830 ;
        RECT 215.225 49.560 215.395 49.980 ;
        RECT 215.630 49.390 216.300 49.800 ;
        RECT 216.515 49.560 216.685 49.980 ;
        RECT 216.885 49.390 217.215 49.800 ;
        RECT 217.410 49.560 217.670 50.530 ;
        RECT 218.085 51.120 221.395 51.290 ;
        RECT 218.085 50.530 219.055 51.120 ;
        RECT 221.995 50.950 222.245 51.760 ;
        RECT 222.425 51.480 222.670 51.940 ;
        RECT 219.225 50.700 222.245 50.950 ;
        RECT 222.415 50.700 222.730 51.310 ;
        RECT 222.900 51.170 224.570 51.940 ;
        RECT 224.745 51.390 225.000 51.680 ;
        RECT 225.170 51.560 225.500 51.940 ;
        RECT 224.745 51.220 225.495 51.390 ;
        RECT 218.085 50.290 221.395 50.530 ;
        RECT 218.090 49.390 218.385 50.120 ;
        RECT 218.555 49.565 218.815 50.290 ;
        RECT 218.985 49.390 219.245 50.120 ;
        RECT 219.415 49.565 219.675 50.290 ;
        RECT 219.845 49.390 220.105 50.120 ;
        RECT 220.275 49.565 220.535 50.290 ;
        RECT 220.705 49.390 220.965 50.120 ;
        RECT 221.135 49.565 221.395 50.290 ;
        RECT 221.565 49.390 221.825 50.500 ;
        RECT 221.995 49.565 222.245 50.700 ;
        RECT 222.900 50.650 223.650 51.170 ;
        RECT 222.425 49.390 222.720 50.500 ;
        RECT 223.820 50.480 224.570 51.000 ;
        RECT 222.900 49.390 224.570 50.480 ;
        RECT 224.745 50.400 225.095 51.050 ;
        RECT 225.265 50.230 225.495 51.220 ;
        RECT 224.745 50.060 225.495 50.230 ;
        RECT 224.745 49.560 225.000 50.060 ;
        RECT 225.170 49.390 225.500 49.890 ;
        RECT 225.670 49.560 225.840 51.680 ;
        RECT 226.200 51.580 226.530 51.940 ;
        RECT 226.700 51.550 227.195 51.720 ;
        RECT 227.400 51.550 228.255 51.720 ;
        RECT 226.070 50.360 226.530 51.410 ;
        RECT 226.010 49.575 226.335 50.360 ;
        RECT 226.700 50.190 226.870 51.550 ;
        RECT 227.040 50.640 227.390 51.260 ;
        RECT 227.560 51.040 227.915 51.260 ;
        RECT 227.560 50.450 227.730 51.040 ;
        RECT 228.085 50.840 228.255 51.550 ;
        RECT 229.130 51.480 229.460 51.940 ;
        RECT 229.670 51.580 230.020 51.750 ;
        RECT 228.460 51.010 229.250 51.260 ;
        RECT 229.670 51.190 229.930 51.580 ;
        RECT 230.240 51.490 231.190 51.770 ;
        RECT 231.360 51.500 231.550 51.940 ;
        RECT 231.720 51.560 232.790 51.730 ;
        RECT 229.420 50.840 229.590 51.020 ;
        RECT 226.700 50.020 227.095 50.190 ;
        RECT 227.265 50.060 227.730 50.450 ;
        RECT 227.900 50.670 229.590 50.840 ;
        RECT 226.925 49.890 227.095 50.020 ;
        RECT 227.900 49.890 228.070 50.670 ;
        RECT 229.760 50.500 229.930 51.190 ;
        RECT 228.430 50.330 229.930 50.500 ;
        RECT 230.120 50.530 230.330 51.320 ;
        RECT 230.500 50.700 230.850 51.320 ;
        RECT 231.020 50.710 231.190 51.490 ;
        RECT 231.720 51.330 231.890 51.560 ;
        RECT 231.360 51.160 231.890 51.330 ;
        RECT 231.360 50.880 231.580 51.160 ;
        RECT 232.060 50.990 232.300 51.390 ;
        RECT 231.020 50.540 231.425 50.710 ;
        RECT 231.760 50.620 232.300 50.990 ;
        RECT 232.470 51.205 232.790 51.560 ;
        RECT 233.035 51.480 233.340 51.940 ;
        RECT 233.510 51.230 233.765 51.760 ;
        RECT 232.470 51.030 232.795 51.205 ;
        RECT 232.470 50.730 233.385 51.030 ;
        RECT 232.645 50.700 233.385 50.730 ;
        RECT 230.120 50.370 230.795 50.530 ;
        RECT 231.255 50.450 231.425 50.540 ;
        RECT 230.120 50.360 231.085 50.370 ;
        RECT 229.760 50.190 229.930 50.330 ;
        RECT 226.505 49.390 226.755 49.850 ;
        RECT 226.925 49.560 227.175 49.890 ;
        RECT 227.390 49.560 228.070 49.890 ;
        RECT 228.240 49.990 229.315 50.160 ;
        RECT 229.760 50.020 230.320 50.190 ;
        RECT 230.625 50.070 231.085 50.360 ;
        RECT 231.255 50.280 232.475 50.450 ;
        RECT 228.240 49.650 228.410 49.990 ;
        RECT 228.645 49.390 228.975 49.820 ;
        RECT 229.145 49.650 229.315 49.990 ;
        RECT 229.610 49.390 229.980 49.850 ;
        RECT 230.150 49.560 230.320 50.020 ;
        RECT 231.255 49.900 231.425 50.280 ;
        RECT 232.645 50.110 232.815 50.700 ;
        RECT 233.555 50.580 233.765 51.230 ;
        RECT 233.940 51.170 235.610 51.940 ;
        RECT 236.240 51.330 236.580 51.745 ;
        RECT 236.750 51.500 236.920 51.940 ;
        RECT 237.090 51.550 238.340 51.730 ;
        RECT 237.090 51.330 237.420 51.550 ;
        RECT 238.610 51.480 238.780 51.940 ;
        RECT 233.940 50.650 234.690 51.170 ;
        RECT 236.240 51.160 237.420 51.330 ;
        RECT 237.590 51.310 237.955 51.380 ;
        RECT 237.590 51.130 238.840 51.310 ;
        RECT 230.555 49.560 231.425 49.900 ;
        RECT 232.015 49.940 232.815 50.110 ;
        RECT 231.595 49.390 231.845 49.850 ;
        RECT 232.015 49.650 232.185 49.940 ;
        RECT 232.365 49.390 232.695 49.770 ;
        RECT 233.035 49.390 233.340 50.530 ;
        RECT 233.510 49.700 233.765 50.580 ;
        RECT 234.860 50.480 235.610 51.000 ;
        RECT 236.240 50.750 236.705 50.950 ;
        RECT 236.880 50.700 237.210 50.950 ;
        RECT 237.380 50.920 237.845 50.950 ;
        RECT 237.380 50.750 237.850 50.920 ;
        RECT 237.380 50.700 237.845 50.750 ;
        RECT 238.040 50.700 238.395 50.950 ;
        RECT 236.880 50.580 237.060 50.700 ;
        RECT 233.940 49.390 235.610 50.480 ;
        RECT 236.240 49.390 236.560 50.570 ;
        RECT 236.730 50.410 237.060 50.580 ;
        RECT 238.565 50.530 238.840 51.130 ;
        RECT 236.730 49.620 236.930 50.410 ;
        RECT 237.230 50.320 238.840 50.530 ;
        RECT 237.230 50.220 237.640 50.320 ;
        RECT 237.255 49.560 237.640 50.220 ;
        RECT 238.035 49.390 238.820 50.150 ;
        RECT 239.010 49.560 239.290 51.660 ;
        RECT 239.460 51.215 239.750 51.940 ;
        RECT 239.920 51.200 240.305 51.770 ;
        RECT 240.475 51.480 240.800 51.940 ;
        RECT 241.320 51.310 241.600 51.770 ;
        RECT 239.460 49.390 239.750 50.555 ;
        RECT 239.920 50.530 240.200 51.200 ;
        RECT 240.475 51.140 241.600 51.310 ;
        RECT 240.475 51.030 240.925 51.140 ;
        RECT 240.370 50.700 240.925 51.030 ;
        RECT 241.790 50.970 242.190 51.770 ;
        RECT 242.590 51.480 242.860 51.940 ;
        RECT 243.030 51.310 243.315 51.770 ;
        RECT 239.920 49.560 240.305 50.530 ;
        RECT 240.475 50.240 240.925 50.700 ;
        RECT 241.095 50.410 242.190 50.970 ;
        RECT 240.475 50.020 241.600 50.240 ;
        RECT 240.475 49.390 240.800 49.850 ;
        RECT 241.320 49.560 241.600 50.020 ;
        RECT 241.790 49.560 242.190 50.410 ;
        RECT 242.360 51.140 243.315 51.310 ;
        RECT 243.600 51.170 245.270 51.940 ;
        RECT 245.440 51.200 245.825 51.770 ;
        RECT 245.995 51.480 246.320 51.940 ;
        RECT 246.840 51.310 247.120 51.770 ;
        RECT 242.360 50.240 242.570 51.140 ;
        RECT 242.740 50.410 243.430 50.970 ;
        RECT 243.600 50.650 244.350 51.170 ;
        RECT 244.520 50.480 245.270 51.000 ;
        RECT 242.360 50.020 243.315 50.240 ;
        RECT 242.590 49.390 242.860 49.850 ;
        RECT 243.030 49.560 243.315 50.020 ;
        RECT 243.600 49.390 245.270 50.480 ;
        RECT 245.440 50.530 245.720 51.200 ;
        RECT 245.995 51.140 247.120 51.310 ;
        RECT 245.995 51.030 246.445 51.140 ;
        RECT 245.890 50.700 246.445 51.030 ;
        RECT 247.310 50.970 247.710 51.770 ;
        RECT 248.110 51.480 248.380 51.940 ;
        RECT 248.550 51.310 248.835 51.770 ;
        RECT 249.120 51.395 254.465 51.940 ;
        RECT 254.885 51.460 255.185 51.940 ;
        RECT 245.440 49.560 245.825 50.530 ;
        RECT 245.995 50.240 246.445 50.700 ;
        RECT 246.615 50.410 247.710 50.970 ;
        RECT 245.995 50.020 247.120 50.240 ;
        RECT 245.995 49.390 246.320 49.850 ;
        RECT 246.840 49.560 247.120 50.020 ;
        RECT 247.310 49.560 247.710 50.410 ;
        RECT 247.880 51.140 248.835 51.310 ;
        RECT 247.880 50.240 248.090 51.140 ;
        RECT 248.260 50.410 248.950 50.970 ;
        RECT 250.705 50.565 251.045 51.395 ;
        RECT 255.355 51.290 255.615 51.745 ;
        RECT 255.785 51.460 256.045 51.940 ;
        RECT 256.215 51.290 256.475 51.745 ;
        RECT 256.645 51.460 256.905 51.940 ;
        RECT 257.075 51.290 257.335 51.745 ;
        RECT 257.505 51.460 257.765 51.940 ;
        RECT 257.935 51.290 258.195 51.745 ;
        RECT 258.365 51.415 258.625 51.940 ;
        RECT 254.885 51.120 258.195 51.290 ;
        RECT 247.880 50.020 248.835 50.240 ;
        RECT 248.110 49.390 248.380 49.850 ;
        RECT 248.550 49.560 248.835 50.020 ;
        RECT 252.525 49.825 252.875 51.075 ;
        RECT 254.885 50.530 255.855 51.120 ;
        RECT 258.795 50.950 259.045 51.760 ;
        RECT 259.225 51.480 259.470 51.940 ;
        RECT 256.025 50.700 259.045 50.950 ;
        RECT 259.215 50.700 259.530 51.310 ;
        RECT 259.700 51.200 260.040 51.770 ;
        RECT 260.235 51.275 260.405 51.940 ;
        RECT 260.685 51.600 260.905 51.645 ;
        RECT 260.680 51.430 260.905 51.600 ;
        RECT 261.075 51.460 261.520 51.630 ;
        RECT 260.685 51.290 260.905 51.430 ;
        RECT 254.885 50.290 258.195 50.530 ;
        RECT 249.120 49.390 254.465 49.825 ;
        RECT 254.890 49.390 255.185 50.120 ;
        RECT 255.355 49.565 255.615 50.290 ;
        RECT 255.785 49.390 256.045 50.120 ;
        RECT 256.215 49.565 256.475 50.290 ;
        RECT 256.645 49.390 256.905 50.120 ;
        RECT 257.075 49.565 257.335 50.290 ;
        RECT 257.505 49.390 257.765 50.120 ;
        RECT 257.935 49.565 258.195 50.290 ;
        RECT 258.365 49.390 258.625 50.500 ;
        RECT 258.795 49.565 259.045 50.700 ;
        RECT 259.225 49.390 259.520 50.500 ;
        RECT 259.700 50.230 259.875 51.200 ;
        RECT 260.685 51.120 261.180 51.290 ;
        RECT 260.045 50.580 260.215 51.030 ;
        RECT 260.385 50.750 260.835 50.950 ;
        RECT 261.005 50.925 261.180 51.120 ;
        RECT 261.350 50.670 261.520 51.460 ;
        RECT 261.690 51.335 261.940 51.705 ;
        RECT 261.770 50.950 261.940 51.335 ;
        RECT 262.110 51.300 262.360 51.705 ;
        RECT 262.530 51.470 262.700 51.940 ;
        RECT 262.870 51.300 263.210 51.705 ;
        RECT 262.110 51.120 263.210 51.300 ;
        RECT 263.380 51.170 265.050 51.940 ;
        RECT 265.220 51.215 265.510 51.940 ;
        RECT 265.685 51.390 265.940 51.680 ;
        RECT 266.110 51.560 266.440 51.940 ;
        RECT 265.685 51.220 266.435 51.390 ;
        RECT 261.770 50.780 261.965 50.950 ;
        RECT 260.045 50.410 260.440 50.580 ;
        RECT 261.350 50.530 261.625 50.670 ;
        RECT 259.700 49.560 259.960 50.230 ;
        RECT 260.270 50.140 260.440 50.410 ;
        RECT 260.610 50.310 261.625 50.530 ;
        RECT 261.795 50.530 261.965 50.780 ;
        RECT 262.135 50.700 262.695 50.950 ;
        RECT 261.795 50.140 262.350 50.530 ;
        RECT 260.270 49.970 262.350 50.140 ;
        RECT 260.130 49.390 260.460 49.790 ;
        RECT 261.330 49.390 261.730 49.790 ;
        RECT 262.020 49.735 262.350 49.970 ;
        RECT 262.520 49.600 262.695 50.700 ;
        RECT 262.865 50.380 263.210 50.950 ;
        RECT 263.380 50.650 264.130 51.170 ;
        RECT 264.300 50.480 265.050 51.000 ;
        RECT 262.865 49.390 263.210 50.210 ;
        RECT 263.380 49.390 265.050 50.480 ;
        RECT 265.220 49.390 265.510 50.555 ;
        RECT 265.685 50.400 266.035 51.050 ;
        RECT 266.205 50.230 266.435 51.220 ;
        RECT 265.685 50.060 266.435 50.230 ;
        RECT 265.685 49.560 265.940 50.060 ;
        RECT 266.110 49.390 266.440 49.890 ;
        RECT 266.610 49.560 266.780 51.680 ;
        RECT 267.140 51.580 267.470 51.940 ;
        RECT 267.640 51.550 268.135 51.720 ;
        RECT 268.340 51.550 269.195 51.720 ;
        RECT 267.010 50.360 267.470 51.410 ;
        RECT 266.950 49.575 267.275 50.360 ;
        RECT 267.640 50.190 267.810 51.550 ;
        RECT 267.980 50.640 268.330 51.260 ;
        RECT 268.500 51.040 268.855 51.260 ;
        RECT 268.500 50.450 268.670 51.040 ;
        RECT 269.025 50.840 269.195 51.550 ;
        RECT 270.070 51.480 270.400 51.940 ;
        RECT 270.610 51.580 270.960 51.750 ;
        RECT 269.400 51.010 270.190 51.260 ;
        RECT 270.610 51.190 270.870 51.580 ;
        RECT 271.180 51.490 272.130 51.770 ;
        RECT 272.300 51.500 272.490 51.940 ;
        RECT 272.660 51.560 273.730 51.730 ;
        RECT 270.360 50.840 270.530 51.020 ;
        RECT 267.640 50.020 268.035 50.190 ;
        RECT 268.205 50.060 268.670 50.450 ;
        RECT 268.840 50.670 270.530 50.840 ;
        RECT 267.865 49.890 268.035 50.020 ;
        RECT 268.840 49.890 269.010 50.670 ;
        RECT 270.700 50.500 270.870 51.190 ;
        RECT 269.370 50.330 270.870 50.500 ;
        RECT 271.060 50.530 271.270 51.320 ;
        RECT 271.440 50.700 271.790 51.320 ;
        RECT 271.960 50.710 272.130 51.490 ;
        RECT 272.660 51.330 272.830 51.560 ;
        RECT 272.300 51.160 272.830 51.330 ;
        RECT 272.300 50.880 272.520 51.160 ;
        RECT 273.000 50.990 273.240 51.390 ;
        RECT 271.960 50.540 272.365 50.710 ;
        RECT 272.700 50.620 273.240 50.990 ;
        RECT 273.410 51.205 273.730 51.560 ;
        RECT 273.975 51.480 274.280 51.940 ;
        RECT 274.450 51.230 274.705 51.760 ;
        RECT 273.410 51.030 273.735 51.205 ;
        RECT 273.410 50.730 274.325 51.030 ;
        RECT 273.585 50.700 274.325 50.730 ;
        RECT 271.060 50.370 271.735 50.530 ;
        RECT 272.195 50.450 272.365 50.540 ;
        RECT 271.060 50.360 272.025 50.370 ;
        RECT 270.700 50.190 270.870 50.330 ;
        RECT 267.445 49.390 267.695 49.850 ;
        RECT 267.865 49.560 268.115 49.890 ;
        RECT 268.330 49.560 269.010 49.890 ;
        RECT 269.180 49.990 270.255 50.160 ;
        RECT 270.700 50.020 271.260 50.190 ;
        RECT 271.565 50.070 272.025 50.360 ;
        RECT 272.195 50.280 273.415 50.450 ;
        RECT 269.180 49.650 269.350 49.990 ;
        RECT 269.585 49.390 269.915 49.820 ;
        RECT 270.085 49.650 270.255 49.990 ;
        RECT 270.550 49.390 270.920 49.850 ;
        RECT 271.090 49.560 271.260 50.020 ;
        RECT 272.195 49.900 272.365 50.280 ;
        RECT 273.585 50.110 273.755 50.700 ;
        RECT 274.495 50.580 274.705 51.230 ;
        RECT 275.080 51.310 275.410 51.670 ;
        RECT 276.030 51.480 276.280 51.940 ;
        RECT 276.450 51.480 277.010 51.770 ;
        RECT 275.080 51.120 276.470 51.310 ;
        RECT 276.300 51.030 276.470 51.120 ;
        RECT 271.495 49.560 272.365 49.900 ;
        RECT 272.955 49.940 273.755 50.110 ;
        RECT 272.535 49.390 272.785 49.850 ;
        RECT 272.955 49.650 273.125 49.940 ;
        RECT 273.305 49.390 273.635 49.770 ;
        RECT 273.975 49.390 274.280 50.530 ;
        RECT 274.450 49.700 274.705 50.580 ;
        RECT 274.895 50.700 275.570 50.950 ;
        RECT 275.790 50.700 276.130 50.950 ;
        RECT 276.300 50.700 276.590 51.030 ;
        RECT 274.895 50.340 275.160 50.700 ;
        RECT 276.300 50.450 276.470 50.700 ;
        RECT 275.530 50.280 276.470 50.450 ;
        RECT 275.080 49.390 275.360 50.060 ;
        RECT 275.530 49.730 275.830 50.280 ;
        RECT 276.760 50.110 277.010 51.480 ;
        RECT 277.295 51.310 277.580 51.770 ;
        RECT 277.750 51.480 278.020 51.940 ;
        RECT 277.295 51.140 278.250 51.310 ;
        RECT 277.180 50.410 277.870 50.970 ;
        RECT 278.040 50.240 278.250 51.140 ;
        RECT 276.030 49.390 276.360 50.110 ;
        RECT 276.550 49.560 277.010 50.110 ;
        RECT 277.295 50.020 278.250 50.240 ;
        RECT 278.420 50.970 278.820 51.770 ;
        RECT 279.010 51.310 279.290 51.770 ;
        RECT 279.810 51.480 280.135 51.940 ;
        RECT 279.010 51.140 280.135 51.310 ;
        RECT 280.305 51.200 280.690 51.770 ;
        RECT 279.685 51.030 280.135 51.140 ;
        RECT 278.420 50.410 279.515 50.970 ;
        RECT 279.685 50.700 280.240 51.030 ;
        RECT 277.295 49.560 277.580 50.020 ;
        RECT 277.750 49.390 278.020 49.850 ;
        RECT 278.420 49.560 278.820 50.410 ;
        RECT 279.685 50.240 280.135 50.700 ;
        RECT 280.410 50.530 280.690 51.200 ;
        RECT 280.950 51.290 281.120 51.770 ;
        RECT 281.290 51.460 281.620 51.940 ;
        RECT 281.845 51.520 283.380 51.770 ;
        RECT 281.845 51.290 282.015 51.520 ;
        RECT 280.950 51.120 282.015 51.290 ;
        RECT 282.195 50.950 282.475 51.350 ;
        RECT 280.865 50.740 281.215 50.950 ;
        RECT 281.385 50.750 281.830 50.950 ;
        RECT 282.000 50.750 282.475 50.950 ;
        RECT 282.745 50.950 283.030 51.350 ;
        RECT 283.210 51.290 283.380 51.520 ;
        RECT 283.550 51.460 283.880 51.940 ;
        RECT 284.095 51.440 284.350 51.770 ;
        RECT 284.600 51.480 284.845 51.940 ;
        RECT 284.165 51.360 284.350 51.440 ;
        RECT 283.210 51.120 284.010 51.290 ;
        RECT 282.745 50.750 283.075 50.950 ;
        RECT 283.245 50.750 283.610 50.950 ;
        RECT 283.840 50.570 284.010 51.120 ;
        RECT 279.010 50.020 280.135 50.240 ;
        RECT 279.010 49.560 279.290 50.020 ;
        RECT 279.810 49.390 280.135 49.850 ;
        RECT 280.305 49.560 280.690 50.530 ;
        RECT 280.950 50.400 284.010 50.570 ;
        RECT 280.950 49.560 281.120 50.400 ;
        RECT 284.180 50.240 284.350 51.360 ;
        RECT 284.540 50.700 284.855 51.310 ;
        RECT 285.025 50.950 285.275 51.760 ;
        RECT 285.445 51.415 285.705 51.940 ;
        RECT 285.875 51.290 286.135 51.745 ;
        RECT 286.305 51.460 286.565 51.940 ;
        RECT 286.735 51.290 286.995 51.745 ;
        RECT 287.165 51.460 287.425 51.940 ;
        RECT 287.595 51.290 287.855 51.745 ;
        RECT 288.025 51.460 288.285 51.940 ;
        RECT 288.455 51.290 288.715 51.745 ;
        RECT 288.885 51.460 289.185 51.940 ;
        RECT 285.875 51.120 289.185 51.290 ;
        RECT 285.025 50.700 288.045 50.950 ;
        RECT 284.140 50.230 284.350 50.240 ;
        RECT 281.290 49.730 281.620 50.230 ;
        RECT 281.790 49.990 283.425 50.230 ;
        RECT 281.790 49.900 282.020 49.990 ;
        RECT 282.130 49.730 282.460 49.770 ;
        RECT 281.290 49.560 282.460 49.730 ;
        RECT 282.650 49.390 283.005 49.810 ;
        RECT 283.175 49.560 283.425 49.990 ;
        RECT 283.595 49.390 283.925 50.150 ;
        RECT 284.095 49.560 284.350 50.230 ;
        RECT 284.550 49.390 284.845 50.500 ;
        RECT 285.025 49.565 285.275 50.700 ;
        RECT 288.215 50.530 289.185 51.120 ;
        RECT 289.600 51.190 290.810 51.940 ;
        RECT 290.980 51.215 291.270 51.940 ;
        RECT 291.555 51.310 291.840 51.770 ;
        RECT 292.010 51.480 292.280 51.940 ;
        RECT 289.600 50.650 290.120 51.190 ;
        RECT 291.555 51.140 292.510 51.310 ;
        RECT 285.445 49.390 285.705 50.500 ;
        RECT 285.875 50.290 289.185 50.530 ;
        RECT 290.290 50.480 290.810 51.020 ;
        RECT 285.875 49.565 286.135 50.290 ;
        RECT 286.305 49.390 286.565 50.120 ;
        RECT 286.735 49.565 286.995 50.290 ;
        RECT 287.165 49.390 287.425 50.120 ;
        RECT 287.595 49.565 287.855 50.290 ;
        RECT 288.025 49.390 288.285 50.120 ;
        RECT 288.455 49.565 288.715 50.290 ;
        RECT 288.885 49.390 289.180 50.120 ;
        RECT 289.600 49.390 290.810 50.480 ;
        RECT 290.980 49.390 291.270 50.555 ;
        RECT 291.440 50.410 292.130 50.970 ;
        RECT 292.300 50.240 292.510 51.140 ;
        RECT 291.555 50.020 292.510 50.240 ;
        RECT 292.680 50.970 293.080 51.770 ;
        RECT 293.270 51.310 293.550 51.770 ;
        RECT 294.070 51.480 294.395 51.940 ;
        RECT 293.270 51.140 294.395 51.310 ;
        RECT 294.565 51.200 294.950 51.770 ;
        RECT 293.945 51.030 294.395 51.140 ;
        RECT 292.680 50.410 293.775 50.970 ;
        RECT 293.945 50.700 294.500 51.030 ;
        RECT 291.555 49.560 291.840 50.020 ;
        RECT 292.010 49.390 292.280 49.850 ;
        RECT 292.680 49.560 293.080 50.410 ;
        RECT 293.945 50.240 294.395 50.700 ;
        RECT 294.670 50.530 294.950 51.200 ;
        RECT 293.270 50.020 294.395 50.240 ;
        RECT 293.270 49.560 293.550 50.020 ;
        RECT 294.070 49.390 294.395 49.850 ;
        RECT 294.565 49.560 294.950 50.530 ;
        RECT 295.585 51.200 295.840 51.770 ;
        RECT 296.010 51.540 296.340 51.940 ;
        RECT 296.765 51.405 297.295 51.770 ;
        RECT 297.485 51.600 297.760 51.770 ;
        RECT 297.480 51.430 297.760 51.600 ;
        RECT 296.765 51.370 296.940 51.405 ;
        RECT 296.010 51.200 296.940 51.370 ;
        RECT 295.585 50.530 295.755 51.200 ;
        RECT 296.010 51.030 296.180 51.200 ;
        RECT 295.925 50.700 296.180 51.030 ;
        RECT 296.405 50.700 296.600 51.030 ;
        RECT 295.585 49.560 295.920 50.530 ;
        RECT 296.090 49.390 296.260 50.530 ;
        RECT 296.430 49.730 296.600 50.700 ;
        RECT 296.770 50.070 296.940 51.200 ;
        RECT 297.110 50.410 297.280 51.210 ;
        RECT 297.485 50.610 297.760 51.430 ;
        RECT 297.930 50.410 298.120 51.770 ;
        RECT 298.300 51.405 298.810 51.940 ;
        RECT 299.030 51.130 299.275 51.735 ;
        RECT 299.810 51.390 299.980 51.680 ;
        RECT 300.150 51.560 300.480 51.940 ;
        RECT 299.810 51.220 300.475 51.390 ;
        RECT 298.320 50.960 299.550 51.130 ;
        RECT 297.110 50.240 298.120 50.410 ;
        RECT 298.290 50.395 299.040 50.585 ;
        RECT 296.770 49.900 297.895 50.070 ;
        RECT 298.290 49.730 298.460 50.395 ;
        RECT 299.210 50.150 299.550 50.960 ;
        RECT 299.725 50.400 300.075 51.050 ;
        RECT 300.245 50.230 300.475 51.220 ;
        RECT 296.430 49.560 298.460 49.730 ;
        RECT 298.630 49.390 298.800 50.150 ;
        RECT 299.035 49.740 299.550 50.150 ;
        RECT 299.810 50.060 300.475 50.230 ;
        RECT 299.810 49.560 299.980 50.060 ;
        RECT 300.150 49.390 300.480 49.890 ;
        RECT 300.650 49.560 300.875 51.680 ;
        RECT 301.090 51.560 301.420 51.940 ;
        RECT 301.590 51.390 301.760 51.720 ;
        RECT 302.060 51.560 303.075 51.760 ;
        RECT 301.065 51.200 301.760 51.390 ;
        RECT 301.065 50.230 301.235 51.200 ;
        RECT 301.405 50.400 301.815 51.020 ;
        RECT 301.985 50.450 302.205 51.320 ;
        RECT 302.385 51.010 302.735 51.380 ;
        RECT 302.905 50.830 303.075 51.560 ;
        RECT 303.245 51.500 303.655 51.940 ;
        RECT 303.945 51.300 304.195 51.730 ;
        RECT 304.395 51.480 304.715 51.940 ;
        RECT 305.275 51.550 306.125 51.720 ;
        RECT 303.245 50.960 303.655 51.290 ;
        RECT 303.945 50.960 304.365 51.300 ;
        RECT 302.655 50.790 303.075 50.830 ;
        RECT 302.655 50.620 304.005 50.790 ;
        RECT 301.065 50.060 301.760 50.230 ;
        RECT 301.985 50.070 302.485 50.450 ;
        RECT 301.090 49.390 301.420 49.890 ;
        RECT 301.590 49.560 301.760 50.060 ;
        RECT 302.655 49.775 302.825 50.620 ;
        RECT 303.755 50.460 304.005 50.620 ;
        RECT 302.995 50.190 303.245 50.450 ;
        RECT 304.175 50.190 304.365 50.960 ;
        RECT 302.995 49.940 304.365 50.190 ;
        RECT 304.535 51.130 305.785 51.300 ;
        RECT 304.535 50.370 304.705 51.130 ;
        RECT 305.455 51.010 305.785 51.130 ;
        RECT 304.875 50.550 305.055 50.960 ;
        RECT 305.955 50.790 306.125 51.550 ;
        RECT 306.325 51.460 306.985 51.940 ;
        RECT 307.165 51.345 307.485 51.675 ;
        RECT 306.315 51.020 306.975 51.290 ;
        RECT 306.315 50.960 306.645 51.020 ;
        RECT 306.795 50.790 307.125 50.850 ;
        RECT 305.225 50.620 307.125 50.790 ;
        RECT 304.535 50.060 305.055 50.370 ;
        RECT 305.225 50.110 305.395 50.620 ;
        RECT 307.295 50.450 307.485 51.345 ;
        RECT 305.565 50.280 307.485 50.450 ;
        RECT 307.165 50.260 307.485 50.280 ;
        RECT 307.685 51.030 307.935 51.680 ;
        RECT 308.115 51.480 308.400 51.940 ;
        RECT 308.580 51.600 308.835 51.760 ;
        RECT 308.580 51.430 308.920 51.600 ;
        RECT 308.580 51.230 308.835 51.430 ;
        RECT 307.685 50.700 308.485 51.030 ;
        RECT 305.225 49.940 306.435 50.110 ;
        RECT 301.995 49.605 302.825 49.775 ;
        RECT 303.065 49.390 303.445 49.770 ;
        RECT 303.625 49.650 303.795 49.940 ;
        RECT 305.225 49.860 305.395 49.940 ;
        RECT 303.965 49.390 304.295 49.770 ;
        RECT 304.765 49.610 305.395 49.860 ;
        RECT 305.575 49.390 305.995 49.770 ;
        RECT 306.195 49.650 306.435 49.940 ;
        RECT 306.665 49.390 306.995 50.080 ;
        RECT 307.165 49.650 307.335 50.260 ;
        RECT 307.685 50.110 307.935 50.700 ;
        RECT 308.655 50.370 308.835 51.230 ;
        RECT 309.840 51.190 311.050 51.940 ;
        RECT 307.605 49.600 307.935 50.110 ;
        RECT 308.115 49.390 308.400 50.190 ;
        RECT 308.580 49.700 308.835 50.370 ;
        RECT 309.840 50.480 310.360 51.020 ;
        RECT 310.530 50.650 311.050 51.190 ;
        RECT 309.840 49.390 311.050 50.480 ;
        RECT 162.095 49.220 311.135 49.390 ;
        RECT 162.180 48.130 163.390 49.220 ;
        RECT 163.560 48.785 168.905 49.220 ;
        RECT 169.080 48.785 174.425 49.220 ;
        RECT 162.180 47.420 162.700 47.960 ;
        RECT 162.870 47.590 163.390 48.130 ;
        RECT 162.180 46.670 163.390 47.420 ;
        RECT 165.145 47.215 165.485 48.045 ;
        RECT 166.965 47.535 167.315 48.785 ;
        RECT 170.665 47.215 171.005 48.045 ;
        RECT 172.485 47.535 172.835 48.785 ;
        RECT 175.060 48.055 175.350 49.220 ;
        RECT 175.520 48.130 176.730 49.220 ;
        RECT 175.520 47.420 176.040 47.960 ;
        RECT 176.210 47.590 176.730 48.130 ;
        RECT 176.990 48.290 177.160 49.050 ;
        RECT 177.340 48.460 177.670 49.220 ;
        RECT 176.990 48.120 177.655 48.290 ;
        RECT 177.840 48.145 178.110 49.050 ;
        RECT 177.485 47.975 177.655 48.120 ;
        RECT 176.920 47.570 177.250 47.940 ;
        RECT 177.485 47.645 177.770 47.975 ;
        RECT 163.560 46.670 168.905 47.215 ;
        RECT 169.080 46.670 174.425 47.215 ;
        RECT 175.060 46.670 175.350 47.395 ;
        RECT 175.520 46.670 176.730 47.420 ;
        RECT 177.485 47.390 177.655 47.645 ;
        RECT 176.990 47.220 177.655 47.390 ;
        RECT 177.940 47.345 178.110 48.145 ;
        RECT 178.280 48.130 179.490 49.220 ;
        RECT 179.665 48.550 179.920 49.050 ;
        RECT 180.090 48.720 180.420 49.220 ;
        RECT 179.665 48.380 180.415 48.550 ;
        RECT 176.990 46.840 177.160 47.220 ;
        RECT 177.340 46.670 177.670 47.050 ;
        RECT 177.850 46.840 178.110 47.345 ;
        RECT 178.280 47.420 178.800 47.960 ;
        RECT 178.970 47.590 179.490 48.130 ;
        RECT 179.665 47.560 180.015 48.210 ;
        RECT 178.280 46.670 179.490 47.420 ;
        RECT 180.185 47.390 180.415 48.380 ;
        RECT 179.665 47.220 180.415 47.390 ;
        RECT 179.665 46.930 179.920 47.220 ;
        RECT 180.090 46.670 180.420 47.050 ;
        RECT 180.590 46.930 180.760 49.050 ;
        RECT 180.930 48.250 181.255 49.035 ;
        RECT 181.425 48.760 181.675 49.220 ;
        RECT 181.845 48.720 182.095 49.050 ;
        RECT 182.310 48.720 182.990 49.050 ;
        RECT 181.845 48.590 182.015 48.720 ;
        RECT 181.620 48.420 182.015 48.590 ;
        RECT 180.990 47.200 181.450 48.250 ;
        RECT 181.620 47.060 181.790 48.420 ;
        RECT 182.185 48.160 182.650 48.550 ;
        RECT 181.960 47.350 182.310 47.970 ;
        RECT 182.480 47.570 182.650 48.160 ;
        RECT 182.820 47.940 182.990 48.720 ;
        RECT 183.160 48.620 183.330 48.960 ;
        RECT 183.565 48.790 183.895 49.220 ;
        RECT 184.065 48.620 184.235 48.960 ;
        RECT 184.530 48.760 184.900 49.220 ;
        RECT 183.160 48.450 184.235 48.620 ;
        RECT 185.070 48.590 185.240 49.050 ;
        RECT 185.475 48.710 186.345 49.050 ;
        RECT 186.515 48.760 186.765 49.220 ;
        RECT 184.680 48.420 185.240 48.590 ;
        RECT 184.680 48.280 184.850 48.420 ;
        RECT 183.350 48.110 184.850 48.280 ;
        RECT 185.545 48.250 186.005 48.540 ;
        RECT 182.820 47.770 184.510 47.940 ;
        RECT 182.480 47.350 182.835 47.570 ;
        RECT 183.005 47.060 183.175 47.770 ;
        RECT 183.380 47.350 184.170 47.600 ;
        RECT 184.340 47.590 184.510 47.770 ;
        RECT 184.680 47.420 184.850 48.110 ;
        RECT 181.120 46.670 181.450 47.030 ;
        RECT 181.620 46.890 182.115 47.060 ;
        RECT 182.320 46.890 183.175 47.060 ;
        RECT 184.050 46.670 184.380 47.130 ;
        RECT 184.590 47.030 184.850 47.420 ;
        RECT 185.040 48.240 186.005 48.250 ;
        RECT 186.175 48.330 186.345 48.710 ;
        RECT 186.935 48.670 187.105 48.960 ;
        RECT 187.285 48.840 187.615 49.220 ;
        RECT 186.935 48.500 187.735 48.670 ;
        RECT 185.040 48.080 185.715 48.240 ;
        RECT 186.175 48.160 187.395 48.330 ;
        RECT 185.040 47.290 185.250 48.080 ;
        RECT 186.175 48.070 186.345 48.160 ;
        RECT 185.420 47.290 185.770 47.910 ;
        RECT 185.940 47.900 186.345 48.070 ;
        RECT 185.940 47.120 186.110 47.900 ;
        RECT 186.280 47.450 186.500 47.730 ;
        RECT 186.680 47.620 187.220 47.990 ;
        RECT 187.565 47.880 187.735 48.500 ;
        RECT 187.910 48.160 188.080 49.220 ;
        RECT 188.290 48.210 188.580 49.050 ;
        RECT 188.750 48.380 188.920 49.220 ;
        RECT 189.130 48.210 189.380 49.050 ;
        RECT 189.590 48.380 189.760 49.220 ;
        RECT 190.330 48.290 190.500 49.050 ;
        RECT 190.680 48.460 191.010 49.220 ;
        RECT 188.290 48.040 190.015 48.210 ;
        RECT 190.330 48.120 190.995 48.290 ;
        RECT 191.180 48.145 191.450 49.050 ;
        RECT 191.625 48.550 191.880 49.050 ;
        RECT 192.050 48.720 192.380 49.220 ;
        RECT 191.625 48.380 192.375 48.550 ;
        RECT 186.280 47.280 186.810 47.450 ;
        RECT 184.590 46.860 184.940 47.030 ;
        RECT 185.160 46.840 186.110 47.120 ;
        RECT 186.280 46.670 186.470 47.110 ;
        RECT 186.640 47.050 186.810 47.280 ;
        RECT 186.980 47.220 187.220 47.620 ;
        RECT 187.390 47.870 187.735 47.880 ;
        RECT 187.390 47.660 189.420 47.870 ;
        RECT 187.390 47.405 187.715 47.660 ;
        RECT 189.605 47.490 190.015 48.040 ;
        RECT 190.825 47.975 190.995 48.120 ;
        RECT 190.260 47.570 190.590 47.940 ;
        RECT 190.825 47.645 191.110 47.975 ;
        RECT 187.390 47.050 187.710 47.405 ;
        RECT 186.640 46.880 187.710 47.050 ;
        RECT 187.910 46.670 188.080 47.480 ;
        RECT 188.250 47.320 190.015 47.490 ;
        RECT 190.825 47.390 190.995 47.645 ;
        RECT 188.250 46.840 188.580 47.320 ;
        RECT 188.750 46.670 188.920 47.140 ;
        RECT 189.090 46.840 189.420 47.320 ;
        RECT 190.330 47.220 190.995 47.390 ;
        RECT 191.280 47.345 191.450 48.145 ;
        RECT 191.625 47.560 191.975 48.210 ;
        RECT 192.145 47.390 192.375 48.380 ;
        RECT 189.590 46.670 189.760 47.140 ;
        RECT 190.330 46.840 190.500 47.220 ;
        RECT 190.680 46.670 191.010 47.050 ;
        RECT 191.190 46.840 191.450 47.345 ;
        RECT 191.625 47.220 192.375 47.390 ;
        RECT 191.625 46.930 191.880 47.220 ;
        RECT 192.050 46.670 192.380 47.050 ;
        RECT 192.550 46.930 192.720 49.050 ;
        RECT 192.890 48.250 193.215 49.035 ;
        RECT 193.385 48.760 193.635 49.220 ;
        RECT 193.805 48.720 194.055 49.050 ;
        RECT 194.270 48.720 194.950 49.050 ;
        RECT 193.805 48.590 193.975 48.720 ;
        RECT 193.580 48.420 193.975 48.590 ;
        RECT 192.950 47.200 193.410 48.250 ;
        RECT 193.580 47.060 193.750 48.420 ;
        RECT 194.145 48.160 194.610 48.550 ;
        RECT 193.920 47.350 194.270 47.970 ;
        RECT 194.440 47.570 194.610 48.160 ;
        RECT 194.780 47.940 194.950 48.720 ;
        RECT 195.120 48.620 195.290 48.960 ;
        RECT 195.525 48.790 195.855 49.220 ;
        RECT 196.025 48.620 196.195 48.960 ;
        RECT 196.490 48.760 196.860 49.220 ;
        RECT 195.120 48.450 196.195 48.620 ;
        RECT 197.030 48.590 197.200 49.050 ;
        RECT 197.435 48.710 198.305 49.050 ;
        RECT 198.475 48.760 198.725 49.220 ;
        RECT 196.640 48.420 197.200 48.590 ;
        RECT 196.640 48.280 196.810 48.420 ;
        RECT 195.310 48.110 196.810 48.280 ;
        RECT 197.505 48.250 197.965 48.540 ;
        RECT 194.780 47.770 196.470 47.940 ;
        RECT 194.440 47.350 194.795 47.570 ;
        RECT 194.965 47.060 195.135 47.770 ;
        RECT 195.340 47.350 196.130 47.600 ;
        RECT 196.300 47.590 196.470 47.770 ;
        RECT 196.640 47.420 196.810 48.110 ;
        RECT 193.080 46.670 193.410 47.030 ;
        RECT 193.580 46.890 194.075 47.060 ;
        RECT 194.280 46.890 195.135 47.060 ;
        RECT 196.010 46.670 196.340 47.130 ;
        RECT 196.550 47.030 196.810 47.420 ;
        RECT 197.000 48.240 197.965 48.250 ;
        RECT 198.135 48.330 198.305 48.710 ;
        RECT 198.895 48.670 199.065 48.960 ;
        RECT 199.245 48.840 199.575 49.220 ;
        RECT 198.895 48.500 199.695 48.670 ;
        RECT 197.000 48.080 197.675 48.240 ;
        RECT 198.135 48.160 199.355 48.330 ;
        RECT 197.000 47.290 197.210 48.080 ;
        RECT 198.135 48.070 198.305 48.160 ;
        RECT 197.380 47.290 197.730 47.910 ;
        RECT 197.900 47.900 198.305 48.070 ;
        RECT 197.900 47.120 198.070 47.900 ;
        RECT 198.240 47.450 198.460 47.730 ;
        RECT 198.640 47.620 199.180 47.990 ;
        RECT 199.525 47.910 199.695 48.500 ;
        RECT 199.915 48.080 200.220 49.220 ;
        RECT 200.390 48.030 200.645 48.910 ;
        RECT 200.820 48.055 201.110 49.220 ;
        RECT 201.335 48.350 201.620 49.220 ;
        RECT 201.790 48.590 202.050 49.050 ;
        RECT 202.225 48.760 202.480 49.220 ;
        RECT 202.650 48.590 202.910 49.050 ;
        RECT 201.790 48.420 202.910 48.590 ;
        RECT 203.080 48.420 203.390 49.220 ;
        RECT 201.790 48.170 202.050 48.420 ;
        RECT 203.560 48.250 203.870 49.050 ;
        RECT 199.525 47.880 200.265 47.910 ;
        RECT 198.240 47.280 198.770 47.450 ;
        RECT 196.550 46.860 196.900 47.030 ;
        RECT 197.120 46.840 198.070 47.120 ;
        RECT 198.240 46.670 198.430 47.110 ;
        RECT 198.600 47.050 198.770 47.280 ;
        RECT 198.940 47.220 199.180 47.620 ;
        RECT 199.350 47.580 200.265 47.880 ;
        RECT 199.350 47.405 199.675 47.580 ;
        RECT 199.350 47.050 199.670 47.405 ;
        RECT 200.435 47.380 200.645 48.030 ;
        RECT 201.295 48.000 202.050 48.170 ;
        RECT 202.840 48.080 203.870 48.250 ;
        RECT 204.510 48.080 204.840 49.220 ;
        RECT 205.370 48.250 205.700 49.035 ;
        RECT 205.020 48.080 205.700 48.250 ;
        RECT 205.880 48.130 208.470 49.220 ;
        RECT 208.890 48.490 209.185 49.220 ;
        RECT 209.355 48.320 209.615 49.045 ;
        RECT 209.785 48.490 210.045 49.220 ;
        RECT 210.215 48.320 210.475 49.045 ;
        RECT 210.645 48.490 210.905 49.220 ;
        RECT 211.075 48.320 211.335 49.045 ;
        RECT 211.505 48.490 211.765 49.220 ;
        RECT 211.935 48.320 212.195 49.045 ;
        RECT 201.295 47.490 201.700 48.000 ;
        RECT 202.840 47.830 203.010 48.080 ;
        RECT 201.870 47.660 203.010 47.830 ;
        RECT 198.600 46.880 199.670 47.050 ;
        RECT 199.915 46.670 200.220 47.130 ;
        RECT 200.390 46.850 200.645 47.380 ;
        RECT 200.820 46.670 201.110 47.395 ;
        RECT 201.295 47.320 202.945 47.490 ;
        RECT 203.180 47.340 203.530 47.910 ;
        RECT 201.340 46.670 201.620 47.150 ;
        RECT 201.790 46.930 202.050 47.320 ;
        RECT 202.225 46.670 202.480 47.150 ;
        RECT 202.650 46.930 202.945 47.320 ;
        RECT 203.700 47.170 203.870 48.080 ;
        RECT 204.500 47.660 204.850 47.910 ;
        RECT 205.020 47.480 205.190 48.080 ;
        RECT 205.360 47.660 205.710 47.910 ;
        RECT 203.125 46.670 203.400 47.150 ;
        RECT 203.570 46.840 203.870 47.170 ;
        RECT 204.510 46.670 204.780 47.480 ;
        RECT 204.950 46.840 205.280 47.480 ;
        RECT 205.450 46.670 205.690 47.480 ;
        RECT 205.880 47.440 207.090 47.960 ;
        RECT 207.260 47.610 208.470 48.130 ;
        RECT 208.885 48.080 212.195 48.320 ;
        RECT 212.365 48.110 212.625 49.220 ;
        RECT 208.885 47.490 209.855 48.080 ;
        RECT 212.795 47.910 213.045 49.045 ;
        RECT 213.225 48.110 213.520 49.220 ;
        RECT 213.700 48.710 213.960 49.220 ;
        RECT 210.025 47.660 213.045 47.910 ;
        RECT 205.880 46.670 208.470 47.440 ;
        RECT 208.885 47.320 212.195 47.490 ;
        RECT 208.885 46.670 209.185 47.150 ;
        RECT 209.355 46.865 209.615 47.320 ;
        RECT 209.785 46.670 210.045 47.150 ;
        RECT 210.215 46.865 210.475 47.320 ;
        RECT 210.645 46.670 210.905 47.150 ;
        RECT 211.075 46.865 211.335 47.320 ;
        RECT 211.505 46.670 211.765 47.150 ;
        RECT 211.935 46.865 212.195 47.320 ;
        RECT 212.365 46.670 212.625 47.195 ;
        RECT 212.795 46.850 213.045 47.660 ;
        RECT 213.215 47.300 213.530 47.910 ;
        RECT 213.700 47.660 214.040 48.540 ;
        RECT 214.210 47.830 214.380 49.050 ;
        RECT 214.620 48.715 215.235 49.220 ;
        RECT 214.620 48.180 214.870 48.545 ;
        RECT 215.040 48.540 215.235 48.715 ;
        RECT 215.405 48.710 215.880 49.050 ;
        RECT 216.050 48.675 216.265 49.220 ;
        RECT 215.040 48.350 215.370 48.540 ;
        RECT 215.590 48.180 216.305 48.475 ;
        RECT 216.475 48.350 216.750 49.050 ;
        RECT 218.040 48.550 218.320 49.220 ;
        RECT 214.620 48.010 216.410 48.180 ;
        RECT 214.210 47.580 215.005 47.830 ;
        RECT 214.210 47.490 214.460 47.580 ;
        RECT 213.225 46.670 213.470 47.130 ;
        RECT 213.700 46.670 213.960 47.490 ;
        RECT 214.130 47.070 214.460 47.490 ;
        RECT 215.175 47.155 215.430 48.010 ;
        RECT 214.640 46.890 215.430 47.155 ;
        RECT 215.600 47.310 216.010 47.830 ;
        RECT 216.180 47.580 216.410 48.010 ;
        RECT 216.580 47.320 216.750 48.350 ;
        RECT 218.490 48.330 218.790 48.880 ;
        RECT 218.990 48.500 219.320 49.220 ;
        RECT 219.510 48.500 219.970 49.050 ;
        RECT 217.855 47.910 218.120 48.270 ;
        RECT 218.490 48.160 219.430 48.330 ;
        RECT 219.260 47.910 219.430 48.160 ;
        RECT 217.855 47.660 218.530 47.910 ;
        RECT 218.750 47.660 219.090 47.910 ;
        RECT 219.260 47.580 219.550 47.910 ;
        RECT 219.260 47.490 219.430 47.580 ;
        RECT 215.600 46.890 215.800 47.310 ;
        RECT 215.990 46.670 216.320 47.130 ;
        RECT 216.490 46.840 216.750 47.320 ;
        RECT 218.040 47.300 219.430 47.490 ;
        RECT 218.040 46.940 218.370 47.300 ;
        RECT 219.720 47.130 219.970 48.500 ;
        RECT 220.140 48.130 221.810 49.220 ;
        RECT 218.990 46.670 219.240 47.130 ;
        RECT 219.410 46.840 219.970 47.130 ;
        RECT 220.140 47.440 220.890 47.960 ;
        RECT 221.060 47.610 221.810 48.130 ;
        RECT 222.530 48.290 222.700 49.050 ;
        RECT 222.915 48.460 223.245 49.220 ;
        RECT 222.530 48.120 223.245 48.290 ;
        RECT 223.415 48.145 223.670 49.050 ;
        RECT 222.440 47.570 222.795 47.940 ;
        RECT 223.075 47.910 223.245 48.120 ;
        RECT 223.075 47.580 223.330 47.910 ;
        RECT 220.140 46.670 221.810 47.440 ;
        RECT 223.075 47.390 223.245 47.580 ;
        RECT 223.500 47.415 223.670 48.145 ;
        RECT 223.845 48.070 224.105 49.220 ;
        RECT 224.740 48.145 225.010 49.050 ;
        RECT 225.180 48.460 225.510 49.220 ;
        RECT 225.690 48.290 225.860 49.050 ;
        RECT 222.530 47.220 223.245 47.390 ;
        RECT 222.530 46.840 222.700 47.220 ;
        RECT 222.915 46.670 223.245 47.050 ;
        RECT 223.415 46.840 223.670 47.415 ;
        RECT 223.845 46.670 224.105 47.510 ;
        RECT 224.740 47.345 224.910 48.145 ;
        RECT 225.195 48.120 225.860 48.290 ;
        RECT 225.195 47.975 225.365 48.120 ;
        RECT 226.580 48.055 226.870 49.220 ;
        RECT 227.130 48.290 227.300 49.050 ;
        RECT 227.515 48.460 227.845 49.220 ;
        RECT 227.130 48.120 227.845 48.290 ;
        RECT 228.015 48.145 228.270 49.050 ;
        RECT 225.080 47.645 225.365 47.975 ;
        RECT 225.195 47.390 225.365 47.645 ;
        RECT 225.600 47.570 225.930 47.940 ;
        RECT 227.040 47.570 227.395 47.940 ;
        RECT 227.675 47.910 227.845 48.120 ;
        RECT 227.675 47.580 227.930 47.910 ;
        RECT 224.740 46.840 225.000 47.345 ;
        RECT 225.195 47.220 225.860 47.390 ;
        RECT 225.180 46.670 225.510 47.050 ;
        RECT 225.690 46.840 225.860 47.220 ;
        RECT 226.580 46.670 226.870 47.395 ;
        RECT 227.675 47.390 227.845 47.580 ;
        RECT 228.100 47.415 228.270 48.145 ;
        RECT 228.445 48.070 228.705 49.220 ;
        RECT 229.805 48.550 230.060 49.050 ;
        RECT 230.230 48.720 230.560 49.220 ;
        RECT 229.805 48.380 230.555 48.550 ;
        RECT 229.805 47.560 230.155 48.210 ;
        RECT 227.130 47.220 227.845 47.390 ;
        RECT 227.130 46.840 227.300 47.220 ;
        RECT 227.515 46.670 227.845 47.050 ;
        RECT 228.015 46.840 228.270 47.415 ;
        RECT 228.445 46.670 228.705 47.510 ;
        RECT 230.325 47.390 230.555 48.380 ;
        RECT 229.805 47.220 230.555 47.390 ;
        RECT 229.805 46.930 230.060 47.220 ;
        RECT 230.230 46.670 230.560 47.050 ;
        RECT 230.730 46.930 230.900 49.050 ;
        RECT 231.070 48.250 231.395 49.035 ;
        RECT 231.565 48.760 231.815 49.220 ;
        RECT 231.985 48.720 232.235 49.050 ;
        RECT 232.450 48.720 233.130 49.050 ;
        RECT 231.985 48.590 232.155 48.720 ;
        RECT 231.760 48.420 232.155 48.590 ;
        RECT 231.130 47.200 231.590 48.250 ;
        RECT 231.760 47.060 231.930 48.420 ;
        RECT 232.325 48.160 232.790 48.550 ;
        RECT 232.100 47.350 232.450 47.970 ;
        RECT 232.620 47.570 232.790 48.160 ;
        RECT 232.960 47.940 233.130 48.720 ;
        RECT 233.300 48.620 233.470 48.960 ;
        RECT 233.705 48.790 234.035 49.220 ;
        RECT 234.205 48.620 234.375 48.960 ;
        RECT 234.670 48.760 235.040 49.220 ;
        RECT 233.300 48.450 234.375 48.620 ;
        RECT 235.210 48.590 235.380 49.050 ;
        RECT 235.615 48.710 236.485 49.050 ;
        RECT 236.655 48.760 236.905 49.220 ;
        RECT 234.820 48.420 235.380 48.590 ;
        RECT 234.820 48.280 234.990 48.420 ;
        RECT 233.490 48.110 234.990 48.280 ;
        RECT 235.685 48.250 236.145 48.540 ;
        RECT 232.960 47.770 234.650 47.940 ;
        RECT 232.620 47.350 232.975 47.570 ;
        RECT 233.145 47.060 233.315 47.770 ;
        RECT 233.520 47.350 234.310 47.600 ;
        RECT 234.480 47.590 234.650 47.770 ;
        RECT 234.820 47.420 234.990 48.110 ;
        RECT 231.260 46.670 231.590 47.030 ;
        RECT 231.760 46.890 232.255 47.060 ;
        RECT 232.460 46.890 233.315 47.060 ;
        RECT 234.190 46.670 234.520 47.130 ;
        RECT 234.730 47.030 234.990 47.420 ;
        RECT 235.180 48.240 236.145 48.250 ;
        RECT 236.315 48.330 236.485 48.710 ;
        RECT 237.075 48.670 237.245 48.960 ;
        RECT 237.425 48.840 237.755 49.220 ;
        RECT 237.075 48.500 237.875 48.670 ;
        RECT 235.180 48.080 235.855 48.240 ;
        RECT 236.315 48.160 237.535 48.330 ;
        RECT 235.180 47.290 235.390 48.080 ;
        RECT 236.315 48.070 236.485 48.160 ;
        RECT 235.560 47.290 235.910 47.910 ;
        RECT 236.080 47.900 236.485 48.070 ;
        RECT 236.080 47.120 236.250 47.900 ;
        RECT 236.420 47.450 236.640 47.730 ;
        RECT 236.820 47.620 237.360 47.990 ;
        RECT 237.705 47.910 237.875 48.500 ;
        RECT 238.095 48.080 238.400 49.220 ;
        RECT 238.570 48.030 238.825 48.910 ;
        RECT 239.005 48.550 239.260 49.050 ;
        RECT 239.430 48.720 239.760 49.220 ;
        RECT 239.005 48.380 239.755 48.550 ;
        RECT 237.705 47.880 238.445 47.910 ;
        RECT 236.420 47.280 236.950 47.450 ;
        RECT 234.730 46.860 235.080 47.030 ;
        RECT 235.300 46.840 236.250 47.120 ;
        RECT 236.420 46.670 236.610 47.110 ;
        RECT 236.780 47.050 236.950 47.280 ;
        RECT 237.120 47.220 237.360 47.620 ;
        RECT 237.530 47.580 238.445 47.880 ;
        RECT 237.530 47.405 237.855 47.580 ;
        RECT 237.530 47.050 237.850 47.405 ;
        RECT 238.615 47.380 238.825 48.030 ;
        RECT 239.005 47.560 239.355 48.210 ;
        RECT 239.525 47.390 239.755 48.380 ;
        RECT 236.780 46.880 237.850 47.050 ;
        RECT 238.095 46.670 238.400 47.130 ;
        RECT 238.570 46.850 238.825 47.380 ;
        RECT 239.005 47.220 239.755 47.390 ;
        RECT 239.005 46.930 239.260 47.220 ;
        RECT 239.430 46.670 239.760 47.050 ;
        RECT 239.930 46.930 240.100 49.050 ;
        RECT 240.270 48.250 240.595 49.035 ;
        RECT 240.765 48.760 241.015 49.220 ;
        RECT 241.185 48.720 241.435 49.050 ;
        RECT 241.650 48.720 242.330 49.050 ;
        RECT 241.185 48.590 241.355 48.720 ;
        RECT 240.960 48.420 241.355 48.590 ;
        RECT 240.330 47.200 240.790 48.250 ;
        RECT 240.960 47.060 241.130 48.420 ;
        RECT 241.525 48.160 241.990 48.550 ;
        RECT 241.300 47.350 241.650 47.970 ;
        RECT 241.820 47.570 241.990 48.160 ;
        RECT 242.160 47.940 242.330 48.720 ;
        RECT 242.500 48.620 242.670 48.960 ;
        RECT 242.905 48.790 243.235 49.220 ;
        RECT 243.405 48.620 243.575 48.960 ;
        RECT 243.870 48.760 244.240 49.220 ;
        RECT 242.500 48.450 243.575 48.620 ;
        RECT 244.410 48.590 244.580 49.050 ;
        RECT 244.815 48.710 245.685 49.050 ;
        RECT 245.855 48.760 246.105 49.220 ;
        RECT 244.020 48.420 244.580 48.590 ;
        RECT 244.020 48.280 244.190 48.420 ;
        RECT 242.690 48.110 244.190 48.280 ;
        RECT 244.885 48.250 245.345 48.540 ;
        RECT 242.160 47.770 243.850 47.940 ;
        RECT 241.820 47.350 242.175 47.570 ;
        RECT 242.345 47.060 242.515 47.770 ;
        RECT 242.720 47.350 243.510 47.600 ;
        RECT 243.680 47.590 243.850 47.770 ;
        RECT 244.020 47.420 244.190 48.110 ;
        RECT 240.460 46.670 240.790 47.030 ;
        RECT 240.960 46.890 241.455 47.060 ;
        RECT 241.660 46.890 242.515 47.060 ;
        RECT 243.390 46.670 243.720 47.130 ;
        RECT 243.930 47.030 244.190 47.420 ;
        RECT 244.380 48.240 245.345 48.250 ;
        RECT 245.515 48.330 245.685 48.710 ;
        RECT 246.275 48.670 246.445 48.960 ;
        RECT 246.625 48.840 246.955 49.220 ;
        RECT 246.275 48.500 247.075 48.670 ;
        RECT 244.380 48.080 245.055 48.240 ;
        RECT 245.515 48.160 246.735 48.330 ;
        RECT 244.380 47.290 244.590 48.080 ;
        RECT 245.515 48.070 245.685 48.160 ;
        RECT 244.760 47.290 245.110 47.910 ;
        RECT 245.280 47.900 245.685 48.070 ;
        RECT 245.280 47.120 245.450 47.900 ;
        RECT 245.620 47.450 245.840 47.730 ;
        RECT 246.020 47.620 246.560 47.990 ;
        RECT 246.905 47.910 247.075 48.500 ;
        RECT 247.295 48.080 247.600 49.220 ;
        RECT 247.770 48.030 248.025 48.910 ;
        RECT 248.200 48.130 251.710 49.220 ;
        RECT 246.905 47.880 247.645 47.910 ;
        RECT 245.620 47.280 246.150 47.450 ;
        RECT 243.930 46.860 244.280 47.030 ;
        RECT 244.500 46.840 245.450 47.120 ;
        RECT 245.620 46.670 245.810 47.110 ;
        RECT 245.980 47.050 246.150 47.280 ;
        RECT 246.320 47.220 246.560 47.620 ;
        RECT 246.730 47.580 247.645 47.880 ;
        RECT 246.730 47.405 247.055 47.580 ;
        RECT 246.730 47.050 247.050 47.405 ;
        RECT 247.815 47.380 248.025 48.030 ;
        RECT 245.980 46.880 247.050 47.050 ;
        RECT 247.295 46.670 247.600 47.130 ;
        RECT 247.770 46.850 248.025 47.380 ;
        RECT 248.200 47.440 249.850 47.960 ;
        RECT 250.020 47.610 251.710 48.130 ;
        RECT 252.340 48.055 252.630 49.220 ;
        RECT 252.800 48.130 255.390 49.220 ;
        RECT 255.565 48.550 255.820 49.050 ;
        RECT 255.990 48.720 256.320 49.220 ;
        RECT 255.565 48.380 256.315 48.550 ;
        RECT 252.800 47.440 254.010 47.960 ;
        RECT 254.180 47.610 255.390 48.130 ;
        RECT 255.565 47.560 255.915 48.210 ;
        RECT 248.200 46.670 251.710 47.440 ;
        RECT 252.340 46.670 252.630 47.395 ;
        RECT 252.800 46.670 255.390 47.440 ;
        RECT 256.085 47.390 256.315 48.380 ;
        RECT 255.565 47.220 256.315 47.390 ;
        RECT 255.565 46.930 255.820 47.220 ;
        RECT 255.990 46.670 256.320 47.050 ;
        RECT 256.490 46.930 256.660 49.050 ;
        RECT 256.830 48.250 257.155 49.035 ;
        RECT 257.325 48.760 257.575 49.220 ;
        RECT 257.745 48.720 257.995 49.050 ;
        RECT 258.210 48.720 258.890 49.050 ;
        RECT 257.745 48.590 257.915 48.720 ;
        RECT 257.520 48.420 257.915 48.590 ;
        RECT 256.890 47.200 257.350 48.250 ;
        RECT 257.520 47.060 257.690 48.420 ;
        RECT 258.085 48.160 258.550 48.550 ;
        RECT 257.860 47.350 258.210 47.970 ;
        RECT 258.380 47.570 258.550 48.160 ;
        RECT 258.720 47.940 258.890 48.720 ;
        RECT 259.060 48.620 259.230 48.960 ;
        RECT 259.465 48.790 259.795 49.220 ;
        RECT 259.965 48.620 260.135 48.960 ;
        RECT 260.430 48.760 260.800 49.220 ;
        RECT 259.060 48.450 260.135 48.620 ;
        RECT 260.970 48.590 261.140 49.050 ;
        RECT 261.375 48.710 262.245 49.050 ;
        RECT 262.415 48.760 262.665 49.220 ;
        RECT 260.580 48.420 261.140 48.590 ;
        RECT 260.580 48.280 260.750 48.420 ;
        RECT 259.250 48.110 260.750 48.280 ;
        RECT 261.445 48.250 261.905 48.540 ;
        RECT 258.720 47.770 260.410 47.940 ;
        RECT 258.380 47.350 258.735 47.570 ;
        RECT 258.905 47.060 259.075 47.770 ;
        RECT 259.280 47.350 260.070 47.600 ;
        RECT 260.240 47.590 260.410 47.770 ;
        RECT 260.580 47.420 260.750 48.110 ;
        RECT 257.020 46.670 257.350 47.030 ;
        RECT 257.520 46.890 258.015 47.060 ;
        RECT 258.220 46.890 259.075 47.060 ;
        RECT 259.950 46.670 260.280 47.130 ;
        RECT 260.490 47.030 260.750 47.420 ;
        RECT 260.940 48.240 261.905 48.250 ;
        RECT 262.075 48.330 262.245 48.710 ;
        RECT 262.835 48.670 263.005 48.960 ;
        RECT 263.185 48.840 263.515 49.220 ;
        RECT 262.835 48.500 263.635 48.670 ;
        RECT 260.940 48.080 261.615 48.240 ;
        RECT 262.075 48.160 263.295 48.330 ;
        RECT 260.940 47.290 261.150 48.080 ;
        RECT 262.075 48.070 262.245 48.160 ;
        RECT 261.320 47.290 261.670 47.910 ;
        RECT 261.840 47.900 262.245 48.070 ;
        RECT 261.840 47.120 262.010 47.900 ;
        RECT 262.180 47.450 262.400 47.730 ;
        RECT 262.580 47.620 263.120 47.990 ;
        RECT 263.465 47.910 263.635 48.500 ;
        RECT 263.855 48.080 264.160 49.220 ;
        RECT 264.330 48.030 264.585 48.910 ;
        RECT 264.875 48.590 265.160 49.050 ;
        RECT 265.330 48.760 265.600 49.220 ;
        RECT 264.875 48.370 265.830 48.590 ;
        RECT 263.465 47.880 264.205 47.910 ;
        RECT 262.180 47.280 262.710 47.450 ;
        RECT 260.490 46.860 260.840 47.030 ;
        RECT 261.060 46.840 262.010 47.120 ;
        RECT 262.180 46.670 262.370 47.110 ;
        RECT 262.540 47.050 262.710 47.280 ;
        RECT 262.880 47.220 263.120 47.620 ;
        RECT 263.290 47.580 264.205 47.880 ;
        RECT 263.290 47.405 263.615 47.580 ;
        RECT 263.290 47.050 263.610 47.405 ;
        RECT 264.375 47.380 264.585 48.030 ;
        RECT 264.760 47.640 265.450 48.200 ;
        RECT 265.620 47.470 265.830 48.370 ;
        RECT 262.540 46.880 263.610 47.050 ;
        RECT 263.855 46.670 264.160 47.130 ;
        RECT 264.330 46.850 264.585 47.380 ;
        RECT 264.875 47.300 265.830 47.470 ;
        RECT 266.000 48.200 266.400 49.050 ;
        RECT 266.590 48.590 266.870 49.050 ;
        RECT 267.390 48.760 267.715 49.220 ;
        RECT 266.590 48.370 267.715 48.590 ;
        RECT 266.000 47.640 267.095 48.200 ;
        RECT 267.265 47.910 267.715 48.370 ;
        RECT 267.885 48.080 268.270 49.050 ;
        RECT 264.875 46.840 265.160 47.300 ;
        RECT 265.330 46.670 265.600 47.130 ;
        RECT 266.000 46.840 266.400 47.640 ;
        RECT 267.265 47.580 267.820 47.910 ;
        RECT 267.265 47.470 267.715 47.580 ;
        RECT 266.590 47.300 267.715 47.470 ;
        RECT 267.990 47.410 268.270 48.080 ;
        RECT 266.590 46.840 266.870 47.300 ;
        RECT 267.390 46.670 267.715 47.130 ;
        RECT 267.885 46.840 268.270 47.410 ;
        RECT 268.460 48.380 268.715 49.050 ;
        RECT 268.885 48.460 269.215 49.220 ;
        RECT 269.385 48.620 269.635 49.050 ;
        RECT 269.805 48.800 270.160 49.220 ;
        RECT 270.350 48.880 271.520 49.050 ;
        RECT 270.350 48.840 270.680 48.880 ;
        RECT 270.790 48.620 271.020 48.710 ;
        RECT 269.385 48.380 271.020 48.620 ;
        RECT 271.190 48.380 271.520 48.880 ;
        RECT 268.460 47.250 268.630 48.380 ;
        RECT 271.690 48.210 271.860 49.050 ;
        RECT 268.800 48.040 271.860 48.210 ;
        RECT 272.140 48.380 272.395 49.050 ;
        RECT 272.565 48.460 272.895 49.220 ;
        RECT 273.065 48.620 273.315 49.050 ;
        RECT 273.485 48.800 273.840 49.220 ;
        RECT 274.030 48.880 275.200 49.050 ;
        RECT 274.030 48.840 274.360 48.880 ;
        RECT 274.470 48.620 274.700 48.710 ;
        RECT 273.065 48.380 274.700 48.620 ;
        RECT 274.870 48.380 275.200 48.880 ;
        RECT 268.800 47.490 268.970 48.040 ;
        RECT 269.200 47.660 269.565 47.860 ;
        RECT 269.735 47.660 270.065 47.860 ;
        RECT 268.800 47.320 269.600 47.490 ;
        RECT 268.460 47.180 268.645 47.250 ;
        RECT 268.460 47.170 268.670 47.180 ;
        RECT 268.460 46.840 268.715 47.170 ;
        RECT 268.930 46.670 269.260 47.150 ;
        RECT 269.430 47.090 269.600 47.320 ;
        RECT 269.780 47.260 270.065 47.660 ;
        RECT 270.335 47.660 270.810 47.860 ;
        RECT 270.980 47.660 271.425 47.860 ;
        RECT 271.595 47.660 271.945 47.870 ;
        RECT 270.335 47.260 270.615 47.660 ;
        RECT 270.795 47.320 271.860 47.490 ;
        RECT 270.795 47.090 270.965 47.320 ;
        RECT 269.430 46.840 270.965 47.090 ;
        RECT 271.190 46.670 271.520 47.150 ;
        RECT 271.690 46.840 271.860 47.320 ;
        RECT 272.140 47.250 272.310 48.380 ;
        RECT 275.370 48.210 275.540 49.050 ;
        RECT 272.480 48.040 275.540 48.210 ;
        RECT 275.800 48.500 276.260 49.050 ;
        RECT 276.450 48.500 276.780 49.220 ;
        RECT 272.480 47.490 272.650 48.040 ;
        RECT 272.870 47.690 273.245 47.860 ;
        RECT 272.880 47.660 273.245 47.690 ;
        RECT 273.415 47.660 273.745 47.860 ;
        RECT 272.480 47.320 273.280 47.490 ;
        RECT 272.140 47.170 272.325 47.250 ;
        RECT 272.140 46.840 272.395 47.170 ;
        RECT 272.610 46.670 272.940 47.150 ;
        RECT 273.110 47.090 273.280 47.320 ;
        RECT 273.460 47.260 273.745 47.660 ;
        RECT 274.015 47.660 274.490 47.860 ;
        RECT 274.660 47.660 275.105 47.860 ;
        RECT 275.275 47.660 275.625 47.870 ;
        RECT 274.015 47.260 274.295 47.660 ;
        RECT 274.475 47.320 275.540 47.490 ;
        RECT 274.475 47.090 274.645 47.320 ;
        RECT 273.110 46.840 274.645 47.090 ;
        RECT 274.870 46.670 275.200 47.150 ;
        RECT 275.370 46.840 275.540 47.320 ;
        RECT 275.800 47.130 276.050 48.500 ;
        RECT 276.980 48.330 277.280 48.880 ;
        RECT 277.450 48.550 277.730 49.220 ;
        RECT 276.340 48.160 277.280 48.330 ;
        RECT 276.340 47.910 276.510 48.160 ;
        RECT 277.650 47.910 277.915 48.270 ;
        RECT 278.100 48.055 278.390 49.220 ;
        RECT 278.560 48.080 278.945 49.050 ;
        RECT 279.115 48.760 279.440 49.220 ;
        RECT 279.960 48.590 280.240 49.050 ;
        RECT 279.115 48.370 280.240 48.590 ;
        RECT 276.220 47.580 276.510 47.910 ;
        RECT 276.680 47.660 277.020 47.910 ;
        RECT 277.240 47.660 277.915 47.910 ;
        RECT 276.340 47.490 276.510 47.580 ;
        RECT 276.340 47.300 277.730 47.490 ;
        RECT 278.560 47.410 278.840 48.080 ;
        RECT 279.115 47.910 279.565 48.370 ;
        RECT 280.430 48.200 280.830 49.050 ;
        RECT 281.230 48.760 281.500 49.220 ;
        RECT 281.670 48.590 281.955 49.050 ;
        RECT 279.010 47.580 279.565 47.910 ;
        RECT 279.735 47.640 280.830 48.200 ;
        RECT 279.115 47.470 279.565 47.580 ;
        RECT 275.800 46.840 276.360 47.130 ;
        RECT 276.530 46.670 276.780 47.130 ;
        RECT 277.400 46.940 277.730 47.300 ;
        RECT 278.100 46.670 278.390 47.395 ;
        RECT 278.560 46.840 278.945 47.410 ;
        RECT 279.115 47.300 280.240 47.470 ;
        RECT 279.115 46.670 279.440 47.130 ;
        RECT 279.960 46.840 280.240 47.300 ;
        RECT 280.430 46.840 280.830 47.640 ;
        RECT 281.000 48.370 281.955 48.590 ;
        RECT 282.240 48.500 282.700 49.050 ;
        RECT 282.890 48.500 283.220 49.220 ;
        RECT 281.000 47.470 281.210 48.370 ;
        RECT 281.380 47.640 282.070 48.200 ;
        RECT 281.000 47.300 281.955 47.470 ;
        RECT 281.230 46.670 281.500 47.130 ;
        RECT 281.670 46.840 281.955 47.300 ;
        RECT 282.240 47.130 282.490 48.500 ;
        RECT 283.420 48.330 283.720 48.880 ;
        RECT 283.890 48.550 284.170 49.220 ;
        RECT 282.780 48.160 283.720 48.330 ;
        RECT 282.780 47.910 282.950 48.160 ;
        RECT 284.090 47.910 284.355 48.270 ;
        RECT 282.660 47.580 282.950 47.910 ;
        RECT 283.120 47.660 283.460 47.910 ;
        RECT 283.680 47.660 284.355 47.910 ;
        RECT 285.465 48.030 285.720 48.910 ;
        RECT 285.890 48.080 286.195 49.220 ;
        RECT 286.535 48.840 286.865 49.220 ;
        RECT 287.045 48.670 287.215 48.960 ;
        RECT 287.385 48.760 287.635 49.220 ;
        RECT 286.415 48.500 287.215 48.670 ;
        RECT 287.805 48.710 288.675 49.050 ;
        RECT 282.780 47.490 282.950 47.580 ;
        RECT 282.780 47.300 284.170 47.490 ;
        RECT 282.240 46.840 282.800 47.130 ;
        RECT 282.970 46.670 283.220 47.130 ;
        RECT 283.840 46.940 284.170 47.300 ;
        RECT 285.465 47.380 285.675 48.030 ;
        RECT 286.415 47.910 286.585 48.500 ;
        RECT 287.805 48.330 287.975 48.710 ;
        RECT 288.910 48.590 289.080 49.050 ;
        RECT 289.250 48.760 289.620 49.220 ;
        RECT 289.915 48.620 290.085 48.960 ;
        RECT 290.255 48.790 290.585 49.220 ;
        RECT 290.820 48.620 290.990 48.960 ;
        RECT 286.755 48.160 287.975 48.330 ;
        RECT 288.145 48.250 288.605 48.540 ;
        RECT 288.910 48.420 289.470 48.590 ;
        RECT 289.915 48.450 290.990 48.620 ;
        RECT 291.160 48.720 291.840 49.050 ;
        RECT 292.055 48.720 292.305 49.050 ;
        RECT 292.475 48.760 292.725 49.220 ;
        RECT 289.300 48.280 289.470 48.420 ;
        RECT 288.145 48.240 289.110 48.250 ;
        RECT 287.805 48.070 287.975 48.160 ;
        RECT 288.435 48.080 289.110 48.240 ;
        RECT 285.845 47.880 286.585 47.910 ;
        RECT 285.845 47.580 286.760 47.880 ;
        RECT 286.435 47.405 286.760 47.580 ;
        RECT 285.465 46.850 285.720 47.380 ;
        RECT 285.890 46.670 286.195 47.130 ;
        RECT 286.440 47.050 286.760 47.405 ;
        RECT 286.930 47.620 287.470 47.990 ;
        RECT 287.805 47.900 288.210 48.070 ;
        RECT 286.930 47.220 287.170 47.620 ;
        RECT 287.650 47.450 287.870 47.730 ;
        RECT 287.340 47.280 287.870 47.450 ;
        RECT 287.340 47.050 287.510 47.280 ;
        RECT 288.040 47.120 288.210 47.900 ;
        RECT 288.380 47.290 288.730 47.910 ;
        RECT 288.900 47.290 289.110 48.080 ;
        RECT 289.300 48.110 290.800 48.280 ;
        RECT 289.300 47.420 289.470 48.110 ;
        RECT 291.160 47.940 291.330 48.720 ;
        RECT 292.135 48.590 292.305 48.720 ;
        RECT 289.640 47.770 291.330 47.940 ;
        RECT 291.500 48.160 291.965 48.550 ;
        RECT 292.135 48.420 292.530 48.590 ;
        RECT 289.640 47.590 289.810 47.770 ;
        RECT 286.440 46.880 287.510 47.050 ;
        RECT 287.680 46.670 287.870 47.110 ;
        RECT 288.040 46.840 288.990 47.120 ;
        RECT 289.300 47.030 289.560 47.420 ;
        RECT 289.980 47.350 290.770 47.600 ;
        RECT 289.210 46.860 289.560 47.030 ;
        RECT 289.770 46.670 290.100 47.130 ;
        RECT 290.975 47.060 291.145 47.770 ;
        RECT 291.500 47.570 291.670 48.160 ;
        RECT 291.315 47.350 291.670 47.570 ;
        RECT 291.840 47.350 292.190 47.970 ;
        RECT 292.360 47.060 292.530 48.420 ;
        RECT 292.895 48.250 293.220 49.035 ;
        RECT 292.700 47.200 293.160 48.250 ;
        RECT 290.975 46.890 291.830 47.060 ;
        RECT 292.035 46.890 292.530 47.060 ;
        RECT 292.700 46.670 293.030 47.030 ;
        RECT 293.390 46.930 293.560 49.050 ;
        RECT 293.730 48.720 294.060 49.220 ;
        RECT 294.230 48.550 294.485 49.050 ;
        RECT 293.735 48.380 294.485 48.550 ;
        RECT 294.665 48.550 294.920 49.050 ;
        RECT 295.090 48.720 295.420 49.220 ;
        RECT 294.665 48.380 295.415 48.550 ;
        RECT 293.735 47.390 293.965 48.380 ;
        RECT 294.135 47.560 294.485 48.210 ;
        RECT 294.665 47.560 295.015 48.210 ;
        RECT 295.185 47.390 295.415 48.380 ;
        RECT 293.735 47.220 294.485 47.390 ;
        RECT 293.730 46.670 294.060 47.050 ;
        RECT 294.230 46.930 294.485 47.220 ;
        RECT 294.665 47.220 295.415 47.390 ;
        RECT 294.665 46.930 294.920 47.220 ;
        RECT 295.090 46.670 295.420 47.050 ;
        RECT 295.590 46.930 295.760 49.050 ;
        RECT 295.930 48.250 296.255 49.035 ;
        RECT 296.425 48.760 296.675 49.220 ;
        RECT 296.845 48.720 297.095 49.050 ;
        RECT 297.310 48.720 297.990 49.050 ;
        RECT 296.845 48.590 297.015 48.720 ;
        RECT 296.620 48.420 297.015 48.590 ;
        RECT 295.990 47.200 296.450 48.250 ;
        RECT 296.620 47.060 296.790 48.420 ;
        RECT 297.185 48.160 297.650 48.550 ;
        RECT 296.960 47.350 297.310 47.970 ;
        RECT 297.480 47.570 297.650 48.160 ;
        RECT 297.820 47.940 297.990 48.720 ;
        RECT 298.160 48.620 298.330 48.960 ;
        RECT 298.565 48.790 298.895 49.220 ;
        RECT 299.065 48.620 299.235 48.960 ;
        RECT 299.530 48.760 299.900 49.220 ;
        RECT 298.160 48.450 299.235 48.620 ;
        RECT 300.070 48.590 300.240 49.050 ;
        RECT 300.475 48.710 301.345 49.050 ;
        RECT 301.515 48.760 301.765 49.220 ;
        RECT 299.680 48.420 300.240 48.590 ;
        RECT 299.680 48.280 299.850 48.420 ;
        RECT 298.350 48.110 299.850 48.280 ;
        RECT 300.545 48.250 301.005 48.540 ;
        RECT 297.820 47.770 299.510 47.940 ;
        RECT 297.480 47.350 297.835 47.570 ;
        RECT 298.005 47.060 298.175 47.770 ;
        RECT 298.380 47.350 299.170 47.600 ;
        RECT 299.340 47.590 299.510 47.770 ;
        RECT 299.680 47.420 299.850 48.110 ;
        RECT 296.120 46.670 296.450 47.030 ;
        RECT 296.620 46.890 297.115 47.060 ;
        RECT 297.320 46.890 298.175 47.060 ;
        RECT 299.050 46.670 299.380 47.130 ;
        RECT 299.590 47.030 299.850 47.420 ;
        RECT 300.040 48.240 301.005 48.250 ;
        RECT 301.175 48.330 301.345 48.710 ;
        RECT 301.935 48.670 302.105 48.960 ;
        RECT 302.285 48.840 302.615 49.220 ;
        RECT 301.935 48.500 302.735 48.670 ;
        RECT 300.040 48.080 300.715 48.240 ;
        RECT 301.175 48.160 302.395 48.330 ;
        RECT 300.040 47.290 300.250 48.080 ;
        RECT 301.175 48.070 301.345 48.160 ;
        RECT 300.420 47.290 300.770 47.910 ;
        RECT 300.940 47.900 301.345 48.070 ;
        RECT 300.940 47.120 301.110 47.900 ;
        RECT 301.280 47.450 301.500 47.730 ;
        RECT 301.680 47.620 302.220 47.990 ;
        RECT 302.565 47.910 302.735 48.500 ;
        RECT 302.955 48.080 303.260 49.220 ;
        RECT 303.430 48.030 303.685 48.910 ;
        RECT 303.860 48.055 304.150 49.220 ;
        RECT 304.320 48.080 304.705 49.050 ;
        RECT 304.875 48.760 305.200 49.220 ;
        RECT 305.720 48.590 306.000 49.050 ;
        RECT 304.875 48.370 306.000 48.590 ;
        RECT 302.565 47.880 303.305 47.910 ;
        RECT 301.280 47.280 301.810 47.450 ;
        RECT 299.590 46.860 299.940 47.030 ;
        RECT 300.160 46.840 301.110 47.120 ;
        RECT 301.280 46.670 301.470 47.110 ;
        RECT 301.640 47.050 301.810 47.280 ;
        RECT 301.980 47.220 302.220 47.620 ;
        RECT 302.390 47.580 303.305 47.880 ;
        RECT 302.390 47.405 302.715 47.580 ;
        RECT 302.390 47.050 302.710 47.405 ;
        RECT 303.475 47.380 303.685 48.030 ;
        RECT 304.320 47.410 304.600 48.080 ;
        RECT 304.875 47.910 305.325 48.370 ;
        RECT 306.190 48.200 306.590 49.050 ;
        RECT 306.990 48.760 307.260 49.220 ;
        RECT 307.430 48.590 307.715 49.050 ;
        RECT 304.770 47.580 305.325 47.910 ;
        RECT 305.495 47.640 306.590 48.200 ;
        RECT 304.875 47.470 305.325 47.580 ;
        RECT 301.640 46.880 302.710 47.050 ;
        RECT 302.955 46.670 303.260 47.130 ;
        RECT 303.430 46.850 303.685 47.380 ;
        RECT 303.860 46.670 304.150 47.395 ;
        RECT 304.320 46.840 304.705 47.410 ;
        RECT 304.875 47.300 306.000 47.470 ;
        RECT 304.875 46.670 305.200 47.130 ;
        RECT 305.720 46.840 306.000 47.300 ;
        RECT 306.190 46.840 306.590 47.640 ;
        RECT 306.760 48.370 307.715 48.590 ;
        RECT 306.760 47.470 306.970 48.370 ;
        RECT 307.140 47.640 307.830 48.200 ;
        RECT 308.000 48.130 309.670 49.220 ;
        RECT 306.760 47.300 307.715 47.470 ;
        RECT 306.990 46.670 307.260 47.130 ;
        RECT 307.430 46.840 307.715 47.300 ;
        RECT 308.000 47.440 308.750 47.960 ;
        RECT 308.920 47.610 309.670 48.130 ;
        RECT 309.840 48.130 311.050 49.220 ;
        RECT 309.840 47.590 310.360 48.130 ;
        RECT 308.000 46.670 309.670 47.440 ;
        RECT 310.530 47.420 311.050 47.960 ;
        RECT 309.840 46.670 311.050 47.420 ;
        RECT 162.095 46.500 311.135 46.670 ;
        RECT 162.180 45.750 163.390 46.500 ;
        RECT 163.560 45.955 168.905 46.500 ;
        RECT 162.180 45.210 162.700 45.750 ;
        RECT 162.870 45.040 163.390 45.580 ;
        RECT 165.145 45.125 165.485 45.955 ;
        RECT 169.080 45.730 172.590 46.500 ;
        RECT 173.680 45.760 174.065 46.330 ;
        RECT 174.235 46.040 174.560 46.500 ;
        RECT 175.080 45.870 175.360 46.330 ;
        RECT 162.180 43.950 163.390 45.040 ;
        RECT 166.965 44.385 167.315 45.635 ;
        RECT 169.080 45.210 170.730 45.730 ;
        RECT 170.900 45.040 172.590 45.560 ;
        RECT 163.560 43.950 168.905 44.385 ;
        RECT 169.080 43.950 172.590 45.040 ;
        RECT 173.680 45.090 173.960 45.760 ;
        RECT 174.235 45.700 175.360 45.870 ;
        RECT 174.235 45.590 174.685 45.700 ;
        RECT 174.130 45.260 174.685 45.590 ;
        RECT 175.550 45.530 175.950 46.330 ;
        RECT 176.350 46.040 176.620 46.500 ;
        RECT 176.790 45.870 177.075 46.330 ;
        RECT 173.680 44.120 174.065 45.090 ;
        RECT 174.235 44.800 174.685 45.260 ;
        RECT 174.855 44.970 175.950 45.530 ;
        RECT 174.235 44.580 175.360 44.800 ;
        RECT 174.235 43.950 174.560 44.410 ;
        RECT 175.080 44.120 175.360 44.580 ;
        RECT 175.550 44.120 175.950 44.970 ;
        RECT 176.120 45.700 177.075 45.870 ;
        RECT 177.365 45.950 177.620 46.240 ;
        RECT 177.790 46.120 178.120 46.500 ;
        RECT 177.365 45.780 178.115 45.950 ;
        RECT 176.120 44.800 176.330 45.700 ;
        RECT 176.500 44.970 177.190 45.530 ;
        RECT 177.365 44.960 177.715 45.610 ;
        RECT 176.120 44.580 177.075 44.800 ;
        RECT 177.885 44.790 178.115 45.780 ;
        RECT 176.350 43.950 176.620 44.410 ;
        RECT 176.790 44.120 177.075 44.580 ;
        RECT 177.365 44.620 178.115 44.790 ;
        RECT 177.365 44.120 177.620 44.620 ;
        RECT 177.790 43.950 178.120 44.450 ;
        RECT 178.290 44.120 178.460 46.240 ;
        RECT 178.820 46.140 179.150 46.500 ;
        RECT 179.320 46.110 179.815 46.280 ;
        RECT 180.020 46.110 180.875 46.280 ;
        RECT 178.690 44.920 179.150 45.970 ;
        RECT 178.630 44.135 178.955 44.920 ;
        RECT 179.320 44.750 179.490 46.110 ;
        RECT 179.660 45.200 180.010 45.820 ;
        RECT 180.180 45.600 180.535 45.820 ;
        RECT 180.180 45.010 180.350 45.600 ;
        RECT 180.705 45.400 180.875 46.110 ;
        RECT 181.750 46.040 182.080 46.500 ;
        RECT 182.290 46.140 182.640 46.310 ;
        RECT 181.080 45.570 181.870 45.820 ;
        RECT 182.290 45.750 182.550 46.140 ;
        RECT 182.860 46.050 183.810 46.330 ;
        RECT 183.980 46.060 184.170 46.500 ;
        RECT 184.340 46.120 185.410 46.290 ;
        RECT 182.040 45.400 182.210 45.580 ;
        RECT 179.320 44.580 179.715 44.750 ;
        RECT 179.885 44.620 180.350 45.010 ;
        RECT 180.520 45.230 182.210 45.400 ;
        RECT 179.545 44.450 179.715 44.580 ;
        RECT 180.520 44.450 180.690 45.230 ;
        RECT 182.380 45.060 182.550 45.750 ;
        RECT 181.050 44.890 182.550 45.060 ;
        RECT 182.740 45.090 182.950 45.880 ;
        RECT 183.120 45.260 183.470 45.880 ;
        RECT 183.640 45.270 183.810 46.050 ;
        RECT 184.340 45.890 184.510 46.120 ;
        RECT 183.980 45.720 184.510 45.890 ;
        RECT 183.980 45.440 184.200 45.720 ;
        RECT 184.680 45.550 184.920 45.950 ;
        RECT 183.640 45.100 184.045 45.270 ;
        RECT 184.380 45.180 184.920 45.550 ;
        RECT 185.090 45.765 185.410 46.120 ;
        RECT 185.090 45.510 185.415 45.765 ;
        RECT 185.610 45.690 185.780 46.500 ;
        RECT 185.950 45.850 186.280 46.330 ;
        RECT 186.450 46.030 186.620 46.500 ;
        RECT 186.790 45.850 187.120 46.330 ;
        RECT 187.290 46.030 187.460 46.500 ;
        RECT 185.950 45.680 187.715 45.850 ;
        RECT 187.940 45.775 188.230 46.500 ;
        RECT 185.090 45.300 187.120 45.510 ;
        RECT 185.090 45.290 185.435 45.300 ;
        RECT 182.740 44.930 183.415 45.090 ;
        RECT 183.875 45.010 184.045 45.100 ;
        RECT 182.740 44.920 183.705 44.930 ;
        RECT 182.380 44.750 182.550 44.890 ;
        RECT 179.125 43.950 179.375 44.410 ;
        RECT 179.545 44.120 179.795 44.450 ;
        RECT 180.010 44.120 180.690 44.450 ;
        RECT 180.860 44.550 181.935 44.720 ;
        RECT 182.380 44.580 182.940 44.750 ;
        RECT 183.245 44.630 183.705 44.920 ;
        RECT 183.875 44.840 185.095 45.010 ;
        RECT 180.860 44.210 181.030 44.550 ;
        RECT 181.265 43.950 181.595 44.380 ;
        RECT 181.765 44.210 181.935 44.550 ;
        RECT 182.230 43.950 182.600 44.410 ;
        RECT 182.770 44.120 182.940 44.580 ;
        RECT 183.875 44.460 184.045 44.840 ;
        RECT 185.265 44.670 185.435 45.290 ;
        RECT 187.305 45.130 187.715 45.680 ;
        RECT 183.175 44.120 184.045 44.460 ;
        RECT 184.635 44.500 185.435 44.670 ;
        RECT 184.215 43.950 184.465 44.410 ;
        RECT 184.635 44.210 184.805 44.500 ;
        RECT 184.985 43.950 185.315 44.330 ;
        RECT 185.610 43.950 185.780 45.010 ;
        RECT 185.990 44.960 187.715 45.130 ;
        RECT 188.405 45.760 188.660 46.330 ;
        RECT 188.830 46.100 189.160 46.500 ;
        RECT 189.585 45.965 190.115 46.330 ;
        RECT 189.585 45.930 189.760 45.965 ;
        RECT 188.830 45.760 189.760 45.930 ;
        RECT 190.305 45.820 190.580 46.330 ;
        RECT 185.990 44.120 186.280 44.960 ;
        RECT 186.450 43.950 186.620 44.790 ;
        RECT 186.830 44.120 187.080 44.960 ;
        RECT 187.290 43.950 187.460 44.790 ;
        RECT 187.940 43.950 188.230 45.115 ;
        RECT 188.405 45.090 188.575 45.760 ;
        RECT 188.830 45.590 189.000 45.760 ;
        RECT 188.745 45.260 189.000 45.590 ;
        RECT 189.225 45.260 189.420 45.590 ;
        RECT 188.405 44.120 188.740 45.090 ;
        RECT 188.910 43.950 189.080 45.090 ;
        RECT 189.250 44.290 189.420 45.260 ;
        RECT 189.590 44.630 189.760 45.760 ;
        RECT 189.930 44.970 190.100 45.770 ;
        RECT 190.300 45.650 190.580 45.820 ;
        RECT 190.305 45.170 190.580 45.650 ;
        RECT 190.750 44.970 190.940 46.330 ;
        RECT 191.120 45.965 191.630 46.500 ;
        RECT 191.850 45.690 192.095 46.295 ;
        RECT 193.465 45.760 193.720 46.330 ;
        RECT 193.890 46.100 194.220 46.500 ;
        RECT 194.645 45.965 195.175 46.330 ;
        RECT 195.365 46.160 195.640 46.330 ;
        RECT 195.360 45.990 195.640 46.160 ;
        RECT 194.645 45.930 194.820 45.965 ;
        RECT 193.890 45.760 194.820 45.930 ;
        RECT 191.140 45.520 192.370 45.690 ;
        RECT 189.930 44.800 190.940 44.970 ;
        RECT 191.110 44.955 191.860 45.145 ;
        RECT 189.590 44.460 190.715 44.630 ;
        RECT 191.110 44.290 191.280 44.955 ;
        RECT 192.030 44.710 192.370 45.520 ;
        RECT 189.250 44.120 191.280 44.290 ;
        RECT 191.450 43.950 191.620 44.710 ;
        RECT 191.855 44.300 192.370 44.710 ;
        RECT 193.465 45.090 193.635 45.760 ;
        RECT 193.890 45.590 194.060 45.760 ;
        RECT 193.805 45.260 194.060 45.590 ;
        RECT 194.285 45.260 194.480 45.590 ;
        RECT 193.465 44.120 193.800 45.090 ;
        RECT 193.970 43.950 194.140 45.090 ;
        RECT 194.310 44.290 194.480 45.260 ;
        RECT 194.650 44.630 194.820 45.760 ;
        RECT 194.990 44.970 195.160 45.770 ;
        RECT 195.365 45.170 195.640 45.990 ;
        RECT 195.810 44.970 196.000 46.330 ;
        RECT 196.180 45.965 196.690 46.500 ;
        RECT 196.910 45.690 197.155 46.295 ;
        RECT 197.600 45.730 199.270 46.500 ;
        RECT 199.905 45.950 200.160 46.240 ;
        RECT 200.330 46.120 200.660 46.500 ;
        RECT 199.905 45.780 200.655 45.950 ;
        RECT 196.200 45.520 197.430 45.690 ;
        RECT 194.990 44.800 196.000 44.970 ;
        RECT 196.170 44.955 196.920 45.145 ;
        RECT 194.650 44.460 195.775 44.630 ;
        RECT 196.170 44.290 196.340 44.955 ;
        RECT 197.090 44.710 197.430 45.520 ;
        RECT 197.600 45.210 198.350 45.730 ;
        RECT 198.520 45.040 199.270 45.560 ;
        RECT 194.310 44.120 196.340 44.290 ;
        RECT 196.510 43.950 196.680 44.710 ;
        RECT 196.915 44.300 197.430 44.710 ;
        RECT 197.600 43.950 199.270 45.040 ;
        RECT 199.905 44.960 200.255 45.610 ;
        RECT 200.425 44.790 200.655 45.780 ;
        RECT 199.905 44.620 200.655 44.790 ;
        RECT 199.905 44.120 200.160 44.620 ;
        RECT 200.330 43.950 200.660 44.450 ;
        RECT 200.830 44.120 201.000 46.240 ;
        RECT 201.360 46.140 201.690 46.500 ;
        RECT 201.860 46.110 202.355 46.280 ;
        RECT 202.560 46.110 203.415 46.280 ;
        RECT 201.230 44.920 201.690 45.970 ;
        RECT 201.170 44.135 201.495 44.920 ;
        RECT 201.860 44.750 202.030 46.110 ;
        RECT 202.200 45.200 202.550 45.820 ;
        RECT 202.720 45.600 203.075 45.820 ;
        RECT 202.720 45.010 202.890 45.600 ;
        RECT 203.245 45.400 203.415 46.110 ;
        RECT 204.290 46.040 204.620 46.500 ;
        RECT 204.830 46.140 205.180 46.310 ;
        RECT 203.620 45.570 204.410 45.820 ;
        RECT 204.830 45.750 205.090 46.140 ;
        RECT 205.400 46.050 206.350 46.330 ;
        RECT 206.520 46.060 206.710 46.500 ;
        RECT 206.880 46.120 207.950 46.290 ;
        RECT 204.580 45.400 204.750 45.580 ;
        RECT 201.860 44.580 202.255 44.750 ;
        RECT 202.425 44.620 202.890 45.010 ;
        RECT 203.060 45.230 204.750 45.400 ;
        RECT 202.085 44.450 202.255 44.580 ;
        RECT 203.060 44.450 203.230 45.230 ;
        RECT 204.920 45.060 205.090 45.750 ;
        RECT 203.590 44.890 205.090 45.060 ;
        RECT 205.280 45.090 205.490 45.880 ;
        RECT 205.660 45.260 206.010 45.880 ;
        RECT 206.180 45.270 206.350 46.050 ;
        RECT 206.880 45.890 207.050 46.120 ;
        RECT 206.520 45.720 207.050 45.890 ;
        RECT 206.520 45.440 206.740 45.720 ;
        RECT 207.220 45.550 207.460 45.950 ;
        RECT 206.180 45.100 206.585 45.270 ;
        RECT 206.920 45.180 207.460 45.550 ;
        RECT 207.630 45.765 207.950 46.120 ;
        RECT 207.630 45.510 207.955 45.765 ;
        RECT 208.150 45.690 208.320 46.500 ;
        RECT 208.490 45.850 208.820 46.330 ;
        RECT 208.990 46.030 209.160 46.500 ;
        RECT 209.330 45.850 209.660 46.330 ;
        RECT 209.830 46.030 210.000 46.500 ;
        RECT 208.490 45.680 210.255 45.850 ;
        RECT 207.630 45.300 209.660 45.510 ;
        RECT 207.630 45.290 207.975 45.300 ;
        RECT 205.280 44.930 205.955 45.090 ;
        RECT 206.415 45.010 206.585 45.100 ;
        RECT 205.280 44.920 206.245 44.930 ;
        RECT 204.920 44.750 205.090 44.890 ;
        RECT 201.665 43.950 201.915 44.410 ;
        RECT 202.085 44.120 202.335 44.450 ;
        RECT 202.550 44.120 203.230 44.450 ;
        RECT 203.400 44.550 204.475 44.720 ;
        RECT 204.920 44.580 205.480 44.750 ;
        RECT 205.785 44.630 206.245 44.920 ;
        RECT 206.415 44.840 207.635 45.010 ;
        RECT 203.400 44.210 203.570 44.550 ;
        RECT 203.805 43.950 204.135 44.380 ;
        RECT 204.305 44.210 204.475 44.550 ;
        RECT 204.770 43.950 205.140 44.410 ;
        RECT 205.310 44.120 205.480 44.580 ;
        RECT 206.415 44.460 206.585 44.840 ;
        RECT 207.805 44.670 207.975 45.290 ;
        RECT 209.845 45.130 210.255 45.680 ;
        RECT 210.480 45.730 213.070 46.500 ;
        RECT 213.700 45.775 213.990 46.500 ;
        RECT 215.080 46.000 215.340 46.330 ;
        RECT 215.550 46.020 215.825 46.500 ;
        RECT 210.480 45.210 211.690 45.730 ;
        RECT 205.715 44.120 206.585 44.460 ;
        RECT 207.175 44.500 207.975 44.670 ;
        RECT 206.755 43.950 207.005 44.410 ;
        RECT 207.175 44.210 207.345 44.500 ;
        RECT 207.525 43.950 207.855 44.330 ;
        RECT 208.150 43.950 208.320 45.010 ;
        RECT 208.530 44.960 210.255 45.130 ;
        RECT 211.860 45.040 213.070 45.560 ;
        RECT 208.530 44.120 208.820 44.960 ;
        RECT 208.990 43.950 209.160 44.790 ;
        RECT 209.370 44.120 209.620 44.960 ;
        RECT 209.830 43.950 210.000 44.790 ;
        RECT 210.480 43.950 213.070 45.040 ;
        RECT 213.700 43.950 213.990 45.115 ;
        RECT 215.080 45.090 215.250 46.000 ;
        RECT 216.035 45.930 216.240 46.330 ;
        RECT 216.410 46.100 216.745 46.500 ;
        RECT 215.420 45.260 215.780 45.840 ;
        RECT 216.035 45.760 216.720 45.930 ;
        RECT 215.960 45.090 216.210 45.590 ;
        RECT 215.080 44.920 216.210 45.090 ;
        RECT 215.080 44.150 215.350 44.920 ;
        RECT 216.380 44.730 216.720 45.760 ;
        RECT 216.960 45.680 217.190 46.500 ;
        RECT 217.360 45.700 217.690 46.330 ;
        RECT 216.940 45.260 217.270 45.510 ;
        RECT 217.440 45.100 217.690 45.700 ;
        RECT 217.860 45.680 218.070 46.500 ;
        RECT 218.300 45.750 219.510 46.500 ;
        RECT 219.685 45.950 219.940 46.240 ;
        RECT 220.110 46.120 220.440 46.500 ;
        RECT 219.685 45.780 220.435 45.950 ;
        RECT 218.300 45.210 218.820 45.750 ;
        RECT 215.520 43.950 215.850 44.730 ;
        RECT 216.055 44.555 216.720 44.730 ;
        RECT 216.055 44.150 216.240 44.555 ;
        RECT 216.410 43.950 216.745 44.375 ;
        RECT 216.960 43.950 217.190 45.090 ;
        RECT 217.360 44.120 217.690 45.100 ;
        RECT 217.860 43.950 218.070 45.090 ;
        RECT 218.990 45.040 219.510 45.580 ;
        RECT 218.300 43.950 219.510 45.040 ;
        RECT 219.685 44.960 220.035 45.610 ;
        RECT 220.205 44.790 220.435 45.780 ;
        RECT 219.685 44.620 220.435 44.790 ;
        RECT 219.685 44.120 219.940 44.620 ;
        RECT 220.110 43.950 220.440 44.450 ;
        RECT 220.610 44.120 220.780 46.240 ;
        RECT 221.140 46.140 221.470 46.500 ;
        RECT 221.640 46.110 222.135 46.280 ;
        RECT 222.340 46.110 223.195 46.280 ;
        RECT 221.010 44.920 221.470 45.970 ;
        RECT 220.950 44.135 221.275 44.920 ;
        RECT 221.640 44.750 221.810 46.110 ;
        RECT 221.980 45.200 222.330 45.820 ;
        RECT 222.500 45.600 222.855 45.820 ;
        RECT 222.500 45.010 222.670 45.600 ;
        RECT 223.025 45.400 223.195 46.110 ;
        RECT 224.070 46.040 224.400 46.500 ;
        RECT 224.610 46.140 224.960 46.310 ;
        RECT 223.400 45.570 224.190 45.820 ;
        RECT 224.610 45.750 224.870 46.140 ;
        RECT 225.180 46.050 226.130 46.330 ;
        RECT 226.300 46.060 226.490 46.500 ;
        RECT 226.660 46.120 227.730 46.290 ;
        RECT 224.360 45.400 224.530 45.580 ;
        RECT 221.640 44.580 222.035 44.750 ;
        RECT 222.205 44.620 222.670 45.010 ;
        RECT 222.840 45.230 224.530 45.400 ;
        RECT 221.865 44.450 222.035 44.580 ;
        RECT 222.840 44.450 223.010 45.230 ;
        RECT 224.700 45.060 224.870 45.750 ;
        RECT 223.370 44.890 224.870 45.060 ;
        RECT 225.060 45.090 225.270 45.880 ;
        RECT 225.440 45.260 225.790 45.880 ;
        RECT 225.960 45.270 226.130 46.050 ;
        RECT 226.660 45.890 226.830 46.120 ;
        RECT 226.300 45.720 226.830 45.890 ;
        RECT 226.300 45.440 226.520 45.720 ;
        RECT 227.000 45.550 227.240 45.950 ;
        RECT 225.960 45.100 226.365 45.270 ;
        RECT 226.700 45.180 227.240 45.550 ;
        RECT 227.410 45.765 227.730 46.120 ;
        RECT 227.410 45.510 227.735 45.765 ;
        RECT 227.930 45.690 228.100 46.500 ;
        RECT 228.270 45.850 228.600 46.330 ;
        RECT 228.770 46.030 228.940 46.500 ;
        RECT 229.110 45.850 229.440 46.330 ;
        RECT 229.610 46.030 229.780 46.500 ;
        RECT 230.260 46.000 230.560 46.330 ;
        RECT 230.730 46.020 231.005 46.500 ;
        RECT 228.270 45.680 230.035 45.850 ;
        RECT 227.410 45.300 229.440 45.510 ;
        RECT 227.410 45.290 227.755 45.300 ;
        RECT 225.060 44.930 225.735 45.090 ;
        RECT 226.195 45.010 226.365 45.100 ;
        RECT 225.060 44.920 226.025 44.930 ;
        RECT 224.700 44.750 224.870 44.890 ;
        RECT 221.445 43.950 221.695 44.410 ;
        RECT 221.865 44.120 222.115 44.450 ;
        RECT 222.330 44.120 223.010 44.450 ;
        RECT 223.180 44.550 224.255 44.720 ;
        RECT 224.700 44.580 225.260 44.750 ;
        RECT 225.565 44.630 226.025 44.920 ;
        RECT 226.195 44.840 227.415 45.010 ;
        RECT 223.180 44.210 223.350 44.550 ;
        RECT 223.585 43.950 223.915 44.380 ;
        RECT 224.085 44.210 224.255 44.550 ;
        RECT 224.550 43.950 224.920 44.410 ;
        RECT 225.090 44.120 225.260 44.580 ;
        RECT 226.195 44.460 226.365 44.840 ;
        RECT 227.585 44.670 227.755 45.290 ;
        RECT 229.625 45.130 230.035 45.680 ;
        RECT 225.495 44.120 226.365 44.460 ;
        RECT 226.955 44.500 227.755 44.670 ;
        RECT 226.535 43.950 226.785 44.410 ;
        RECT 226.955 44.210 227.125 44.500 ;
        RECT 227.305 43.950 227.635 44.330 ;
        RECT 227.930 43.950 228.100 45.010 ;
        RECT 228.310 44.960 230.035 45.130 ;
        RECT 230.260 45.090 230.430 46.000 ;
        RECT 231.185 45.850 231.480 46.240 ;
        RECT 231.650 46.020 231.905 46.500 ;
        RECT 232.080 45.850 232.340 46.240 ;
        RECT 232.510 46.020 232.790 46.500 ;
        RECT 233.020 45.955 238.365 46.500 ;
        RECT 230.600 45.260 230.950 45.830 ;
        RECT 231.185 45.680 232.835 45.850 ;
        RECT 231.120 45.340 232.260 45.510 ;
        RECT 231.120 45.090 231.290 45.340 ;
        RECT 232.430 45.170 232.835 45.680 ;
        RECT 228.310 44.120 228.600 44.960 ;
        RECT 228.770 43.950 228.940 44.790 ;
        RECT 229.150 44.120 229.400 44.960 ;
        RECT 230.260 44.920 231.290 45.090 ;
        RECT 232.080 45.000 232.835 45.170 ;
        RECT 234.605 45.125 234.945 45.955 ;
        RECT 239.460 45.775 239.750 46.500 ;
        RECT 239.920 45.730 243.430 46.500 ;
        RECT 243.605 45.950 243.860 46.240 ;
        RECT 244.030 46.120 244.360 46.500 ;
        RECT 243.605 45.780 244.355 45.950 ;
        RECT 229.610 43.950 229.780 44.790 ;
        RECT 230.260 44.120 230.570 44.920 ;
        RECT 232.080 44.750 232.340 45.000 ;
        RECT 230.740 43.950 231.050 44.750 ;
        RECT 231.220 44.580 232.340 44.750 ;
        RECT 231.220 44.120 231.480 44.580 ;
        RECT 231.650 43.950 231.905 44.410 ;
        RECT 232.080 44.120 232.340 44.580 ;
        RECT 232.510 43.950 232.795 44.820 ;
        RECT 236.425 44.385 236.775 45.635 ;
        RECT 239.920 45.210 241.570 45.730 ;
        RECT 233.020 43.950 238.365 44.385 ;
        RECT 239.460 43.950 239.750 45.115 ;
        RECT 241.740 45.040 243.430 45.560 ;
        RECT 239.920 43.950 243.430 45.040 ;
        RECT 243.605 44.960 243.955 45.610 ;
        RECT 244.125 44.790 244.355 45.780 ;
        RECT 243.605 44.620 244.355 44.790 ;
        RECT 243.605 44.120 243.860 44.620 ;
        RECT 244.030 43.950 244.360 44.450 ;
        RECT 244.530 44.120 244.700 46.240 ;
        RECT 245.060 46.140 245.390 46.500 ;
        RECT 245.560 46.110 246.055 46.280 ;
        RECT 246.260 46.110 247.115 46.280 ;
        RECT 244.930 44.920 245.390 45.970 ;
        RECT 244.870 44.135 245.195 44.920 ;
        RECT 245.560 44.750 245.730 46.110 ;
        RECT 245.900 45.200 246.250 45.820 ;
        RECT 246.420 45.600 246.775 45.820 ;
        RECT 246.420 45.010 246.590 45.600 ;
        RECT 246.945 45.400 247.115 46.110 ;
        RECT 247.990 46.040 248.320 46.500 ;
        RECT 248.530 46.140 248.880 46.310 ;
        RECT 247.320 45.570 248.110 45.820 ;
        RECT 248.530 45.750 248.790 46.140 ;
        RECT 249.100 46.050 250.050 46.330 ;
        RECT 250.220 46.060 250.410 46.500 ;
        RECT 250.580 46.120 251.650 46.290 ;
        RECT 248.280 45.400 248.450 45.580 ;
        RECT 245.560 44.580 245.955 44.750 ;
        RECT 246.125 44.620 246.590 45.010 ;
        RECT 246.760 45.230 248.450 45.400 ;
        RECT 245.785 44.450 245.955 44.580 ;
        RECT 246.760 44.450 246.930 45.230 ;
        RECT 248.620 45.060 248.790 45.750 ;
        RECT 247.290 44.890 248.790 45.060 ;
        RECT 248.980 45.090 249.190 45.880 ;
        RECT 249.360 45.260 249.710 45.880 ;
        RECT 249.880 45.270 250.050 46.050 ;
        RECT 250.580 45.890 250.750 46.120 ;
        RECT 250.220 45.720 250.750 45.890 ;
        RECT 250.220 45.440 250.440 45.720 ;
        RECT 250.920 45.550 251.160 45.950 ;
        RECT 249.880 45.100 250.285 45.270 ;
        RECT 250.620 45.180 251.160 45.550 ;
        RECT 251.330 45.765 251.650 46.120 ;
        RECT 251.895 46.040 252.200 46.500 ;
        RECT 252.370 45.790 252.625 46.320 ;
        RECT 251.330 45.590 251.655 45.765 ;
        RECT 251.330 45.290 252.245 45.590 ;
        RECT 251.505 45.260 252.245 45.290 ;
        RECT 248.980 44.930 249.655 45.090 ;
        RECT 250.115 45.010 250.285 45.100 ;
        RECT 248.980 44.920 249.945 44.930 ;
        RECT 248.620 44.750 248.790 44.890 ;
        RECT 245.365 43.950 245.615 44.410 ;
        RECT 245.785 44.120 246.035 44.450 ;
        RECT 246.250 44.120 246.930 44.450 ;
        RECT 247.100 44.550 248.175 44.720 ;
        RECT 248.620 44.580 249.180 44.750 ;
        RECT 249.485 44.630 249.945 44.920 ;
        RECT 250.115 44.840 251.335 45.010 ;
        RECT 247.100 44.210 247.270 44.550 ;
        RECT 247.505 43.950 247.835 44.380 ;
        RECT 248.005 44.210 248.175 44.550 ;
        RECT 248.470 43.950 248.840 44.410 ;
        RECT 249.010 44.120 249.180 44.580 ;
        RECT 250.115 44.460 250.285 44.840 ;
        RECT 251.505 44.670 251.675 45.260 ;
        RECT 252.415 45.140 252.625 45.790 ;
        RECT 249.415 44.120 250.285 44.460 ;
        RECT 250.875 44.500 251.675 44.670 ;
        RECT 250.455 43.950 250.705 44.410 ;
        RECT 250.875 44.210 251.045 44.500 ;
        RECT 251.225 43.950 251.555 44.330 ;
        RECT 251.895 43.950 252.200 45.090 ;
        RECT 252.370 44.260 252.625 45.140 ;
        RECT 253.260 45.760 253.645 46.330 ;
        RECT 253.815 46.040 254.140 46.500 ;
        RECT 254.660 45.870 254.940 46.330 ;
        RECT 253.260 45.090 253.540 45.760 ;
        RECT 253.815 45.700 254.940 45.870 ;
        RECT 253.815 45.590 254.265 45.700 ;
        RECT 253.710 45.260 254.265 45.590 ;
        RECT 255.130 45.530 255.530 46.330 ;
        RECT 255.930 46.040 256.200 46.500 ;
        RECT 256.370 45.870 256.655 46.330 ;
        RECT 253.260 44.120 253.645 45.090 ;
        RECT 253.815 44.800 254.265 45.260 ;
        RECT 254.435 44.970 255.530 45.530 ;
        RECT 253.815 44.580 254.940 44.800 ;
        RECT 253.815 43.950 254.140 44.410 ;
        RECT 254.660 44.120 254.940 44.580 ;
        RECT 255.130 44.120 255.530 44.970 ;
        RECT 255.700 45.700 256.655 45.870 ;
        RECT 256.940 46.040 257.500 46.330 ;
        RECT 257.670 46.040 257.920 46.500 ;
        RECT 255.700 44.800 255.910 45.700 ;
        RECT 256.080 44.970 256.770 45.530 ;
        RECT 255.700 44.580 256.655 44.800 ;
        RECT 255.930 43.950 256.200 44.410 ;
        RECT 256.370 44.120 256.655 44.580 ;
        RECT 256.940 44.670 257.190 46.040 ;
        RECT 258.540 45.870 258.870 46.230 ;
        RECT 260.405 46.020 260.705 46.500 ;
        RECT 257.480 45.680 258.870 45.870 ;
        RECT 260.875 45.850 261.135 46.305 ;
        RECT 261.305 46.020 261.565 46.500 ;
        RECT 261.735 45.850 261.995 46.305 ;
        RECT 262.165 46.020 262.425 46.500 ;
        RECT 262.595 45.850 262.855 46.305 ;
        RECT 263.025 46.020 263.285 46.500 ;
        RECT 263.455 45.850 263.715 46.305 ;
        RECT 263.885 45.975 264.145 46.500 ;
        RECT 260.405 45.680 263.715 45.850 ;
        RECT 257.480 45.590 257.650 45.680 ;
        RECT 257.360 45.260 257.650 45.590 ;
        RECT 257.820 45.260 258.160 45.510 ;
        RECT 258.380 45.260 259.055 45.510 ;
        RECT 257.480 45.010 257.650 45.260 ;
        RECT 257.480 44.840 258.420 45.010 ;
        RECT 258.790 44.900 259.055 45.260 ;
        RECT 260.405 45.090 261.375 45.680 ;
        RECT 264.315 45.510 264.565 46.320 ;
        RECT 264.745 46.040 264.990 46.500 ;
        RECT 261.545 45.260 264.565 45.510 ;
        RECT 264.735 45.260 265.050 45.870 ;
        RECT 265.220 45.775 265.510 46.500 ;
        RECT 265.680 45.760 266.065 46.330 ;
        RECT 266.235 46.040 266.560 46.500 ;
        RECT 267.080 45.870 267.360 46.330 ;
        RECT 260.405 44.850 263.715 45.090 ;
        RECT 256.940 44.120 257.400 44.670 ;
        RECT 257.590 43.950 257.920 44.670 ;
        RECT 258.120 44.290 258.420 44.840 ;
        RECT 258.590 43.950 258.870 44.620 ;
        RECT 260.410 43.950 260.705 44.680 ;
        RECT 260.875 44.125 261.135 44.850 ;
        RECT 261.305 43.950 261.565 44.680 ;
        RECT 261.735 44.125 261.995 44.850 ;
        RECT 262.165 43.950 262.425 44.680 ;
        RECT 262.595 44.125 262.855 44.850 ;
        RECT 263.025 43.950 263.285 44.680 ;
        RECT 263.455 44.125 263.715 44.850 ;
        RECT 263.885 43.950 264.145 45.060 ;
        RECT 264.315 44.125 264.565 45.260 ;
        RECT 264.745 43.950 265.040 45.060 ;
        RECT 265.220 43.950 265.510 45.115 ;
        RECT 265.680 45.090 265.960 45.760 ;
        RECT 266.235 45.700 267.360 45.870 ;
        RECT 266.235 45.590 266.685 45.700 ;
        RECT 266.130 45.260 266.685 45.590 ;
        RECT 267.550 45.530 267.950 46.330 ;
        RECT 268.350 46.040 268.620 46.500 ;
        RECT 268.790 45.870 269.075 46.330 ;
        RECT 265.680 44.120 266.065 45.090 ;
        RECT 266.235 44.800 266.685 45.260 ;
        RECT 266.855 44.970 267.950 45.530 ;
        RECT 266.235 44.580 267.360 44.800 ;
        RECT 266.235 43.950 266.560 44.410 ;
        RECT 267.080 44.120 267.360 44.580 ;
        RECT 267.550 44.120 267.950 44.970 ;
        RECT 268.120 45.700 269.075 45.870 ;
        RECT 269.560 45.870 269.890 46.230 ;
        RECT 270.510 46.040 270.760 46.500 ;
        RECT 270.930 46.040 271.490 46.330 ;
        RECT 268.120 44.800 268.330 45.700 ;
        RECT 269.560 45.680 270.950 45.870 ;
        RECT 270.780 45.590 270.950 45.680 ;
        RECT 268.500 44.970 269.190 45.530 ;
        RECT 269.375 45.260 270.050 45.510 ;
        RECT 270.270 45.260 270.610 45.510 ;
        RECT 270.780 45.260 271.070 45.590 ;
        RECT 269.375 44.900 269.640 45.260 ;
        RECT 270.780 45.010 270.950 45.260 ;
        RECT 270.010 44.840 270.950 45.010 ;
        RECT 268.120 44.580 269.075 44.800 ;
        RECT 268.350 43.950 268.620 44.410 ;
        RECT 268.790 44.120 269.075 44.580 ;
        RECT 269.560 43.950 269.840 44.620 ;
        RECT 270.010 44.290 270.310 44.840 ;
        RECT 271.240 44.670 271.490 46.040 ;
        RECT 272.585 45.950 272.840 46.240 ;
        RECT 273.010 46.120 273.340 46.500 ;
        RECT 272.585 45.780 273.335 45.950 ;
        RECT 272.585 44.960 272.935 45.610 ;
        RECT 273.105 44.790 273.335 45.780 ;
        RECT 270.510 43.950 270.840 44.670 ;
        RECT 271.030 44.120 271.490 44.670 ;
        RECT 272.585 44.620 273.335 44.790 ;
        RECT 272.585 44.120 272.840 44.620 ;
        RECT 273.010 43.950 273.340 44.450 ;
        RECT 273.510 44.120 273.680 46.240 ;
        RECT 274.040 46.140 274.370 46.500 ;
        RECT 274.540 46.110 275.035 46.280 ;
        RECT 275.240 46.110 276.095 46.280 ;
        RECT 273.910 44.920 274.370 45.970 ;
        RECT 273.850 44.135 274.175 44.920 ;
        RECT 274.540 44.750 274.710 46.110 ;
        RECT 274.880 45.200 275.230 45.820 ;
        RECT 275.400 45.600 275.755 45.820 ;
        RECT 275.400 45.010 275.570 45.600 ;
        RECT 275.925 45.400 276.095 46.110 ;
        RECT 276.970 46.040 277.300 46.500 ;
        RECT 277.510 46.140 277.860 46.310 ;
        RECT 276.300 45.570 277.090 45.820 ;
        RECT 277.510 45.750 277.770 46.140 ;
        RECT 278.080 46.050 279.030 46.330 ;
        RECT 279.200 46.060 279.390 46.500 ;
        RECT 279.560 46.120 280.630 46.290 ;
        RECT 277.260 45.400 277.430 45.580 ;
        RECT 274.540 44.580 274.935 44.750 ;
        RECT 275.105 44.620 275.570 45.010 ;
        RECT 275.740 45.230 277.430 45.400 ;
        RECT 274.765 44.450 274.935 44.580 ;
        RECT 275.740 44.450 275.910 45.230 ;
        RECT 277.600 45.060 277.770 45.750 ;
        RECT 276.270 44.890 277.770 45.060 ;
        RECT 277.960 45.090 278.170 45.880 ;
        RECT 278.340 45.260 278.690 45.880 ;
        RECT 278.860 45.270 279.030 46.050 ;
        RECT 279.560 45.890 279.730 46.120 ;
        RECT 279.200 45.720 279.730 45.890 ;
        RECT 279.200 45.440 279.420 45.720 ;
        RECT 279.900 45.550 280.140 45.950 ;
        RECT 278.860 45.100 279.265 45.270 ;
        RECT 279.600 45.180 280.140 45.550 ;
        RECT 280.310 45.765 280.630 46.120 ;
        RECT 280.875 46.040 281.180 46.500 ;
        RECT 281.350 45.790 281.605 46.320 ;
        RECT 280.310 45.590 280.635 45.765 ;
        RECT 280.310 45.290 281.225 45.590 ;
        RECT 280.485 45.260 281.225 45.290 ;
        RECT 277.960 44.930 278.635 45.090 ;
        RECT 279.095 45.010 279.265 45.100 ;
        RECT 277.960 44.920 278.925 44.930 ;
        RECT 277.600 44.750 277.770 44.890 ;
        RECT 274.345 43.950 274.595 44.410 ;
        RECT 274.765 44.120 275.015 44.450 ;
        RECT 275.230 44.120 275.910 44.450 ;
        RECT 276.080 44.550 277.155 44.720 ;
        RECT 277.600 44.580 278.160 44.750 ;
        RECT 278.465 44.630 278.925 44.920 ;
        RECT 279.095 44.840 280.315 45.010 ;
        RECT 276.080 44.210 276.250 44.550 ;
        RECT 276.485 43.950 276.815 44.380 ;
        RECT 276.985 44.210 277.155 44.550 ;
        RECT 277.450 43.950 277.820 44.410 ;
        RECT 277.990 44.120 278.160 44.580 ;
        RECT 279.095 44.460 279.265 44.840 ;
        RECT 280.485 44.670 280.655 45.260 ;
        RECT 281.395 45.140 281.605 45.790 ;
        RECT 278.395 44.120 279.265 44.460 ;
        RECT 279.855 44.500 280.655 44.670 ;
        RECT 279.435 43.950 279.685 44.410 ;
        RECT 279.855 44.210 280.025 44.500 ;
        RECT 280.205 43.950 280.535 44.330 ;
        RECT 280.875 43.950 281.180 45.090 ;
        RECT 281.350 44.260 281.605 45.140 ;
        RECT 281.785 45.790 282.040 46.320 ;
        RECT 282.210 46.040 282.515 46.500 ;
        RECT 282.760 46.120 283.830 46.290 ;
        RECT 281.785 45.140 281.995 45.790 ;
        RECT 282.760 45.765 283.080 46.120 ;
        RECT 282.755 45.590 283.080 45.765 ;
        RECT 282.165 45.290 283.080 45.590 ;
        RECT 283.250 45.550 283.490 45.950 ;
        RECT 283.660 45.890 283.830 46.120 ;
        RECT 284.000 46.060 284.190 46.500 ;
        RECT 284.360 46.050 285.310 46.330 ;
        RECT 285.530 46.140 285.880 46.310 ;
        RECT 283.660 45.720 284.190 45.890 ;
        RECT 282.165 45.260 282.905 45.290 ;
        RECT 281.785 44.260 282.040 45.140 ;
        RECT 282.210 43.950 282.515 45.090 ;
        RECT 282.735 44.670 282.905 45.260 ;
        RECT 283.250 45.180 283.790 45.550 ;
        RECT 283.970 45.440 284.190 45.720 ;
        RECT 284.360 45.270 284.530 46.050 ;
        RECT 284.125 45.100 284.530 45.270 ;
        RECT 284.700 45.260 285.050 45.880 ;
        RECT 284.125 45.010 284.295 45.100 ;
        RECT 285.220 45.090 285.430 45.880 ;
        RECT 283.075 44.840 284.295 45.010 ;
        RECT 284.755 44.930 285.430 45.090 ;
        RECT 282.735 44.500 283.535 44.670 ;
        RECT 282.855 43.950 283.185 44.330 ;
        RECT 283.365 44.210 283.535 44.500 ;
        RECT 284.125 44.460 284.295 44.840 ;
        RECT 284.465 44.920 285.430 44.930 ;
        RECT 285.620 45.750 285.880 46.140 ;
        RECT 286.090 46.040 286.420 46.500 ;
        RECT 287.295 46.110 288.150 46.280 ;
        RECT 288.355 46.110 288.850 46.280 ;
        RECT 289.020 46.140 289.350 46.500 ;
        RECT 285.620 45.060 285.790 45.750 ;
        RECT 285.960 45.400 286.130 45.580 ;
        RECT 286.300 45.570 287.090 45.820 ;
        RECT 287.295 45.400 287.465 46.110 ;
        RECT 287.635 45.600 287.990 45.820 ;
        RECT 285.960 45.230 287.650 45.400 ;
        RECT 284.465 44.630 284.925 44.920 ;
        RECT 285.620 44.890 287.120 45.060 ;
        RECT 285.620 44.750 285.790 44.890 ;
        RECT 285.230 44.580 285.790 44.750 ;
        RECT 283.705 43.950 283.955 44.410 ;
        RECT 284.125 44.120 284.995 44.460 ;
        RECT 285.230 44.120 285.400 44.580 ;
        RECT 286.235 44.550 287.310 44.720 ;
        RECT 285.570 43.950 285.940 44.410 ;
        RECT 286.235 44.210 286.405 44.550 ;
        RECT 286.575 43.950 286.905 44.380 ;
        RECT 287.140 44.210 287.310 44.550 ;
        RECT 287.480 44.450 287.650 45.230 ;
        RECT 287.820 45.010 287.990 45.600 ;
        RECT 288.160 45.200 288.510 45.820 ;
        RECT 287.820 44.620 288.285 45.010 ;
        RECT 288.680 44.750 288.850 46.110 ;
        RECT 289.020 44.920 289.480 45.970 ;
        RECT 288.455 44.580 288.850 44.750 ;
        RECT 288.455 44.450 288.625 44.580 ;
        RECT 287.480 44.120 288.160 44.450 ;
        RECT 288.375 44.120 288.625 44.450 ;
        RECT 288.795 43.950 289.045 44.410 ;
        RECT 289.215 44.135 289.540 44.920 ;
        RECT 289.710 44.120 289.880 46.240 ;
        RECT 290.050 46.120 290.380 46.500 ;
        RECT 290.550 45.950 290.805 46.240 ;
        RECT 290.055 45.780 290.805 45.950 ;
        RECT 290.055 44.790 290.285 45.780 ;
        RECT 290.980 45.775 291.270 46.500 ;
        RECT 291.530 45.850 291.700 46.330 ;
        RECT 291.870 46.020 292.200 46.500 ;
        RECT 292.425 46.080 293.960 46.330 ;
        RECT 292.425 45.850 292.595 46.080 ;
        RECT 291.530 45.680 292.595 45.850 ;
        RECT 290.455 44.960 290.805 45.610 ;
        RECT 292.775 45.510 293.055 45.910 ;
        RECT 291.445 45.300 291.795 45.510 ;
        RECT 291.965 45.310 292.410 45.510 ;
        RECT 292.580 45.310 293.055 45.510 ;
        RECT 293.325 45.510 293.610 45.910 ;
        RECT 293.790 45.850 293.960 46.080 ;
        RECT 294.130 46.020 294.460 46.500 ;
        RECT 294.675 46.000 294.930 46.330 ;
        RECT 294.745 45.920 294.930 46.000 ;
        RECT 293.790 45.680 294.590 45.850 ;
        RECT 293.325 45.310 293.655 45.510 ;
        RECT 293.825 45.310 294.190 45.510 ;
        RECT 294.420 45.130 294.590 45.680 ;
        RECT 290.055 44.620 290.805 44.790 ;
        RECT 290.050 43.950 290.380 44.450 ;
        RECT 290.550 44.120 290.805 44.620 ;
        RECT 290.980 43.950 291.270 45.115 ;
        RECT 291.530 44.960 294.590 45.130 ;
        RECT 291.530 44.120 291.700 44.960 ;
        RECT 294.760 44.800 294.930 45.920 ;
        RECT 295.695 45.870 295.980 46.330 ;
        RECT 296.150 46.040 296.420 46.500 ;
        RECT 295.695 45.700 296.650 45.870 ;
        RECT 295.580 44.970 296.270 45.530 ;
        RECT 296.440 44.800 296.650 45.700 ;
        RECT 294.720 44.790 294.930 44.800 ;
        RECT 291.870 44.290 292.200 44.790 ;
        RECT 292.370 44.550 294.005 44.790 ;
        RECT 292.370 44.460 292.600 44.550 ;
        RECT 292.710 44.290 293.040 44.330 ;
        RECT 291.870 44.120 293.040 44.290 ;
        RECT 293.230 43.950 293.585 44.370 ;
        RECT 293.755 44.120 294.005 44.550 ;
        RECT 294.175 43.950 294.505 44.710 ;
        RECT 294.675 44.120 294.930 44.790 ;
        RECT 295.695 44.580 296.650 44.800 ;
        RECT 296.820 45.530 297.220 46.330 ;
        RECT 297.410 45.870 297.690 46.330 ;
        RECT 298.210 46.040 298.535 46.500 ;
        RECT 297.410 45.700 298.535 45.870 ;
        RECT 298.705 45.760 299.090 46.330 ;
        RECT 298.085 45.590 298.535 45.700 ;
        RECT 296.820 44.970 297.915 45.530 ;
        RECT 298.085 45.260 298.640 45.590 ;
        RECT 295.695 44.120 295.980 44.580 ;
        RECT 296.150 43.950 296.420 44.410 ;
        RECT 296.820 44.120 297.220 44.970 ;
        RECT 298.085 44.800 298.535 45.260 ;
        RECT 298.810 45.090 299.090 45.760 ;
        RECT 300.095 45.790 300.350 46.320 ;
        RECT 300.530 46.040 300.815 46.500 ;
        RECT 300.095 45.140 300.275 45.790 ;
        RECT 300.995 45.590 301.245 46.240 ;
        RECT 300.445 45.260 301.245 45.590 ;
        RECT 297.410 44.580 298.535 44.800 ;
        RECT 297.410 44.120 297.690 44.580 ;
        RECT 298.210 43.950 298.535 44.410 ;
        RECT 298.705 44.120 299.090 45.090 ;
        RECT 300.010 44.970 300.275 45.140 ;
        RECT 300.095 44.930 300.275 44.970 ;
        RECT 300.095 44.260 300.350 44.930 ;
        RECT 300.530 43.950 300.815 44.750 ;
        RECT 300.995 44.670 301.245 45.260 ;
        RECT 301.445 45.905 301.765 46.235 ;
        RECT 301.945 46.020 302.605 46.500 ;
        RECT 302.805 46.110 303.655 46.280 ;
        RECT 301.445 45.010 301.635 45.905 ;
        RECT 301.955 45.580 302.615 45.850 ;
        RECT 302.285 45.520 302.615 45.580 ;
        RECT 301.805 45.350 302.135 45.410 ;
        RECT 302.805 45.350 302.975 46.110 ;
        RECT 304.215 46.040 304.535 46.500 ;
        RECT 304.735 45.860 304.985 46.290 ;
        RECT 305.275 46.060 305.685 46.500 ;
        RECT 305.855 46.120 306.870 46.320 ;
        RECT 303.145 45.690 304.395 45.860 ;
        RECT 303.145 45.570 303.475 45.690 ;
        RECT 301.805 45.180 303.705 45.350 ;
        RECT 301.445 44.840 303.365 45.010 ;
        RECT 301.445 44.820 301.765 44.840 ;
        RECT 300.995 44.160 301.325 44.670 ;
        RECT 301.595 44.210 301.765 44.820 ;
        RECT 303.535 44.670 303.705 45.180 ;
        RECT 303.875 45.110 304.055 45.520 ;
        RECT 304.225 44.930 304.395 45.690 ;
        RECT 301.935 43.950 302.265 44.640 ;
        RECT 302.495 44.500 303.705 44.670 ;
        RECT 303.875 44.620 304.395 44.930 ;
        RECT 304.565 45.520 304.985 45.860 ;
        RECT 305.275 45.520 305.685 45.850 ;
        RECT 304.565 44.750 304.755 45.520 ;
        RECT 305.855 45.390 306.025 46.120 ;
        RECT 307.170 45.950 307.340 46.280 ;
        RECT 307.510 46.120 307.840 46.500 ;
        RECT 306.195 45.570 306.545 45.940 ;
        RECT 305.855 45.350 306.275 45.390 ;
        RECT 304.925 45.180 306.275 45.350 ;
        RECT 304.925 45.020 305.175 45.180 ;
        RECT 305.685 44.750 305.935 45.010 ;
        RECT 304.565 44.500 305.935 44.750 ;
        RECT 302.495 44.210 302.735 44.500 ;
        RECT 303.535 44.420 303.705 44.500 ;
        RECT 302.935 43.950 303.355 44.330 ;
        RECT 303.535 44.170 304.165 44.420 ;
        RECT 304.635 43.950 304.965 44.330 ;
        RECT 305.135 44.210 305.305 44.500 ;
        RECT 306.105 44.335 306.275 45.180 ;
        RECT 306.725 45.010 306.945 45.880 ;
        RECT 307.170 45.760 307.865 45.950 ;
        RECT 306.445 44.630 306.945 45.010 ;
        RECT 307.115 44.960 307.525 45.580 ;
        RECT 307.695 44.790 307.865 45.760 ;
        RECT 307.170 44.620 307.865 44.790 ;
        RECT 305.485 43.950 305.865 44.330 ;
        RECT 306.105 44.165 306.935 44.335 ;
        RECT 307.170 44.120 307.340 44.620 ;
        RECT 307.510 43.950 307.840 44.450 ;
        RECT 308.055 44.120 308.280 46.240 ;
        RECT 308.450 46.120 308.780 46.500 ;
        RECT 308.950 45.950 309.120 46.240 ;
        RECT 308.455 45.780 309.120 45.950 ;
        RECT 308.455 44.790 308.685 45.780 ;
        RECT 309.840 45.750 311.050 46.500 ;
        RECT 308.855 44.960 309.205 45.610 ;
        RECT 309.840 45.040 310.360 45.580 ;
        RECT 310.530 45.210 311.050 45.750 ;
        RECT 308.455 44.620 309.120 44.790 ;
        RECT 308.450 43.950 308.780 44.450 ;
        RECT 308.950 44.120 309.120 44.620 ;
        RECT 309.840 43.950 311.050 45.040 ;
        RECT 162.095 43.780 311.135 43.950 ;
        RECT 162.180 42.690 163.390 43.780 ;
        RECT 163.560 43.345 168.905 43.780 ;
        RECT 162.180 41.980 162.700 42.520 ;
        RECT 162.870 42.150 163.390 42.690 ;
        RECT 162.180 41.230 163.390 41.980 ;
        RECT 165.145 41.775 165.485 42.605 ;
        RECT 166.965 42.095 167.315 43.345 ;
        RECT 170.000 42.705 170.270 43.610 ;
        RECT 170.440 43.020 170.770 43.780 ;
        RECT 170.950 42.850 171.120 43.610 ;
        RECT 171.495 43.150 171.780 43.610 ;
        RECT 171.950 43.320 172.220 43.780 ;
        RECT 171.495 42.930 172.450 43.150 ;
        RECT 170.000 41.905 170.170 42.705 ;
        RECT 170.455 42.680 171.120 42.850 ;
        RECT 170.455 42.535 170.625 42.680 ;
        RECT 170.340 42.205 170.625 42.535 ;
        RECT 170.455 41.950 170.625 42.205 ;
        RECT 170.860 42.130 171.190 42.500 ;
        RECT 171.380 42.200 172.070 42.760 ;
        RECT 172.240 42.030 172.450 42.930 ;
        RECT 163.560 41.230 168.905 41.775 ;
        RECT 170.000 41.400 170.260 41.905 ;
        RECT 170.455 41.780 171.120 41.950 ;
        RECT 170.440 41.230 170.770 41.610 ;
        RECT 170.950 41.400 171.120 41.780 ;
        RECT 171.495 41.860 172.450 42.030 ;
        RECT 172.620 42.760 173.020 43.610 ;
        RECT 173.210 43.150 173.490 43.610 ;
        RECT 174.010 43.320 174.335 43.780 ;
        RECT 173.210 42.930 174.335 43.150 ;
        RECT 172.620 42.200 173.715 42.760 ;
        RECT 173.885 42.470 174.335 42.930 ;
        RECT 174.505 42.640 174.890 43.610 ;
        RECT 171.495 41.400 171.780 41.860 ;
        RECT 171.950 41.230 172.220 41.690 ;
        RECT 172.620 41.400 173.020 42.200 ;
        RECT 173.885 42.140 174.440 42.470 ;
        RECT 173.885 42.030 174.335 42.140 ;
        RECT 173.210 41.860 174.335 42.030 ;
        RECT 174.610 41.970 174.890 42.640 ;
        RECT 175.060 42.615 175.350 43.780 ;
        RECT 175.525 42.640 175.860 43.610 ;
        RECT 176.030 42.640 176.200 43.780 ;
        RECT 176.370 43.440 178.400 43.610 ;
        RECT 173.210 41.400 173.490 41.860 ;
        RECT 174.010 41.230 174.335 41.690 ;
        RECT 174.505 41.400 174.890 41.970 ;
        RECT 175.525 41.970 175.695 42.640 ;
        RECT 176.370 42.470 176.540 43.440 ;
        RECT 175.865 42.140 176.120 42.470 ;
        RECT 176.345 42.140 176.540 42.470 ;
        RECT 176.710 43.100 177.835 43.270 ;
        RECT 175.950 41.970 176.120 42.140 ;
        RECT 176.710 41.970 176.880 43.100 ;
        RECT 175.060 41.230 175.350 41.955 ;
        RECT 175.525 41.400 175.780 41.970 ;
        RECT 175.950 41.800 176.880 41.970 ;
        RECT 177.050 42.760 178.060 42.930 ;
        RECT 177.050 41.960 177.220 42.760 ;
        RECT 177.425 42.080 177.700 42.560 ;
        RECT 177.420 41.910 177.700 42.080 ;
        RECT 176.705 41.765 176.880 41.800 ;
        RECT 175.950 41.230 176.280 41.630 ;
        RECT 176.705 41.400 177.235 41.765 ;
        RECT 177.425 41.400 177.700 41.910 ;
        RECT 177.870 41.400 178.060 42.760 ;
        RECT 178.230 42.775 178.400 43.440 ;
        RECT 178.570 43.020 178.740 43.780 ;
        RECT 178.975 43.020 179.490 43.430 ;
        RECT 178.230 42.585 178.980 42.775 ;
        RECT 179.150 42.210 179.490 43.020 ;
        RECT 178.260 42.040 179.490 42.210 ;
        RECT 180.120 42.705 180.390 43.610 ;
        RECT 180.560 43.020 180.890 43.780 ;
        RECT 181.070 42.850 181.240 43.610 ;
        RECT 178.240 41.230 178.750 41.765 ;
        RECT 178.970 41.435 179.215 42.040 ;
        RECT 180.120 41.905 180.290 42.705 ;
        RECT 180.575 42.680 181.240 42.850 ;
        RECT 180.575 42.535 180.745 42.680 ;
        RECT 180.460 42.205 180.745 42.535 ;
        RECT 181.965 42.640 182.300 43.610 ;
        RECT 182.470 42.640 182.640 43.780 ;
        RECT 182.810 43.440 184.840 43.610 ;
        RECT 180.575 41.950 180.745 42.205 ;
        RECT 180.980 42.130 181.310 42.500 ;
        RECT 181.965 41.970 182.135 42.640 ;
        RECT 182.810 42.470 182.980 43.440 ;
        RECT 182.305 42.140 182.560 42.470 ;
        RECT 182.785 42.140 182.980 42.470 ;
        RECT 183.150 43.100 184.275 43.270 ;
        RECT 182.390 41.970 182.560 42.140 ;
        RECT 183.150 41.970 183.320 43.100 ;
        RECT 180.120 41.400 180.380 41.905 ;
        RECT 180.575 41.780 181.240 41.950 ;
        RECT 180.560 41.230 180.890 41.610 ;
        RECT 181.070 41.400 181.240 41.780 ;
        RECT 181.965 41.400 182.220 41.970 ;
        RECT 182.390 41.800 183.320 41.970 ;
        RECT 183.490 42.760 184.500 42.930 ;
        RECT 183.490 41.960 183.660 42.760 ;
        RECT 183.145 41.765 183.320 41.800 ;
        RECT 182.390 41.230 182.720 41.630 ;
        RECT 183.145 41.400 183.675 41.765 ;
        RECT 183.865 41.740 184.140 42.560 ;
        RECT 183.860 41.570 184.140 41.740 ;
        RECT 183.865 41.400 184.140 41.570 ;
        RECT 184.310 41.400 184.500 42.760 ;
        RECT 184.670 42.775 184.840 43.440 ;
        RECT 185.010 43.020 185.180 43.780 ;
        RECT 185.415 43.020 185.930 43.430 ;
        RECT 184.670 42.585 185.420 42.775 ;
        RECT 185.590 42.210 185.930 43.020 ;
        RECT 186.215 43.150 186.500 43.610 ;
        RECT 186.670 43.320 186.940 43.780 ;
        RECT 186.215 42.930 187.170 43.150 ;
        RECT 184.700 42.040 185.930 42.210 ;
        RECT 186.100 42.200 186.790 42.760 ;
        RECT 184.680 41.230 185.190 41.765 ;
        RECT 185.410 41.435 185.655 42.040 ;
        RECT 186.960 42.030 187.170 42.930 ;
        RECT 186.215 41.860 187.170 42.030 ;
        RECT 187.340 42.760 187.740 43.610 ;
        RECT 187.930 43.150 188.210 43.610 ;
        RECT 188.730 43.320 189.055 43.780 ;
        RECT 187.930 42.930 189.055 43.150 ;
        RECT 187.340 42.200 188.435 42.760 ;
        RECT 188.605 42.470 189.055 42.930 ;
        RECT 189.225 42.640 189.610 43.610 ;
        RECT 190.245 43.110 190.500 43.610 ;
        RECT 190.670 43.280 191.000 43.780 ;
        RECT 190.245 42.940 190.995 43.110 ;
        RECT 186.215 41.400 186.500 41.860 ;
        RECT 186.670 41.230 186.940 41.690 ;
        RECT 187.340 41.400 187.740 42.200 ;
        RECT 188.605 42.140 189.160 42.470 ;
        RECT 188.605 42.030 189.055 42.140 ;
        RECT 187.930 41.860 189.055 42.030 ;
        RECT 189.330 41.970 189.610 42.640 ;
        RECT 190.245 42.120 190.595 42.770 ;
        RECT 187.930 41.400 188.210 41.860 ;
        RECT 188.730 41.230 189.055 41.690 ;
        RECT 189.225 41.400 189.610 41.970 ;
        RECT 190.765 41.950 190.995 42.940 ;
        RECT 190.245 41.780 190.995 41.950 ;
        RECT 190.245 41.490 190.500 41.780 ;
        RECT 190.670 41.230 191.000 41.610 ;
        RECT 191.170 41.490 191.340 43.610 ;
        RECT 191.510 42.810 191.835 43.595 ;
        RECT 192.005 43.320 192.255 43.780 ;
        RECT 192.425 43.280 192.675 43.610 ;
        RECT 192.890 43.280 193.570 43.610 ;
        RECT 192.425 43.150 192.595 43.280 ;
        RECT 192.200 42.980 192.595 43.150 ;
        RECT 191.570 41.760 192.030 42.810 ;
        RECT 192.200 41.620 192.370 42.980 ;
        RECT 192.765 42.720 193.230 43.110 ;
        RECT 192.540 41.910 192.890 42.530 ;
        RECT 193.060 42.130 193.230 42.720 ;
        RECT 193.400 42.500 193.570 43.280 ;
        RECT 193.740 43.180 193.910 43.520 ;
        RECT 194.145 43.350 194.475 43.780 ;
        RECT 194.645 43.180 194.815 43.520 ;
        RECT 195.110 43.320 195.480 43.780 ;
        RECT 193.740 43.010 194.815 43.180 ;
        RECT 195.650 43.150 195.820 43.610 ;
        RECT 196.055 43.270 196.925 43.610 ;
        RECT 197.095 43.320 197.345 43.780 ;
        RECT 195.260 42.980 195.820 43.150 ;
        RECT 195.260 42.840 195.430 42.980 ;
        RECT 193.930 42.670 195.430 42.840 ;
        RECT 196.125 42.810 196.585 43.100 ;
        RECT 193.400 42.330 195.090 42.500 ;
        RECT 193.060 41.910 193.415 42.130 ;
        RECT 193.585 41.620 193.755 42.330 ;
        RECT 193.960 41.910 194.750 42.160 ;
        RECT 194.920 42.150 195.090 42.330 ;
        RECT 195.260 41.980 195.430 42.670 ;
        RECT 191.700 41.230 192.030 41.590 ;
        RECT 192.200 41.450 192.695 41.620 ;
        RECT 192.900 41.450 193.755 41.620 ;
        RECT 194.630 41.230 194.960 41.690 ;
        RECT 195.170 41.590 195.430 41.980 ;
        RECT 195.620 42.800 196.585 42.810 ;
        RECT 196.755 42.890 196.925 43.270 ;
        RECT 197.515 43.230 197.685 43.520 ;
        RECT 197.865 43.400 198.195 43.780 ;
        RECT 197.515 43.060 198.315 43.230 ;
        RECT 195.620 42.640 196.295 42.800 ;
        RECT 196.755 42.720 197.975 42.890 ;
        RECT 195.620 41.850 195.830 42.640 ;
        RECT 196.755 42.630 196.925 42.720 ;
        RECT 196.000 41.850 196.350 42.470 ;
        RECT 196.520 42.460 196.925 42.630 ;
        RECT 196.520 41.680 196.690 42.460 ;
        RECT 196.860 42.010 197.080 42.290 ;
        RECT 197.260 42.180 197.800 42.550 ;
        RECT 198.145 42.440 198.315 43.060 ;
        RECT 198.490 42.720 198.660 43.780 ;
        RECT 198.870 42.770 199.160 43.610 ;
        RECT 199.330 42.940 199.500 43.780 ;
        RECT 199.710 42.770 199.960 43.610 ;
        RECT 200.170 42.940 200.340 43.780 ;
        RECT 198.870 42.600 200.595 42.770 ;
        RECT 200.820 42.615 201.110 43.780 ;
        RECT 201.285 43.110 201.540 43.610 ;
        RECT 201.710 43.280 202.040 43.780 ;
        RECT 201.285 42.940 202.035 43.110 ;
        RECT 196.860 41.840 197.390 42.010 ;
        RECT 195.170 41.420 195.520 41.590 ;
        RECT 195.740 41.400 196.690 41.680 ;
        RECT 196.860 41.230 197.050 41.670 ;
        RECT 197.220 41.610 197.390 41.840 ;
        RECT 197.560 41.780 197.800 42.180 ;
        RECT 197.970 42.430 198.315 42.440 ;
        RECT 197.970 42.220 200.000 42.430 ;
        RECT 197.970 41.965 198.295 42.220 ;
        RECT 200.185 42.050 200.595 42.600 ;
        RECT 201.285 42.120 201.635 42.770 ;
        RECT 197.970 41.610 198.290 41.965 ;
        RECT 197.220 41.440 198.290 41.610 ;
        RECT 198.490 41.230 198.660 42.040 ;
        RECT 198.830 41.880 200.595 42.050 ;
        RECT 198.830 41.400 199.160 41.880 ;
        RECT 199.330 41.230 199.500 41.700 ;
        RECT 199.670 41.400 200.000 41.880 ;
        RECT 200.170 41.230 200.340 41.700 ;
        RECT 200.820 41.230 201.110 41.955 ;
        RECT 201.805 41.950 202.035 42.940 ;
        RECT 201.285 41.780 202.035 41.950 ;
        RECT 201.285 41.490 201.540 41.780 ;
        RECT 201.710 41.230 202.040 41.610 ;
        RECT 202.210 41.490 202.380 43.610 ;
        RECT 202.550 42.810 202.875 43.595 ;
        RECT 203.045 43.320 203.295 43.780 ;
        RECT 203.465 43.280 203.715 43.610 ;
        RECT 203.930 43.280 204.610 43.610 ;
        RECT 203.465 43.150 203.635 43.280 ;
        RECT 203.240 42.980 203.635 43.150 ;
        RECT 202.610 41.760 203.070 42.810 ;
        RECT 203.240 41.620 203.410 42.980 ;
        RECT 203.805 42.720 204.270 43.110 ;
        RECT 203.580 41.910 203.930 42.530 ;
        RECT 204.100 42.130 204.270 42.720 ;
        RECT 204.440 42.500 204.610 43.280 ;
        RECT 204.780 43.180 204.950 43.520 ;
        RECT 205.185 43.350 205.515 43.780 ;
        RECT 205.685 43.180 205.855 43.520 ;
        RECT 206.150 43.320 206.520 43.780 ;
        RECT 204.780 43.010 205.855 43.180 ;
        RECT 206.690 43.150 206.860 43.610 ;
        RECT 207.095 43.270 207.965 43.610 ;
        RECT 208.135 43.320 208.385 43.780 ;
        RECT 206.300 42.980 206.860 43.150 ;
        RECT 206.300 42.840 206.470 42.980 ;
        RECT 204.970 42.670 206.470 42.840 ;
        RECT 207.165 42.810 207.625 43.100 ;
        RECT 204.440 42.330 206.130 42.500 ;
        RECT 204.100 41.910 204.455 42.130 ;
        RECT 204.625 41.620 204.795 42.330 ;
        RECT 205.000 41.910 205.790 42.160 ;
        RECT 205.960 42.150 206.130 42.330 ;
        RECT 206.300 41.980 206.470 42.670 ;
        RECT 202.740 41.230 203.070 41.590 ;
        RECT 203.240 41.450 203.735 41.620 ;
        RECT 203.940 41.450 204.795 41.620 ;
        RECT 205.670 41.230 206.000 41.690 ;
        RECT 206.210 41.590 206.470 41.980 ;
        RECT 206.660 42.800 207.625 42.810 ;
        RECT 207.795 42.890 207.965 43.270 ;
        RECT 208.555 43.230 208.725 43.520 ;
        RECT 208.905 43.400 209.235 43.780 ;
        RECT 208.555 43.060 209.355 43.230 ;
        RECT 206.660 42.640 207.335 42.800 ;
        RECT 207.795 42.720 209.015 42.890 ;
        RECT 206.660 41.850 206.870 42.640 ;
        RECT 207.795 42.630 207.965 42.720 ;
        RECT 207.040 41.850 207.390 42.470 ;
        RECT 207.560 42.460 207.965 42.630 ;
        RECT 207.560 41.680 207.730 42.460 ;
        RECT 207.900 42.010 208.120 42.290 ;
        RECT 208.300 42.180 208.840 42.550 ;
        RECT 209.185 42.440 209.355 43.060 ;
        RECT 209.530 42.720 209.700 43.780 ;
        RECT 209.910 42.770 210.200 43.610 ;
        RECT 210.370 42.940 210.540 43.780 ;
        RECT 210.750 42.770 211.000 43.610 ;
        RECT 211.210 42.940 211.380 43.780 ;
        RECT 211.950 43.160 212.120 43.590 ;
        RECT 212.290 43.330 212.620 43.780 ;
        RECT 211.950 42.930 212.625 43.160 ;
        RECT 209.910 42.600 211.635 42.770 ;
        RECT 207.900 41.840 208.430 42.010 ;
        RECT 206.210 41.420 206.560 41.590 ;
        RECT 206.780 41.400 207.730 41.680 ;
        RECT 207.900 41.230 208.090 41.670 ;
        RECT 208.260 41.610 208.430 41.840 ;
        RECT 208.600 41.780 208.840 42.180 ;
        RECT 209.010 42.430 209.355 42.440 ;
        RECT 209.010 42.220 211.040 42.430 ;
        RECT 209.010 41.965 209.335 42.220 ;
        RECT 211.225 42.050 211.635 42.600 ;
        RECT 209.010 41.610 209.330 41.965 ;
        RECT 208.260 41.440 209.330 41.610 ;
        RECT 209.530 41.230 209.700 42.040 ;
        RECT 209.870 41.880 211.635 42.050 ;
        RECT 211.920 41.910 212.220 42.760 ;
        RECT 212.390 42.280 212.625 42.930 ;
        RECT 212.795 42.620 213.080 43.565 ;
        RECT 213.260 43.310 213.945 43.780 ;
        RECT 213.255 42.790 213.950 43.100 ;
        RECT 214.125 42.725 214.430 43.510 ;
        RECT 212.795 42.470 213.655 42.620 ;
        RECT 212.795 42.450 214.080 42.470 ;
        RECT 212.390 41.950 212.925 42.280 ;
        RECT 213.095 42.090 214.080 42.450 ;
        RECT 209.870 41.400 210.200 41.880 ;
        RECT 210.370 41.230 210.540 41.700 ;
        RECT 210.710 41.400 211.040 41.880 ;
        RECT 212.390 41.800 212.610 41.950 ;
        RECT 211.210 41.230 211.380 41.700 ;
        RECT 211.865 41.230 212.200 41.735 ;
        RECT 212.370 41.425 212.610 41.800 ;
        RECT 213.095 41.755 213.265 42.090 ;
        RECT 214.255 41.920 214.430 42.725 ;
        RECT 212.890 41.560 213.265 41.755 ;
        RECT 212.890 41.415 213.060 41.560 ;
        RECT 213.625 41.230 214.020 41.725 ;
        RECT 214.190 41.400 214.430 41.920 ;
        RECT 214.620 42.810 214.930 43.610 ;
        RECT 215.100 42.980 215.410 43.780 ;
        RECT 215.580 43.150 215.840 43.610 ;
        RECT 216.010 43.320 216.265 43.780 ;
        RECT 216.440 43.150 216.700 43.610 ;
        RECT 215.580 42.980 216.700 43.150 ;
        RECT 214.620 42.640 215.650 42.810 ;
        RECT 214.620 41.730 214.790 42.640 ;
        RECT 214.960 41.900 215.310 42.470 ;
        RECT 215.480 42.390 215.650 42.640 ;
        RECT 216.440 42.730 216.700 42.980 ;
        RECT 216.870 42.910 217.155 43.780 ;
        RECT 217.385 43.110 217.640 43.610 ;
        RECT 217.810 43.280 218.140 43.780 ;
        RECT 217.385 42.940 218.135 43.110 ;
        RECT 216.440 42.560 217.195 42.730 ;
        RECT 215.480 42.220 216.620 42.390 ;
        RECT 216.790 42.050 217.195 42.560 ;
        RECT 217.385 42.120 217.735 42.770 ;
        RECT 215.545 41.880 217.195 42.050 ;
        RECT 217.905 41.950 218.135 42.940 ;
        RECT 214.620 41.400 214.920 41.730 ;
        RECT 215.090 41.230 215.365 41.710 ;
        RECT 215.545 41.490 215.840 41.880 ;
        RECT 216.010 41.230 216.265 41.710 ;
        RECT 216.440 41.490 216.700 41.880 ;
        RECT 217.385 41.780 218.135 41.950 ;
        RECT 216.870 41.230 217.150 41.710 ;
        RECT 217.385 41.490 217.640 41.780 ;
        RECT 217.810 41.230 218.140 41.610 ;
        RECT 218.310 41.490 218.480 43.610 ;
        RECT 218.650 42.810 218.975 43.595 ;
        RECT 219.145 43.320 219.395 43.780 ;
        RECT 219.565 43.280 219.815 43.610 ;
        RECT 220.030 43.280 220.710 43.610 ;
        RECT 219.565 43.150 219.735 43.280 ;
        RECT 219.340 42.980 219.735 43.150 ;
        RECT 218.710 41.760 219.170 42.810 ;
        RECT 219.340 41.620 219.510 42.980 ;
        RECT 219.905 42.720 220.370 43.110 ;
        RECT 219.680 41.910 220.030 42.530 ;
        RECT 220.200 42.130 220.370 42.720 ;
        RECT 220.540 42.500 220.710 43.280 ;
        RECT 220.880 43.180 221.050 43.520 ;
        RECT 221.285 43.350 221.615 43.780 ;
        RECT 221.785 43.180 221.955 43.520 ;
        RECT 222.250 43.320 222.620 43.780 ;
        RECT 220.880 43.010 221.955 43.180 ;
        RECT 222.790 43.150 222.960 43.610 ;
        RECT 223.195 43.270 224.065 43.610 ;
        RECT 224.235 43.320 224.485 43.780 ;
        RECT 222.400 42.980 222.960 43.150 ;
        RECT 222.400 42.840 222.570 42.980 ;
        RECT 221.070 42.670 222.570 42.840 ;
        RECT 223.265 42.810 223.725 43.100 ;
        RECT 220.540 42.330 222.230 42.500 ;
        RECT 220.200 41.910 220.555 42.130 ;
        RECT 220.725 41.620 220.895 42.330 ;
        RECT 221.100 41.910 221.890 42.160 ;
        RECT 222.060 42.150 222.230 42.330 ;
        RECT 222.400 41.980 222.570 42.670 ;
        RECT 218.840 41.230 219.170 41.590 ;
        RECT 219.340 41.450 219.835 41.620 ;
        RECT 220.040 41.450 220.895 41.620 ;
        RECT 221.770 41.230 222.100 41.690 ;
        RECT 222.310 41.590 222.570 41.980 ;
        RECT 222.760 42.800 223.725 42.810 ;
        RECT 223.895 42.890 224.065 43.270 ;
        RECT 224.655 43.230 224.825 43.520 ;
        RECT 225.005 43.400 225.335 43.780 ;
        RECT 224.655 43.060 225.455 43.230 ;
        RECT 222.760 42.640 223.435 42.800 ;
        RECT 223.895 42.720 225.115 42.890 ;
        RECT 222.760 41.850 222.970 42.640 ;
        RECT 223.895 42.630 224.065 42.720 ;
        RECT 223.140 41.850 223.490 42.470 ;
        RECT 223.660 42.460 224.065 42.630 ;
        RECT 223.660 41.680 223.830 42.460 ;
        RECT 224.000 42.010 224.220 42.290 ;
        RECT 224.400 42.180 224.940 42.550 ;
        RECT 225.285 42.470 225.455 43.060 ;
        RECT 225.675 42.640 225.980 43.780 ;
        RECT 226.150 42.590 226.405 43.470 ;
        RECT 226.580 42.615 226.870 43.780 ;
        RECT 227.350 42.940 227.520 43.780 ;
        RECT 227.730 42.770 227.980 43.610 ;
        RECT 228.190 42.940 228.360 43.780 ;
        RECT 228.530 42.770 228.820 43.610 ;
        RECT 225.285 42.440 226.025 42.470 ;
        RECT 224.000 41.840 224.530 42.010 ;
        RECT 222.310 41.420 222.660 41.590 ;
        RECT 222.880 41.400 223.830 41.680 ;
        RECT 224.000 41.230 224.190 41.670 ;
        RECT 224.360 41.610 224.530 41.840 ;
        RECT 224.700 41.780 224.940 42.180 ;
        RECT 225.110 42.140 226.025 42.440 ;
        RECT 225.110 41.965 225.435 42.140 ;
        RECT 225.110 41.610 225.430 41.965 ;
        RECT 226.195 41.940 226.405 42.590 ;
        RECT 227.095 42.600 228.820 42.770 ;
        RECT 229.030 42.720 229.200 43.780 ;
        RECT 229.495 43.400 229.825 43.780 ;
        RECT 230.005 43.230 230.175 43.520 ;
        RECT 230.345 43.320 230.595 43.780 ;
        RECT 229.375 43.060 230.175 43.230 ;
        RECT 230.765 43.270 231.635 43.610 ;
        RECT 227.095 42.050 227.505 42.600 ;
        RECT 229.375 42.440 229.545 43.060 ;
        RECT 230.765 42.890 230.935 43.270 ;
        RECT 231.870 43.150 232.040 43.610 ;
        RECT 232.210 43.320 232.580 43.780 ;
        RECT 232.875 43.180 233.045 43.520 ;
        RECT 233.215 43.350 233.545 43.780 ;
        RECT 233.780 43.180 233.950 43.520 ;
        RECT 229.715 42.720 230.935 42.890 ;
        RECT 231.105 42.810 231.565 43.100 ;
        RECT 231.870 42.980 232.430 43.150 ;
        RECT 232.875 43.010 233.950 43.180 ;
        RECT 234.120 43.280 234.800 43.610 ;
        RECT 235.015 43.280 235.265 43.610 ;
        RECT 235.435 43.320 235.685 43.780 ;
        RECT 232.260 42.840 232.430 42.980 ;
        RECT 231.105 42.800 232.070 42.810 ;
        RECT 230.765 42.630 230.935 42.720 ;
        RECT 231.395 42.640 232.070 42.800 ;
        RECT 229.375 42.430 229.720 42.440 ;
        RECT 227.690 42.220 229.720 42.430 ;
        RECT 224.360 41.440 225.430 41.610 ;
        RECT 225.675 41.230 225.980 41.690 ;
        RECT 226.150 41.410 226.405 41.940 ;
        RECT 226.580 41.230 226.870 41.955 ;
        RECT 227.095 41.880 228.860 42.050 ;
        RECT 227.350 41.230 227.520 41.700 ;
        RECT 227.690 41.400 228.020 41.880 ;
        RECT 228.190 41.230 228.360 41.700 ;
        RECT 228.530 41.400 228.860 41.880 ;
        RECT 229.030 41.230 229.200 42.040 ;
        RECT 229.395 41.965 229.720 42.220 ;
        RECT 229.400 41.610 229.720 41.965 ;
        RECT 229.890 42.180 230.430 42.550 ;
        RECT 230.765 42.460 231.170 42.630 ;
        RECT 229.890 41.780 230.130 42.180 ;
        RECT 230.610 42.010 230.830 42.290 ;
        RECT 230.300 41.840 230.830 42.010 ;
        RECT 230.300 41.610 230.470 41.840 ;
        RECT 231.000 41.680 231.170 42.460 ;
        RECT 231.340 41.850 231.690 42.470 ;
        RECT 231.860 41.850 232.070 42.640 ;
        RECT 232.260 42.670 233.760 42.840 ;
        RECT 232.260 41.980 232.430 42.670 ;
        RECT 234.120 42.500 234.290 43.280 ;
        RECT 235.095 43.150 235.265 43.280 ;
        RECT 232.600 42.330 234.290 42.500 ;
        RECT 234.460 42.720 234.925 43.110 ;
        RECT 235.095 42.980 235.490 43.150 ;
        RECT 232.600 42.150 232.770 42.330 ;
        RECT 229.400 41.440 230.470 41.610 ;
        RECT 230.640 41.230 230.830 41.670 ;
        RECT 231.000 41.400 231.950 41.680 ;
        RECT 232.260 41.590 232.520 41.980 ;
        RECT 232.940 41.910 233.730 42.160 ;
        RECT 232.170 41.420 232.520 41.590 ;
        RECT 232.730 41.230 233.060 41.690 ;
        RECT 233.935 41.620 234.105 42.330 ;
        RECT 234.460 42.130 234.630 42.720 ;
        RECT 234.275 41.910 234.630 42.130 ;
        RECT 234.800 41.910 235.150 42.530 ;
        RECT 235.320 41.620 235.490 42.980 ;
        RECT 235.855 42.810 236.180 43.595 ;
        RECT 235.660 41.760 236.120 42.810 ;
        RECT 233.935 41.450 234.790 41.620 ;
        RECT 234.995 41.450 235.490 41.620 ;
        RECT 235.660 41.230 235.990 41.590 ;
        RECT 236.350 41.490 236.520 43.610 ;
        RECT 236.690 43.280 237.020 43.780 ;
        RECT 237.190 43.110 237.445 43.610 ;
        RECT 236.695 42.940 237.445 43.110 ;
        RECT 236.695 41.950 236.925 42.940 ;
        RECT 237.095 42.120 237.445 42.770 ;
        RECT 237.620 42.640 238.005 43.610 ;
        RECT 238.175 43.320 238.500 43.780 ;
        RECT 239.020 43.150 239.300 43.610 ;
        RECT 238.175 42.930 239.300 43.150 ;
        RECT 237.620 41.970 237.900 42.640 ;
        RECT 238.175 42.470 238.625 42.930 ;
        RECT 239.490 42.760 239.890 43.610 ;
        RECT 240.290 43.320 240.560 43.780 ;
        RECT 240.730 43.150 241.015 43.610 ;
        RECT 238.070 42.140 238.625 42.470 ;
        RECT 238.795 42.200 239.890 42.760 ;
        RECT 238.175 42.030 238.625 42.140 ;
        RECT 236.695 41.780 237.445 41.950 ;
        RECT 236.690 41.230 237.020 41.610 ;
        RECT 237.190 41.490 237.445 41.780 ;
        RECT 237.620 41.400 238.005 41.970 ;
        RECT 238.175 41.860 239.300 42.030 ;
        RECT 238.175 41.230 238.500 41.690 ;
        RECT 239.020 41.400 239.300 41.860 ;
        RECT 239.490 41.400 239.890 42.200 ;
        RECT 240.060 42.930 241.015 43.150 ;
        RECT 240.060 42.030 240.270 42.930 ;
        RECT 240.440 42.200 241.130 42.760 ;
        RECT 241.300 42.690 242.970 43.780 ;
        RECT 240.060 41.860 241.015 42.030 ;
        RECT 240.290 41.230 240.560 41.690 ;
        RECT 240.730 41.400 241.015 41.860 ;
        RECT 241.300 42.000 242.050 42.520 ;
        RECT 242.220 42.170 242.970 42.690 ;
        RECT 243.600 42.640 243.985 43.610 ;
        RECT 244.155 43.320 244.480 43.780 ;
        RECT 245.000 43.150 245.280 43.610 ;
        RECT 244.155 42.930 245.280 43.150 ;
        RECT 241.300 41.230 242.970 42.000 ;
        RECT 243.600 41.970 243.880 42.640 ;
        RECT 244.155 42.470 244.605 42.930 ;
        RECT 245.470 42.760 245.870 43.610 ;
        RECT 246.270 43.320 246.540 43.780 ;
        RECT 246.710 43.150 246.995 43.610 ;
        RECT 244.050 42.140 244.605 42.470 ;
        RECT 244.775 42.200 245.870 42.760 ;
        RECT 244.155 42.030 244.605 42.140 ;
        RECT 243.600 41.400 243.985 41.970 ;
        RECT 244.155 41.860 245.280 42.030 ;
        RECT 244.155 41.230 244.480 41.690 ;
        RECT 245.000 41.400 245.280 41.860 ;
        RECT 245.470 41.400 245.870 42.200 ;
        RECT 246.040 42.930 246.995 43.150 ;
        RECT 246.040 42.030 246.250 42.930 ;
        RECT 246.420 42.200 247.110 42.760 ;
        RECT 247.280 42.690 250.790 43.780 ;
        RECT 250.960 42.690 252.170 43.780 ;
        RECT 246.040 41.860 246.995 42.030 ;
        RECT 246.270 41.230 246.540 41.690 ;
        RECT 246.710 41.400 246.995 41.860 ;
        RECT 247.280 42.000 248.930 42.520 ;
        RECT 249.100 42.170 250.790 42.690 ;
        RECT 247.280 41.230 250.790 42.000 ;
        RECT 250.960 41.980 251.480 42.520 ;
        RECT 251.650 42.150 252.170 42.690 ;
        RECT 252.340 42.615 252.630 43.780 ;
        RECT 252.800 42.930 253.060 43.610 ;
        RECT 253.230 43.000 253.480 43.780 ;
        RECT 253.730 43.230 253.980 43.610 ;
        RECT 254.150 43.400 254.505 43.780 ;
        RECT 255.510 43.390 255.845 43.610 ;
        RECT 255.110 43.230 255.340 43.270 ;
        RECT 253.730 43.030 255.340 43.230 ;
        RECT 253.730 43.020 254.565 43.030 ;
        RECT 255.155 42.940 255.340 43.030 ;
        RECT 250.960 41.230 252.170 41.980 ;
        RECT 252.340 41.230 252.630 41.955 ;
        RECT 252.800 41.740 252.970 42.930 ;
        RECT 254.670 42.830 255.000 42.860 ;
        RECT 253.200 42.770 255.000 42.830 ;
        RECT 255.590 42.770 255.845 43.390 ;
        RECT 253.140 42.660 255.845 42.770 ;
        RECT 253.140 42.625 253.340 42.660 ;
        RECT 253.140 42.050 253.310 42.625 ;
        RECT 254.670 42.600 255.845 42.660 ;
        RECT 256.570 42.770 256.740 43.610 ;
        RECT 256.910 43.440 258.080 43.610 ;
        RECT 256.910 42.940 257.240 43.440 ;
        RECT 257.750 43.400 258.080 43.440 ;
        RECT 258.270 43.360 258.625 43.780 ;
        RECT 257.410 43.180 257.640 43.270 ;
        RECT 258.795 43.180 259.045 43.610 ;
        RECT 257.410 42.940 259.045 43.180 ;
        RECT 259.215 43.020 259.545 43.780 ;
        RECT 259.715 42.940 259.970 43.610 ;
        RECT 261.085 43.110 261.340 43.610 ;
        RECT 261.510 43.280 261.840 43.780 ;
        RECT 261.085 42.940 261.835 43.110 ;
        RECT 256.570 42.600 259.630 42.770 ;
        RECT 253.540 42.185 253.950 42.490 ;
        RECT 254.120 42.220 254.450 42.430 ;
        RECT 253.140 41.930 253.410 42.050 ;
        RECT 253.140 41.885 253.985 41.930 ;
        RECT 253.230 41.760 253.985 41.885 ;
        RECT 254.240 41.820 254.450 42.220 ;
        RECT 254.695 42.220 255.170 42.430 ;
        RECT 255.360 42.220 255.850 42.420 ;
        RECT 256.485 42.220 256.835 42.430 ;
        RECT 257.005 42.220 257.450 42.420 ;
        RECT 257.620 42.220 258.095 42.420 ;
        RECT 254.695 41.820 254.915 42.220 ;
        RECT 252.800 41.730 253.030 41.740 ;
        RECT 252.800 41.400 253.060 41.730 ;
        RECT 253.815 41.610 253.985 41.760 ;
        RECT 253.230 41.230 253.560 41.590 ;
        RECT 253.815 41.400 255.115 41.610 ;
        RECT 255.390 41.230 255.845 41.995 ;
        RECT 256.570 41.880 257.635 42.050 ;
        RECT 256.570 41.400 256.740 41.880 ;
        RECT 256.910 41.230 257.240 41.710 ;
        RECT 257.465 41.650 257.635 41.880 ;
        RECT 257.815 41.820 258.095 42.220 ;
        RECT 258.365 42.220 258.695 42.420 ;
        RECT 258.865 42.220 259.230 42.420 ;
        RECT 258.365 41.820 258.650 42.220 ;
        RECT 259.460 42.050 259.630 42.600 ;
        RECT 258.830 41.880 259.630 42.050 ;
        RECT 258.830 41.650 259.000 41.880 ;
        RECT 259.800 41.810 259.970 42.940 ;
        RECT 261.085 42.120 261.435 42.770 ;
        RECT 261.605 41.950 261.835 42.940 ;
        RECT 259.785 41.740 259.970 41.810 ;
        RECT 259.760 41.730 259.970 41.740 ;
        RECT 257.465 41.400 259.000 41.650 ;
        RECT 259.170 41.230 259.500 41.710 ;
        RECT 259.715 41.400 259.970 41.730 ;
        RECT 261.085 41.780 261.835 41.950 ;
        RECT 261.085 41.490 261.340 41.780 ;
        RECT 261.510 41.230 261.840 41.610 ;
        RECT 262.010 41.490 262.180 43.610 ;
        RECT 262.350 42.810 262.675 43.595 ;
        RECT 262.845 43.320 263.095 43.780 ;
        RECT 263.265 43.280 263.515 43.610 ;
        RECT 263.730 43.280 264.410 43.610 ;
        RECT 263.265 43.150 263.435 43.280 ;
        RECT 263.040 42.980 263.435 43.150 ;
        RECT 262.410 41.760 262.870 42.810 ;
        RECT 263.040 41.620 263.210 42.980 ;
        RECT 263.605 42.720 264.070 43.110 ;
        RECT 263.380 41.910 263.730 42.530 ;
        RECT 263.900 42.130 264.070 42.720 ;
        RECT 264.240 42.500 264.410 43.280 ;
        RECT 264.580 43.180 264.750 43.520 ;
        RECT 264.985 43.350 265.315 43.780 ;
        RECT 265.485 43.180 265.655 43.520 ;
        RECT 265.950 43.320 266.320 43.780 ;
        RECT 264.580 43.010 265.655 43.180 ;
        RECT 266.490 43.150 266.660 43.610 ;
        RECT 266.895 43.270 267.765 43.610 ;
        RECT 267.935 43.320 268.185 43.780 ;
        RECT 266.100 42.980 266.660 43.150 ;
        RECT 266.100 42.840 266.270 42.980 ;
        RECT 264.770 42.670 266.270 42.840 ;
        RECT 266.965 42.810 267.425 43.100 ;
        RECT 264.240 42.330 265.930 42.500 ;
        RECT 263.900 41.910 264.255 42.130 ;
        RECT 264.425 41.620 264.595 42.330 ;
        RECT 264.800 41.910 265.590 42.160 ;
        RECT 265.760 42.150 265.930 42.330 ;
        RECT 266.100 41.980 266.270 42.670 ;
        RECT 262.540 41.230 262.870 41.590 ;
        RECT 263.040 41.450 263.535 41.620 ;
        RECT 263.740 41.450 264.595 41.620 ;
        RECT 265.470 41.230 265.800 41.690 ;
        RECT 266.010 41.590 266.270 41.980 ;
        RECT 266.460 42.800 267.425 42.810 ;
        RECT 267.595 42.890 267.765 43.270 ;
        RECT 268.355 43.230 268.525 43.520 ;
        RECT 268.705 43.400 269.035 43.780 ;
        RECT 268.355 43.060 269.155 43.230 ;
        RECT 266.460 42.640 267.135 42.800 ;
        RECT 267.595 42.720 268.815 42.890 ;
        RECT 266.460 41.850 266.670 42.640 ;
        RECT 267.595 42.630 267.765 42.720 ;
        RECT 266.840 41.850 267.190 42.470 ;
        RECT 267.360 42.460 267.765 42.630 ;
        RECT 267.360 41.680 267.530 42.460 ;
        RECT 267.700 42.010 267.920 42.290 ;
        RECT 268.100 42.180 268.640 42.550 ;
        RECT 268.985 42.470 269.155 43.060 ;
        RECT 269.375 42.640 269.680 43.780 ;
        RECT 269.850 42.590 270.105 43.470 ;
        RECT 268.985 42.440 269.725 42.470 ;
        RECT 267.700 41.840 268.230 42.010 ;
        RECT 266.010 41.420 266.360 41.590 ;
        RECT 266.580 41.400 267.530 41.680 ;
        RECT 267.700 41.230 267.890 41.670 ;
        RECT 268.060 41.610 268.230 41.840 ;
        RECT 268.400 41.780 268.640 42.180 ;
        RECT 268.810 42.140 269.725 42.440 ;
        RECT 268.810 41.965 269.135 42.140 ;
        RECT 268.810 41.610 269.130 41.965 ;
        RECT 269.895 41.940 270.105 42.590 ;
        RECT 268.060 41.440 269.130 41.610 ;
        RECT 269.375 41.230 269.680 41.690 ;
        RECT 269.850 41.410 270.105 41.940 ;
        RECT 270.280 42.640 270.665 43.610 ;
        RECT 270.835 43.320 271.160 43.780 ;
        RECT 271.680 43.150 271.960 43.610 ;
        RECT 270.835 42.930 271.960 43.150 ;
        RECT 270.280 41.970 270.560 42.640 ;
        RECT 270.835 42.470 271.285 42.930 ;
        RECT 272.150 42.760 272.550 43.610 ;
        RECT 272.950 43.320 273.220 43.780 ;
        RECT 273.390 43.150 273.675 43.610 ;
        RECT 270.730 42.140 271.285 42.470 ;
        RECT 271.455 42.200 272.550 42.760 ;
        RECT 270.835 42.030 271.285 42.140 ;
        RECT 270.280 41.400 270.665 41.970 ;
        RECT 270.835 41.860 271.960 42.030 ;
        RECT 270.835 41.230 271.160 41.690 ;
        RECT 271.680 41.400 271.960 41.860 ;
        RECT 272.150 41.400 272.550 42.200 ;
        RECT 272.720 42.930 273.675 43.150 ;
        RECT 274.075 43.150 274.360 43.610 ;
        RECT 274.530 43.320 274.800 43.780 ;
        RECT 274.075 42.930 275.030 43.150 ;
        RECT 272.720 42.030 272.930 42.930 ;
        RECT 273.100 42.200 273.790 42.760 ;
        RECT 273.960 42.200 274.650 42.760 ;
        RECT 274.820 42.030 275.030 42.930 ;
        RECT 272.720 41.860 273.675 42.030 ;
        RECT 272.950 41.230 273.220 41.690 ;
        RECT 273.390 41.400 273.675 41.860 ;
        RECT 274.075 41.860 275.030 42.030 ;
        RECT 275.200 42.760 275.600 43.610 ;
        RECT 275.790 43.150 276.070 43.610 ;
        RECT 276.590 43.320 276.915 43.780 ;
        RECT 275.790 42.930 276.915 43.150 ;
        RECT 275.200 42.200 276.295 42.760 ;
        RECT 276.465 42.470 276.915 42.930 ;
        RECT 277.085 42.640 277.470 43.610 ;
        RECT 274.075 41.400 274.360 41.860 ;
        RECT 274.530 41.230 274.800 41.690 ;
        RECT 275.200 41.400 275.600 42.200 ;
        RECT 276.465 42.140 277.020 42.470 ;
        RECT 276.465 42.030 276.915 42.140 ;
        RECT 275.790 41.860 276.915 42.030 ;
        RECT 277.190 41.970 277.470 42.640 ;
        RECT 278.100 42.615 278.390 43.780 ;
        RECT 278.650 42.770 278.820 43.610 ;
        RECT 278.990 43.440 280.160 43.610 ;
        RECT 278.990 42.940 279.320 43.440 ;
        RECT 279.830 43.400 280.160 43.440 ;
        RECT 280.350 43.360 280.705 43.780 ;
        RECT 279.490 43.180 279.720 43.270 ;
        RECT 280.875 43.180 281.125 43.610 ;
        RECT 279.490 42.940 281.125 43.180 ;
        RECT 281.295 43.020 281.625 43.780 ;
        RECT 281.795 42.940 282.050 43.610 ;
        RECT 278.650 42.600 281.710 42.770 ;
        RECT 278.565 42.220 278.915 42.430 ;
        RECT 279.085 42.220 279.530 42.420 ;
        RECT 279.700 42.220 280.175 42.420 ;
        RECT 275.790 41.400 276.070 41.860 ;
        RECT 276.590 41.230 276.915 41.690 ;
        RECT 277.085 41.400 277.470 41.970 ;
        RECT 278.100 41.230 278.390 41.955 ;
        RECT 278.650 41.880 279.715 42.050 ;
        RECT 278.650 41.400 278.820 41.880 ;
        RECT 278.990 41.230 279.320 41.710 ;
        RECT 279.545 41.650 279.715 41.880 ;
        RECT 279.895 41.820 280.175 42.220 ;
        RECT 280.445 42.220 280.775 42.420 ;
        RECT 280.945 42.220 281.310 42.420 ;
        RECT 280.445 41.820 280.730 42.220 ;
        RECT 281.540 42.050 281.710 42.600 ;
        RECT 280.910 41.880 281.710 42.050 ;
        RECT 280.910 41.650 281.080 41.880 ;
        RECT 281.880 41.810 282.050 42.940 ;
        RECT 281.865 41.740 282.050 41.810 ;
        RECT 281.840 41.730 282.050 41.740 ;
        RECT 279.545 41.400 281.080 41.650 ;
        RECT 281.250 41.230 281.580 41.710 ;
        RECT 281.795 41.400 282.050 41.730 ;
        RECT 282.240 42.640 282.625 43.610 ;
        RECT 282.795 43.320 283.120 43.780 ;
        RECT 283.640 43.150 283.920 43.610 ;
        RECT 282.795 42.930 283.920 43.150 ;
        RECT 282.240 41.970 282.520 42.640 ;
        RECT 282.795 42.470 283.245 42.930 ;
        RECT 284.110 42.760 284.510 43.610 ;
        RECT 284.910 43.320 285.180 43.780 ;
        RECT 285.350 43.150 285.635 43.610 ;
        RECT 282.690 42.140 283.245 42.470 ;
        RECT 283.415 42.200 284.510 42.760 ;
        RECT 282.795 42.030 283.245 42.140 ;
        RECT 282.240 41.400 282.625 41.970 ;
        RECT 282.795 41.860 283.920 42.030 ;
        RECT 282.795 41.230 283.120 41.690 ;
        RECT 283.640 41.400 283.920 41.860 ;
        RECT 284.110 41.400 284.510 42.200 ;
        RECT 284.680 42.930 285.635 43.150 ;
        RECT 286.035 43.150 286.320 43.610 ;
        RECT 286.490 43.320 286.760 43.780 ;
        RECT 286.035 42.930 286.990 43.150 ;
        RECT 284.680 42.030 284.890 42.930 ;
        RECT 285.060 42.200 285.750 42.760 ;
        RECT 285.920 42.200 286.610 42.760 ;
        RECT 286.780 42.030 286.990 42.930 ;
        RECT 284.680 41.860 285.635 42.030 ;
        RECT 284.910 41.230 285.180 41.690 ;
        RECT 285.350 41.400 285.635 41.860 ;
        RECT 286.035 41.860 286.990 42.030 ;
        RECT 287.160 42.760 287.560 43.610 ;
        RECT 287.750 43.150 288.030 43.610 ;
        RECT 288.550 43.320 288.875 43.780 ;
        RECT 287.750 42.930 288.875 43.150 ;
        RECT 287.160 42.200 288.255 42.760 ;
        RECT 288.425 42.470 288.875 42.930 ;
        RECT 289.045 42.640 289.430 43.610 ;
        RECT 290.575 42.910 290.860 43.780 ;
        RECT 291.030 43.150 291.290 43.610 ;
        RECT 291.465 43.320 291.720 43.780 ;
        RECT 291.890 43.150 292.150 43.610 ;
        RECT 291.030 42.980 292.150 43.150 ;
        RECT 292.320 42.980 292.630 43.780 ;
        RECT 291.030 42.730 291.290 42.980 ;
        RECT 292.800 42.810 293.110 43.610 ;
        RECT 286.035 41.400 286.320 41.860 ;
        RECT 286.490 41.230 286.760 41.690 ;
        RECT 287.160 41.400 287.560 42.200 ;
        RECT 288.425 42.140 288.980 42.470 ;
        RECT 288.425 42.030 288.875 42.140 ;
        RECT 287.750 41.860 288.875 42.030 ;
        RECT 289.150 41.970 289.430 42.640 ;
        RECT 287.750 41.400 288.030 41.860 ;
        RECT 288.550 41.230 288.875 41.690 ;
        RECT 289.045 41.400 289.430 41.970 ;
        RECT 290.535 42.560 291.290 42.730 ;
        RECT 292.080 42.640 293.110 42.810 ;
        RECT 293.280 42.690 294.950 43.780 ;
        RECT 295.175 42.910 295.460 43.780 ;
        RECT 295.630 43.150 295.890 43.610 ;
        RECT 296.065 43.320 296.320 43.780 ;
        RECT 296.490 43.150 296.750 43.610 ;
        RECT 295.630 42.980 296.750 43.150 ;
        RECT 296.920 42.980 297.230 43.780 ;
        RECT 295.630 42.730 295.890 42.980 ;
        RECT 297.400 42.810 297.710 43.610 ;
        RECT 290.535 42.050 290.940 42.560 ;
        RECT 292.080 42.390 292.250 42.640 ;
        RECT 291.110 42.220 292.250 42.390 ;
        RECT 290.535 41.880 292.185 42.050 ;
        RECT 292.420 41.900 292.770 42.470 ;
        RECT 290.580 41.230 290.860 41.710 ;
        RECT 291.030 41.490 291.290 41.880 ;
        RECT 291.465 41.230 291.720 41.710 ;
        RECT 291.890 41.490 292.185 41.880 ;
        RECT 292.940 41.730 293.110 42.640 ;
        RECT 292.365 41.230 292.640 41.710 ;
        RECT 292.810 41.400 293.110 41.730 ;
        RECT 293.280 42.000 294.030 42.520 ;
        RECT 294.200 42.170 294.950 42.690 ;
        RECT 295.135 42.560 295.890 42.730 ;
        RECT 296.680 42.640 297.710 42.810 ;
        RECT 295.135 42.050 295.540 42.560 ;
        RECT 296.680 42.390 296.850 42.640 ;
        RECT 295.710 42.220 296.850 42.390 ;
        RECT 293.280 41.230 294.950 42.000 ;
        RECT 295.135 41.880 296.785 42.050 ;
        RECT 297.020 41.900 297.370 42.470 ;
        RECT 295.180 41.230 295.460 41.710 ;
        RECT 295.630 41.490 295.890 41.880 ;
        RECT 296.065 41.230 296.320 41.710 ;
        RECT 296.490 41.490 296.785 41.880 ;
        RECT 297.540 41.730 297.710 42.640 ;
        RECT 296.965 41.230 297.240 41.710 ;
        RECT 297.410 41.400 297.710 41.730 ;
        RECT 297.880 42.640 298.265 43.610 ;
        RECT 298.435 43.320 298.760 43.780 ;
        RECT 299.280 43.150 299.560 43.610 ;
        RECT 298.435 42.930 299.560 43.150 ;
        RECT 297.880 41.970 298.160 42.640 ;
        RECT 298.435 42.470 298.885 42.930 ;
        RECT 299.750 42.760 300.150 43.610 ;
        RECT 300.550 43.320 300.820 43.780 ;
        RECT 300.990 43.150 301.275 43.610 ;
        RECT 298.330 42.140 298.885 42.470 ;
        RECT 299.055 42.200 300.150 42.760 ;
        RECT 298.435 42.030 298.885 42.140 ;
        RECT 297.880 41.400 298.265 41.970 ;
        RECT 298.435 41.860 299.560 42.030 ;
        RECT 298.435 41.230 298.760 41.690 ;
        RECT 299.280 41.400 299.560 41.860 ;
        RECT 299.750 41.400 300.150 42.200 ;
        RECT 300.320 42.930 301.275 43.150 ;
        RECT 300.320 42.030 300.530 42.930 ;
        RECT 302.020 42.810 302.290 43.580 ;
        RECT 302.460 43.000 302.790 43.780 ;
        RECT 302.995 43.175 303.180 43.580 ;
        RECT 303.350 43.355 303.685 43.780 ;
        RECT 302.995 43.000 303.660 43.175 ;
        RECT 300.700 42.200 301.390 42.760 ;
        RECT 302.020 42.640 303.150 42.810 ;
        RECT 300.320 41.860 301.275 42.030 ;
        RECT 300.550 41.230 300.820 41.690 ;
        RECT 300.990 41.400 301.275 41.860 ;
        RECT 302.020 41.730 302.190 42.640 ;
        RECT 302.360 41.890 302.720 42.470 ;
        RECT 302.900 42.140 303.150 42.640 ;
        RECT 303.320 41.970 303.660 43.000 ;
        RECT 303.860 42.615 304.150 43.780 ;
        RECT 305.240 42.810 305.550 43.610 ;
        RECT 305.720 42.980 306.030 43.780 ;
        RECT 306.200 43.150 306.460 43.610 ;
        RECT 306.630 43.320 306.885 43.780 ;
        RECT 307.060 43.150 307.320 43.610 ;
        RECT 306.200 42.980 307.320 43.150 ;
        RECT 305.240 42.640 306.270 42.810 ;
        RECT 302.975 41.800 303.660 41.970 ;
        RECT 302.020 41.400 302.280 41.730 ;
        RECT 302.490 41.230 302.765 41.710 ;
        RECT 302.975 41.400 303.180 41.800 ;
        RECT 303.350 41.230 303.685 41.630 ;
        RECT 303.860 41.230 304.150 41.955 ;
        RECT 305.240 41.730 305.410 42.640 ;
        RECT 305.580 41.900 305.930 42.470 ;
        RECT 306.100 42.390 306.270 42.640 ;
        RECT 307.060 42.730 307.320 42.980 ;
        RECT 307.490 42.910 307.775 43.780 ;
        RECT 307.060 42.560 307.815 42.730 ;
        RECT 308.000 42.690 309.670 43.780 ;
        RECT 306.100 42.220 307.240 42.390 ;
        RECT 307.410 42.050 307.815 42.560 ;
        RECT 306.165 41.880 307.815 42.050 ;
        RECT 308.000 42.000 308.750 42.520 ;
        RECT 308.920 42.170 309.670 42.690 ;
        RECT 309.840 42.690 311.050 43.780 ;
        RECT 309.840 42.150 310.360 42.690 ;
        RECT 305.240 41.400 305.540 41.730 ;
        RECT 305.710 41.230 305.985 41.710 ;
        RECT 306.165 41.490 306.460 41.880 ;
        RECT 306.630 41.230 306.885 41.710 ;
        RECT 307.060 41.490 307.320 41.880 ;
        RECT 307.490 41.230 307.770 41.710 ;
        RECT 308.000 41.230 309.670 42.000 ;
        RECT 310.530 41.980 311.050 42.520 ;
        RECT 309.840 41.230 311.050 41.980 ;
        RECT 162.095 41.060 311.135 41.230 ;
        RECT 162.180 40.310 163.390 41.060 ;
        RECT 164.485 40.510 164.740 40.800 ;
        RECT 164.910 40.680 165.240 41.060 ;
        RECT 164.485 40.340 165.235 40.510 ;
        RECT 162.180 39.770 162.700 40.310 ;
        RECT 162.870 39.600 163.390 40.140 ;
        RECT 162.180 38.510 163.390 39.600 ;
        RECT 164.485 39.520 164.835 40.170 ;
        RECT 165.005 39.350 165.235 40.340 ;
        RECT 164.485 39.180 165.235 39.350 ;
        RECT 164.485 38.680 164.740 39.180 ;
        RECT 164.910 38.510 165.240 39.010 ;
        RECT 165.410 38.680 165.580 40.800 ;
        RECT 165.940 40.700 166.270 41.060 ;
        RECT 166.440 40.670 166.935 40.840 ;
        RECT 167.140 40.670 167.995 40.840 ;
        RECT 165.810 39.480 166.270 40.530 ;
        RECT 165.750 38.695 166.075 39.480 ;
        RECT 166.440 39.310 166.610 40.670 ;
        RECT 166.780 39.760 167.130 40.380 ;
        RECT 167.300 40.160 167.655 40.380 ;
        RECT 167.300 39.570 167.470 40.160 ;
        RECT 167.825 39.960 167.995 40.670 ;
        RECT 168.870 40.600 169.200 41.060 ;
        RECT 169.410 40.700 169.760 40.870 ;
        RECT 168.200 40.130 168.990 40.380 ;
        RECT 169.410 40.310 169.670 40.700 ;
        RECT 169.980 40.610 170.930 40.890 ;
        RECT 171.100 40.620 171.290 41.060 ;
        RECT 171.460 40.680 172.530 40.850 ;
        RECT 169.160 39.960 169.330 40.140 ;
        RECT 166.440 39.140 166.835 39.310 ;
        RECT 167.005 39.180 167.470 39.570 ;
        RECT 167.640 39.790 169.330 39.960 ;
        RECT 166.665 39.010 166.835 39.140 ;
        RECT 167.640 39.010 167.810 39.790 ;
        RECT 169.500 39.620 169.670 40.310 ;
        RECT 168.170 39.450 169.670 39.620 ;
        RECT 169.860 39.650 170.070 40.440 ;
        RECT 170.240 39.820 170.590 40.440 ;
        RECT 170.760 39.830 170.930 40.610 ;
        RECT 171.460 40.450 171.630 40.680 ;
        RECT 171.100 40.280 171.630 40.450 ;
        RECT 171.100 40.000 171.320 40.280 ;
        RECT 171.800 40.110 172.040 40.510 ;
        RECT 170.760 39.660 171.165 39.830 ;
        RECT 171.500 39.740 172.040 40.110 ;
        RECT 172.210 40.325 172.530 40.680 ;
        RECT 172.775 40.600 173.080 41.060 ;
        RECT 173.250 40.350 173.505 40.880 ;
        RECT 172.210 40.150 172.535 40.325 ;
        RECT 172.210 39.850 173.125 40.150 ;
        RECT 172.385 39.820 173.125 39.850 ;
        RECT 169.860 39.490 170.535 39.650 ;
        RECT 170.995 39.570 171.165 39.660 ;
        RECT 169.860 39.480 170.825 39.490 ;
        RECT 169.500 39.310 169.670 39.450 ;
        RECT 166.245 38.510 166.495 38.970 ;
        RECT 166.665 38.680 166.915 39.010 ;
        RECT 167.130 38.680 167.810 39.010 ;
        RECT 167.980 39.110 169.055 39.280 ;
        RECT 169.500 39.140 170.060 39.310 ;
        RECT 170.365 39.190 170.825 39.480 ;
        RECT 170.995 39.400 172.215 39.570 ;
        RECT 167.980 38.770 168.150 39.110 ;
        RECT 168.385 38.510 168.715 38.940 ;
        RECT 168.885 38.770 169.055 39.110 ;
        RECT 169.350 38.510 169.720 38.970 ;
        RECT 169.890 38.680 170.060 39.140 ;
        RECT 170.995 39.020 171.165 39.400 ;
        RECT 172.385 39.230 172.555 39.820 ;
        RECT 173.295 39.700 173.505 40.350 ;
        RECT 170.295 38.680 171.165 39.020 ;
        RECT 171.755 39.060 172.555 39.230 ;
        RECT 171.335 38.510 171.585 38.970 ;
        RECT 171.755 38.770 171.925 39.060 ;
        RECT 172.105 38.510 172.435 38.890 ;
        RECT 172.775 38.510 173.080 39.650 ;
        RECT 173.250 38.820 173.505 39.700 ;
        RECT 173.685 40.350 173.940 40.880 ;
        RECT 174.110 40.600 174.415 41.060 ;
        RECT 174.660 40.680 175.730 40.850 ;
        RECT 173.685 39.700 173.895 40.350 ;
        RECT 174.660 40.325 174.980 40.680 ;
        RECT 174.655 40.150 174.980 40.325 ;
        RECT 174.065 39.850 174.980 40.150 ;
        RECT 175.150 40.110 175.390 40.510 ;
        RECT 175.560 40.450 175.730 40.680 ;
        RECT 175.900 40.620 176.090 41.060 ;
        RECT 176.260 40.610 177.210 40.890 ;
        RECT 177.430 40.700 177.780 40.870 ;
        RECT 175.560 40.280 176.090 40.450 ;
        RECT 174.065 39.820 174.805 39.850 ;
        RECT 173.685 38.820 173.940 39.700 ;
        RECT 174.110 38.510 174.415 39.650 ;
        RECT 174.635 39.230 174.805 39.820 ;
        RECT 175.150 39.740 175.690 40.110 ;
        RECT 175.870 40.000 176.090 40.280 ;
        RECT 176.260 39.830 176.430 40.610 ;
        RECT 176.025 39.660 176.430 39.830 ;
        RECT 176.600 39.820 176.950 40.440 ;
        RECT 176.025 39.570 176.195 39.660 ;
        RECT 177.120 39.650 177.330 40.440 ;
        RECT 174.975 39.400 176.195 39.570 ;
        RECT 176.655 39.490 177.330 39.650 ;
        RECT 174.635 39.060 175.435 39.230 ;
        RECT 174.755 38.510 175.085 38.890 ;
        RECT 175.265 38.770 175.435 39.060 ;
        RECT 176.025 39.020 176.195 39.400 ;
        RECT 176.365 39.480 177.330 39.490 ;
        RECT 177.520 40.310 177.780 40.700 ;
        RECT 177.990 40.600 178.320 41.060 ;
        RECT 179.195 40.670 180.050 40.840 ;
        RECT 180.255 40.670 180.750 40.840 ;
        RECT 180.920 40.700 181.250 41.060 ;
        RECT 177.520 39.620 177.690 40.310 ;
        RECT 177.860 39.960 178.030 40.140 ;
        RECT 178.200 40.130 178.990 40.380 ;
        RECT 179.195 39.960 179.365 40.670 ;
        RECT 179.535 40.160 179.890 40.380 ;
        RECT 177.860 39.790 179.550 39.960 ;
        RECT 176.365 39.190 176.825 39.480 ;
        RECT 177.520 39.450 179.020 39.620 ;
        RECT 177.520 39.310 177.690 39.450 ;
        RECT 177.130 39.140 177.690 39.310 ;
        RECT 175.605 38.510 175.855 38.970 ;
        RECT 176.025 38.680 176.895 39.020 ;
        RECT 177.130 38.680 177.300 39.140 ;
        RECT 178.135 39.110 179.210 39.280 ;
        RECT 177.470 38.510 177.840 38.970 ;
        RECT 178.135 38.770 178.305 39.110 ;
        RECT 178.475 38.510 178.805 38.940 ;
        RECT 179.040 38.770 179.210 39.110 ;
        RECT 179.380 39.010 179.550 39.790 ;
        RECT 179.720 39.570 179.890 40.160 ;
        RECT 180.060 39.760 180.410 40.380 ;
        RECT 179.720 39.180 180.185 39.570 ;
        RECT 180.580 39.310 180.750 40.670 ;
        RECT 180.920 39.480 181.380 40.530 ;
        RECT 180.355 39.140 180.750 39.310 ;
        RECT 180.355 39.010 180.525 39.140 ;
        RECT 179.380 38.680 180.060 39.010 ;
        RECT 180.275 38.680 180.525 39.010 ;
        RECT 180.695 38.510 180.945 38.970 ;
        RECT 181.115 38.695 181.440 39.480 ;
        RECT 181.610 38.680 181.780 40.800 ;
        RECT 181.950 40.680 182.280 41.060 ;
        RECT 182.450 40.510 182.705 40.800 ;
        RECT 181.955 40.340 182.705 40.510 ;
        RECT 181.955 39.350 182.185 40.340 ;
        RECT 182.880 40.320 183.265 40.890 ;
        RECT 183.435 40.600 183.760 41.060 ;
        RECT 184.280 40.430 184.560 40.890 ;
        RECT 182.355 39.520 182.705 40.170 ;
        RECT 182.880 39.650 183.160 40.320 ;
        RECT 183.435 40.260 184.560 40.430 ;
        RECT 183.435 40.150 183.885 40.260 ;
        RECT 183.330 39.820 183.885 40.150 ;
        RECT 184.750 40.090 185.150 40.890 ;
        RECT 185.550 40.600 185.820 41.060 ;
        RECT 185.990 40.430 186.275 40.890 ;
        RECT 181.955 39.180 182.705 39.350 ;
        RECT 181.950 38.510 182.280 39.010 ;
        RECT 182.450 38.680 182.705 39.180 ;
        RECT 182.880 38.680 183.265 39.650 ;
        RECT 183.435 39.360 183.885 39.820 ;
        RECT 184.055 39.530 185.150 40.090 ;
        RECT 183.435 39.140 184.560 39.360 ;
        RECT 183.435 38.510 183.760 38.970 ;
        RECT 184.280 38.680 184.560 39.140 ;
        RECT 184.750 38.680 185.150 39.530 ;
        RECT 185.320 40.260 186.275 40.430 ;
        RECT 186.560 40.385 186.820 40.890 ;
        RECT 187.000 40.680 187.330 41.060 ;
        RECT 187.510 40.510 187.680 40.890 ;
        RECT 185.320 39.360 185.530 40.260 ;
        RECT 185.700 39.530 186.390 40.090 ;
        RECT 186.560 39.585 186.730 40.385 ;
        RECT 187.015 40.340 187.680 40.510 ;
        RECT 187.015 40.085 187.185 40.340 ;
        RECT 187.940 40.335 188.230 41.060 ;
        RECT 188.400 40.310 189.610 41.060 ;
        RECT 189.870 40.510 190.040 40.890 ;
        RECT 190.220 40.680 190.550 41.060 ;
        RECT 189.870 40.340 190.535 40.510 ;
        RECT 190.730 40.385 190.990 40.890 ;
        RECT 186.900 39.755 187.185 40.085 ;
        RECT 187.420 39.790 187.750 40.160 ;
        RECT 188.400 39.770 188.920 40.310 ;
        RECT 187.015 39.610 187.185 39.755 ;
        RECT 185.320 39.140 186.275 39.360 ;
        RECT 185.550 38.510 185.820 38.970 ;
        RECT 185.990 38.680 186.275 39.140 ;
        RECT 186.560 38.680 186.830 39.585 ;
        RECT 187.015 39.440 187.680 39.610 ;
        RECT 187.000 38.510 187.330 39.270 ;
        RECT 187.510 38.680 187.680 39.440 ;
        RECT 187.940 38.510 188.230 39.675 ;
        RECT 189.090 39.600 189.610 40.140 ;
        RECT 189.800 39.790 190.130 40.160 ;
        RECT 190.365 40.085 190.535 40.340 ;
        RECT 190.365 39.755 190.650 40.085 ;
        RECT 190.365 39.610 190.535 39.755 ;
        RECT 188.400 38.510 189.610 39.600 ;
        RECT 189.870 39.440 190.535 39.610 ;
        RECT 190.820 39.585 190.990 40.385 ;
        RECT 189.870 38.680 190.040 39.440 ;
        RECT 190.220 38.510 190.550 39.270 ;
        RECT 190.720 38.680 190.990 39.585 ;
        RECT 191.160 40.385 191.420 40.890 ;
        RECT 191.600 40.680 191.930 41.060 ;
        RECT 192.110 40.510 192.280 40.890 ;
        RECT 191.160 39.585 191.330 40.385 ;
        RECT 191.615 40.340 192.280 40.510 ;
        RECT 191.615 40.085 191.785 40.340 ;
        RECT 192.540 40.310 193.750 41.060 ;
        RECT 193.925 40.320 194.180 40.890 ;
        RECT 194.350 40.660 194.680 41.060 ;
        RECT 195.105 40.525 195.635 40.890 ;
        RECT 195.825 40.720 196.100 40.890 ;
        RECT 195.820 40.550 196.100 40.720 ;
        RECT 195.105 40.490 195.280 40.525 ;
        RECT 194.350 40.320 195.280 40.490 ;
        RECT 191.500 39.755 191.785 40.085 ;
        RECT 192.020 39.790 192.350 40.160 ;
        RECT 192.540 39.770 193.060 40.310 ;
        RECT 191.615 39.610 191.785 39.755 ;
        RECT 191.160 38.680 191.430 39.585 ;
        RECT 191.615 39.440 192.280 39.610 ;
        RECT 193.230 39.600 193.750 40.140 ;
        RECT 191.600 38.510 191.930 39.270 ;
        RECT 192.110 38.680 192.280 39.440 ;
        RECT 192.540 38.510 193.750 39.600 ;
        RECT 193.925 39.650 194.095 40.320 ;
        RECT 194.350 40.150 194.520 40.320 ;
        RECT 194.265 39.820 194.520 40.150 ;
        RECT 194.745 39.820 194.940 40.150 ;
        RECT 193.925 38.680 194.260 39.650 ;
        RECT 194.430 38.510 194.600 39.650 ;
        RECT 194.770 38.850 194.940 39.820 ;
        RECT 195.110 39.190 195.280 40.320 ;
        RECT 195.450 39.530 195.620 40.330 ;
        RECT 195.825 39.730 196.100 40.550 ;
        RECT 196.270 39.530 196.460 40.890 ;
        RECT 196.640 40.525 197.150 41.060 ;
        RECT 197.370 40.250 197.615 40.855 ;
        RECT 198.060 40.320 198.445 40.890 ;
        RECT 198.615 40.600 198.940 41.060 ;
        RECT 199.460 40.430 199.740 40.890 ;
        RECT 196.660 40.080 197.890 40.250 ;
        RECT 195.450 39.360 196.460 39.530 ;
        RECT 196.630 39.515 197.380 39.705 ;
        RECT 195.110 39.020 196.235 39.190 ;
        RECT 196.630 38.850 196.800 39.515 ;
        RECT 197.550 39.270 197.890 40.080 ;
        RECT 194.770 38.680 196.800 38.850 ;
        RECT 196.970 38.510 197.140 39.270 ;
        RECT 197.375 38.860 197.890 39.270 ;
        RECT 198.060 39.650 198.340 40.320 ;
        RECT 198.615 40.260 199.740 40.430 ;
        RECT 198.615 40.150 199.065 40.260 ;
        RECT 198.510 39.820 199.065 40.150 ;
        RECT 199.930 40.090 200.330 40.890 ;
        RECT 200.730 40.600 201.000 41.060 ;
        RECT 201.170 40.430 201.455 40.890 ;
        RECT 198.060 38.680 198.445 39.650 ;
        RECT 198.615 39.360 199.065 39.820 ;
        RECT 199.235 39.530 200.330 40.090 ;
        RECT 198.615 39.140 199.740 39.360 ;
        RECT 198.615 38.510 198.940 38.970 ;
        RECT 199.460 38.680 199.740 39.140 ;
        RECT 199.930 38.680 200.330 39.530 ;
        RECT 200.500 40.260 201.455 40.430 ;
        RECT 201.740 40.310 202.950 41.060 ;
        RECT 200.500 39.360 200.710 40.260 ;
        RECT 200.880 39.530 201.570 40.090 ;
        RECT 201.740 39.770 202.260 40.310 ;
        RECT 203.160 40.240 203.390 41.060 ;
        RECT 203.560 40.260 203.890 40.890 ;
        RECT 202.430 39.600 202.950 40.140 ;
        RECT 203.140 39.820 203.470 40.070 ;
        RECT 203.640 39.660 203.890 40.260 ;
        RECT 204.060 40.240 204.270 41.060 ;
        RECT 204.505 40.510 204.760 40.800 ;
        RECT 204.930 40.680 205.260 41.060 ;
        RECT 204.505 40.340 205.255 40.510 ;
        RECT 200.500 39.140 201.455 39.360 ;
        RECT 200.730 38.510 201.000 38.970 ;
        RECT 201.170 38.680 201.455 39.140 ;
        RECT 201.740 38.510 202.950 39.600 ;
        RECT 203.160 38.510 203.390 39.650 ;
        RECT 203.560 38.680 203.890 39.660 ;
        RECT 204.060 38.510 204.270 39.650 ;
        RECT 204.505 39.520 204.855 40.170 ;
        RECT 205.025 39.350 205.255 40.340 ;
        RECT 204.505 39.180 205.255 39.350 ;
        RECT 204.505 38.680 204.760 39.180 ;
        RECT 204.930 38.510 205.260 39.010 ;
        RECT 205.430 38.680 205.600 40.800 ;
        RECT 205.960 40.700 206.290 41.060 ;
        RECT 206.460 40.670 206.955 40.840 ;
        RECT 207.160 40.670 208.015 40.840 ;
        RECT 205.830 39.480 206.290 40.530 ;
        RECT 205.770 38.695 206.095 39.480 ;
        RECT 206.460 39.310 206.630 40.670 ;
        RECT 206.800 39.760 207.150 40.380 ;
        RECT 207.320 40.160 207.675 40.380 ;
        RECT 207.320 39.570 207.490 40.160 ;
        RECT 207.845 39.960 208.015 40.670 ;
        RECT 208.890 40.600 209.220 41.060 ;
        RECT 209.430 40.700 209.780 40.870 ;
        RECT 208.220 40.130 209.010 40.380 ;
        RECT 209.430 40.310 209.690 40.700 ;
        RECT 210.000 40.610 210.950 40.890 ;
        RECT 211.120 40.620 211.310 41.060 ;
        RECT 211.480 40.680 212.550 40.850 ;
        RECT 209.180 39.960 209.350 40.140 ;
        RECT 206.460 39.140 206.855 39.310 ;
        RECT 207.025 39.180 207.490 39.570 ;
        RECT 207.660 39.790 209.350 39.960 ;
        RECT 206.685 39.010 206.855 39.140 ;
        RECT 207.660 39.010 207.830 39.790 ;
        RECT 209.520 39.620 209.690 40.310 ;
        RECT 208.190 39.450 209.690 39.620 ;
        RECT 209.880 39.650 210.090 40.440 ;
        RECT 210.260 39.820 210.610 40.440 ;
        RECT 210.780 39.830 210.950 40.610 ;
        RECT 211.480 40.450 211.650 40.680 ;
        RECT 211.120 40.280 211.650 40.450 ;
        RECT 211.120 40.000 211.340 40.280 ;
        RECT 211.820 40.110 212.060 40.510 ;
        RECT 210.780 39.660 211.185 39.830 ;
        RECT 211.520 39.740 212.060 40.110 ;
        RECT 212.230 40.325 212.550 40.680 ;
        RECT 212.795 40.600 213.100 41.060 ;
        RECT 213.270 40.350 213.525 40.880 ;
        RECT 212.230 40.150 212.555 40.325 ;
        RECT 212.230 39.850 213.145 40.150 ;
        RECT 212.405 39.820 213.145 39.850 ;
        RECT 209.880 39.490 210.555 39.650 ;
        RECT 211.015 39.570 211.185 39.660 ;
        RECT 209.880 39.480 210.845 39.490 ;
        RECT 209.520 39.310 209.690 39.450 ;
        RECT 206.265 38.510 206.515 38.970 ;
        RECT 206.685 38.680 206.935 39.010 ;
        RECT 207.150 38.680 207.830 39.010 ;
        RECT 208.000 39.110 209.075 39.280 ;
        RECT 209.520 39.140 210.080 39.310 ;
        RECT 210.385 39.190 210.845 39.480 ;
        RECT 211.015 39.400 212.235 39.570 ;
        RECT 208.000 38.770 208.170 39.110 ;
        RECT 208.405 38.510 208.735 38.940 ;
        RECT 208.905 38.770 209.075 39.110 ;
        RECT 209.370 38.510 209.740 38.970 ;
        RECT 209.910 38.680 210.080 39.140 ;
        RECT 211.015 39.020 211.185 39.400 ;
        RECT 212.405 39.230 212.575 39.820 ;
        RECT 213.315 39.700 213.525 40.350 ;
        RECT 213.700 40.335 213.990 41.060 ;
        RECT 214.160 40.515 219.505 41.060 ;
        RECT 210.315 38.680 211.185 39.020 ;
        RECT 211.775 39.060 212.575 39.230 ;
        RECT 211.355 38.510 211.605 38.970 ;
        RECT 211.775 38.770 211.945 39.060 ;
        RECT 212.125 38.510 212.455 38.890 ;
        RECT 212.795 38.510 213.100 39.650 ;
        RECT 213.270 38.820 213.525 39.700 ;
        RECT 215.745 39.685 216.085 40.515 ;
        RECT 219.680 40.385 219.940 40.890 ;
        RECT 220.120 40.680 220.450 41.060 ;
        RECT 220.630 40.510 220.800 40.890 ;
        RECT 213.700 38.510 213.990 39.675 ;
        RECT 217.565 38.945 217.915 40.195 ;
        RECT 219.680 39.585 219.850 40.385 ;
        RECT 220.135 40.340 220.800 40.510 ;
        RECT 221.150 40.510 221.320 40.890 ;
        RECT 221.500 40.680 221.830 41.060 ;
        RECT 221.150 40.340 221.815 40.510 ;
        RECT 222.010 40.385 222.270 40.890 ;
        RECT 220.135 40.085 220.305 40.340 ;
        RECT 220.020 39.755 220.305 40.085 ;
        RECT 220.540 39.790 220.870 40.160 ;
        RECT 221.080 39.790 221.410 40.160 ;
        RECT 221.645 40.085 221.815 40.340 ;
        RECT 220.135 39.610 220.305 39.755 ;
        RECT 221.645 39.755 221.930 40.085 ;
        RECT 221.645 39.610 221.815 39.755 ;
        RECT 214.160 38.510 219.505 38.945 ;
        RECT 219.680 38.680 219.950 39.585 ;
        RECT 220.135 39.440 220.800 39.610 ;
        RECT 220.120 38.510 220.450 39.270 ;
        RECT 220.630 38.680 220.800 39.440 ;
        RECT 221.150 39.440 221.815 39.610 ;
        RECT 222.100 39.585 222.270 40.385 ;
        RECT 221.150 38.680 221.320 39.440 ;
        RECT 221.500 38.510 221.830 39.270 ;
        RECT 222.000 38.680 222.270 39.585 ;
        RECT 222.445 40.320 222.700 40.890 ;
        RECT 222.870 40.660 223.200 41.060 ;
        RECT 223.625 40.525 224.155 40.890 ;
        RECT 224.345 40.720 224.620 40.890 ;
        RECT 224.340 40.550 224.620 40.720 ;
        RECT 223.625 40.490 223.800 40.525 ;
        RECT 222.870 40.320 223.800 40.490 ;
        RECT 222.445 39.650 222.615 40.320 ;
        RECT 222.870 40.150 223.040 40.320 ;
        RECT 222.785 39.820 223.040 40.150 ;
        RECT 223.265 39.820 223.460 40.150 ;
        RECT 222.445 38.680 222.780 39.650 ;
        RECT 222.950 38.510 223.120 39.650 ;
        RECT 223.290 38.850 223.460 39.820 ;
        RECT 223.630 39.190 223.800 40.320 ;
        RECT 223.970 39.530 224.140 40.330 ;
        RECT 224.345 39.730 224.620 40.550 ;
        RECT 224.790 39.530 224.980 40.890 ;
        RECT 225.160 40.525 225.670 41.060 ;
        RECT 225.890 40.250 226.135 40.855 ;
        RECT 227.130 40.510 227.300 40.890 ;
        RECT 227.480 40.680 227.810 41.060 ;
        RECT 227.130 40.340 227.795 40.510 ;
        RECT 227.990 40.385 228.250 40.890 ;
        RECT 225.180 40.080 226.410 40.250 ;
        RECT 223.970 39.360 224.980 39.530 ;
        RECT 225.150 39.515 225.900 39.705 ;
        RECT 223.630 39.020 224.755 39.190 ;
        RECT 225.150 38.850 225.320 39.515 ;
        RECT 226.070 39.270 226.410 40.080 ;
        RECT 227.060 39.790 227.390 40.160 ;
        RECT 227.625 40.085 227.795 40.340 ;
        RECT 227.625 39.755 227.910 40.085 ;
        RECT 227.625 39.610 227.795 39.755 ;
        RECT 223.290 38.680 225.320 38.850 ;
        RECT 225.490 38.510 225.660 39.270 ;
        RECT 225.895 38.860 226.410 39.270 ;
        RECT 227.130 39.440 227.795 39.610 ;
        RECT 228.080 39.585 228.250 40.385 ;
        RECT 227.130 38.680 227.300 39.440 ;
        RECT 227.480 38.510 227.810 39.270 ;
        RECT 227.980 38.680 228.250 39.585 ;
        RECT 228.425 40.320 228.680 40.890 ;
        RECT 228.850 40.660 229.180 41.060 ;
        RECT 229.605 40.525 230.135 40.890 ;
        RECT 230.325 40.720 230.600 40.890 ;
        RECT 230.320 40.550 230.600 40.720 ;
        RECT 229.605 40.490 229.780 40.525 ;
        RECT 228.850 40.320 229.780 40.490 ;
        RECT 228.425 39.650 228.595 40.320 ;
        RECT 228.850 40.150 229.020 40.320 ;
        RECT 228.765 39.820 229.020 40.150 ;
        RECT 229.245 39.820 229.440 40.150 ;
        RECT 228.425 38.680 228.760 39.650 ;
        RECT 228.930 38.510 229.100 39.650 ;
        RECT 229.270 38.850 229.440 39.820 ;
        RECT 229.610 39.190 229.780 40.320 ;
        RECT 229.950 39.530 230.120 40.330 ;
        RECT 230.325 39.730 230.600 40.550 ;
        RECT 230.770 39.530 230.960 40.890 ;
        RECT 231.140 40.525 231.650 41.060 ;
        RECT 231.870 40.250 232.115 40.855 ;
        RECT 232.565 40.320 232.820 40.890 ;
        RECT 232.990 40.660 233.320 41.060 ;
        RECT 233.745 40.525 234.275 40.890 ;
        RECT 234.465 40.720 234.740 40.890 ;
        RECT 234.460 40.550 234.740 40.720 ;
        RECT 233.745 40.490 233.920 40.525 ;
        RECT 232.990 40.320 233.920 40.490 ;
        RECT 231.160 40.080 232.390 40.250 ;
        RECT 229.950 39.360 230.960 39.530 ;
        RECT 231.130 39.515 231.880 39.705 ;
        RECT 229.610 39.020 230.735 39.190 ;
        RECT 231.130 38.850 231.300 39.515 ;
        RECT 232.050 39.270 232.390 40.080 ;
        RECT 229.270 38.680 231.300 38.850 ;
        RECT 231.470 38.510 231.640 39.270 ;
        RECT 231.875 38.860 232.390 39.270 ;
        RECT 232.565 39.650 232.735 40.320 ;
        RECT 232.990 40.150 233.160 40.320 ;
        RECT 232.905 39.820 233.160 40.150 ;
        RECT 233.385 39.820 233.580 40.150 ;
        RECT 232.565 38.680 232.900 39.650 ;
        RECT 233.070 38.510 233.240 39.650 ;
        RECT 233.410 38.850 233.580 39.820 ;
        RECT 233.750 39.190 233.920 40.320 ;
        RECT 234.090 39.530 234.260 40.330 ;
        RECT 234.465 39.730 234.740 40.550 ;
        RECT 234.910 39.530 235.100 40.890 ;
        RECT 235.280 40.525 235.790 41.060 ;
        RECT 236.010 40.250 236.255 40.855 ;
        RECT 236.700 40.290 239.290 41.060 ;
        RECT 239.460 40.335 239.750 41.060 ;
        RECT 240.495 40.430 240.780 40.890 ;
        RECT 240.950 40.600 241.220 41.060 ;
        RECT 235.300 40.080 236.530 40.250 ;
        RECT 234.090 39.360 235.100 39.530 ;
        RECT 235.270 39.515 236.020 39.705 ;
        RECT 233.750 39.020 234.875 39.190 ;
        RECT 235.270 38.850 235.440 39.515 ;
        RECT 236.190 39.270 236.530 40.080 ;
        RECT 236.700 39.770 237.910 40.290 ;
        RECT 240.495 40.260 241.450 40.430 ;
        RECT 238.080 39.600 239.290 40.120 ;
        RECT 233.410 38.680 235.440 38.850 ;
        RECT 235.610 38.510 235.780 39.270 ;
        RECT 236.015 38.860 236.530 39.270 ;
        RECT 236.700 38.510 239.290 39.600 ;
        RECT 239.460 38.510 239.750 39.675 ;
        RECT 240.380 39.530 241.070 40.090 ;
        RECT 241.240 39.360 241.450 40.260 ;
        RECT 240.495 39.140 241.450 39.360 ;
        RECT 241.620 40.090 242.020 40.890 ;
        RECT 242.210 40.430 242.490 40.890 ;
        RECT 243.010 40.600 243.335 41.060 ;
        RECT 242.210 40.260 243.335 40.430 ;
        RECT 243.505 40.320 243.890 40.890 ;
        RECT 242.885 40.150 243.335 40.260 ;
        RECT 241.620 39.530 242.715 40.090 ;
        RECT 242.885 39.820 243.440 40.150 ;
        RECT 240.495 38.680 240.780 39.140 ;
        RECT 240.950 38.510 241.220 38.970 ;
        RECT 241.620 38.680 242.020 39.530 ;
        RECT 242.885 39.360 243.335 39.820 ;
        RECT 243.610 39.650 243.890 40.320 ;
        RECT 242.210 39.140 243.335 39.360 ;
        RECT 242.210 38.680 242.490 39.140 ;
        RECT 243.010 38.510 243.335 38.970 ;
        RECT 243.505 38.680 243.890 39.650 ;
        RECT 244.525 40.320 244.780 40.890 ;
        RECT 244.950 40.660 245.280 41.060 ;
        RECT 245.705 40.525 246.235 40.890 ;
        RECT 245.705 40.490 245.880 40.525 ;
        RECT 244.950 40.320 245.880 40.490 ;
        RECT 244.525 39.650 244.695 40.320 ;
        RECT 244.950 40.150 245.120 40.320 ;
        RECT 244.865 39.820 245.120 40.150 ;
        RECT 245.345 39.820 245.540 40.150 ;
        RECT 244.525 38.680 244.860 39.650 ;
        RECT 245.030 38.510 245.200 39.650 ;
        RECT 245.370 38.850 245.540 39.820 ;
        RECT 245.710 39.190 245.880 40.320 ;
        RECT 246.050 39.530 246.220 40.330 ;
        RECT 246.425 40.040 246.700 40.890 ;
        RECT 246.420 39.870 246.700 40.040 ;
        RECT 246.425 39.730 246.700 39.870 ;
        RECT 246.870 39.530 247.060 40.890 ;
        RECT 247.240 40.525 247.750 41.060 ;
        RECT 247.970 40.250 248.215 40.855 ;
        RECT 248.665 40.510 248.920 40.800 ;
        RECT 249.090 40.680 249.420 41.060 ;
        RECT 248.665 40.340 249.415 40.510 ;
        RECT 247.260 40.080 248.490 40.250 ;
        RECT 246.050 39.360 247.060 39.530 ;
        RECT 247.230 39.515 247.980 39.705 ;
        RECT 245.710 39.020 246.835 39.190 ;
        RECT 247.230 38.850 247.400 39.515 ;
        RECT 248.150 39.270 248.490 40.080 ;
        RECT 248.665 39.520 249.015 40.170 ;
        RECT 249.185 39.350 249.415 40.340 ;
        RECT 245.370 38.680 247.400 38.850 ;
        RECT 247.570 38.510 247.740 39.270 ;
        RECT 247.975 38.860 248.490 39.270 ;
        RECT 248.665 39.180 249.415 39.350 ;
        RECT 248.665 38.680 248.920 39.180 ;
        RECT 249.090 38.510 249.420 39.010 ;
        RECT 249.590 38.680 249.760 40.800 ;
        RECT 250.120 40.700 250.450 41.060 ;
        RECT 250.620 40.670 251.115 40.840 ;
        RECT 251.320 40.670 252.175 40.840 ;
        RECT 249.990 39.480 250.450 40.530 ;
        RECT 249.930 38.695 250.255 39.480 ;
        RECT 250.620 39.310 250.790 40.670 ;
        RECT 250.960 39.760 251.310 40.380 ;
        RECT 251.480 40.160 251.835 40.380 ;
        RECT 251.480 39.570 251.650 40.160 ;
        RECT 252.005 39.960 252.175 40.670 ;
        RECT 253.050 40.600 253.380 41.060 ;
        RECT 253.590 40.700 253.940 40.870 ;
        RECT 252.380 40.130 253.170 40.380 ;
        RECT 253.590 40.310 253.850 40.700 ;
        RECT 254.160 40.610 255.110 40.890 ;
        RECT 255.280 40.620 255.470 41.060 ;
        RECT 255.640 40.680 256.710 40.850 ;
        RECT 253.340 39.960 253.510 40.140 ;
        RECT 250.620 39.140 251.015 39.310 ;
        RECT 251.185 39.180 251.650 39.570 ;
        RECT 251.820 39.790 253.510 39.960 ;
        RECT 250.845 39.010 251.015 39.140 ;
        RECT 251.820 39.010 251.990 39.790 ;
        RECT 253.680 39.620 253.850 40.310 ;
        RECT 252.350 39.450 253.850 39.620 ;
        RECT 254.040 39.650 254.250 40.440 ;
        RECT 254.420 39.820 254.770 40.440 ;
        RECT 254.940 39.830 255.110 40.610 ;
        RECT 255.640 40.450 255.810 40.680 ;
        RECT 255.280 40.280 255.810 40.450 ;
        RECT 255.280 40.000 255.500 40.280 ;
        RECT 255.980 40.110 256.220 40.510 ;
        RECT 254.940 39.660 255.345 39.830 ;
        RECT 255.680 39.740 256.220 40.110 ;
        RECT 256.390 40.325 256.710 40.680 ;
        RECT 256.955 40.600 257.260 41.060 ;
        RECT 257.430 40.350 257.685 40.880 ;
        RECT 256.390 40.150 256.715 40.325 ;
        RECT 256.390 39.850 257.305 40.150 ;
        RECT 256.565 39.820 257.305 39.850 ;
        RECT 254.040 39.490 254.715 39.650 ;
        RECT 255.175 39.570 255.345 39.660 ;
        RECT 254.040 39.480 255.005 39.490 ;
        RECT 253.680 39.310 253.850 39.450 ;
        RECT 250.425 38.510 250.675 38.970 ;
        RECT 250.845 38.680 251.095 39.010 ;
        RECT 251.310 38.680 251.990 39.010 ;
        RECT 252.160 39.110 253.235 39.280 ;
        RECT 253.680 39.140 254.240 39.310 ;
        RECT 254.545 39.190 255.005 39.480 ;
        RECT 255.175 39.400 256.395 39.570 ;
        RECT 252.160 38.770 252.330 39.110 ;
        RECT 252.565 38.510 252.895 38.940 ;
        RECT 253.065 38.770 253.235 39.110 ;
        RECT 253.530 38.510 253.900 38.970 ;
        RECT 254.070 38.680 254.240 39.140 ;
        RECT 255.175 39.020 255.345 39.400 ;
        RECT 256.565 39.230 256.735 39.820 ;
        RECT 257.475 39.700 257.685 40.350 ;
        RECT 254.475 38.680 255.345 39.020 ;
        RECT 255.935 39.060 256.735 39.230 ;
        RECT 255.515 38.510 255.765 38.970 ;
        RECT 255.935 38.770 256.105 39.060 ;
        RECT 256.285 38.510 256.615 38.890 ;
        RECT 256.955 38.510 257.260 39.650 ;
        RECT 257.430 38.820 257.685 39.700 ;
        RECT 257.860 40.320 258.245 40.890 ;
        RECT 258.415 40.600 258.740 41.060 ;
        RECT 259.260 40.430 259.540 40.890 ;
        RECT 257.860 39.650 258.140 40.320 ;
        RECT 258.415 40.260 259.540 40.430 ;
        RECT 258.415 40.150 258.865 40.260 ;
        RECT 258.310 39.820 258.865 40.150 ;
        RECT 259.730 40.090 260.130 40.890 ;
        RECT 260.530 40.600 260.800 41.060 ;
        RECT 260.970 40.430 261.255 40.890 ;
        RECT 257.860 38.680 258.245 39.650 ;
        RECT 258.415 39.360 258.865 39.820 ;
        RECT 259.035 39.530 260.130 40.090 ;
        RECT 258.415 39.140 259.540 39.360 ;
        RECT 258.415 38.510 258.740 38.970 ;
        RECT 259.260 38.680 259.540 39.140 ;
        RECT 259.730 38.680 260.130 39.530 ;
        RECT 260.300 40.260 261.255 40.430 ;
        RECT 261.540 40.320 261.925 40.890 ;
        RECT 262.095 40.600 262.420 41.060 ;
        RECT 262.940 40.430 263.220 40.890 ;
        RECT 260.300 39.360 260.510 40.260 ;
        RECT 260.680 39.530 261.370 40.090 ;
        RECT 261.540 39.650 261.820 40.320 ;
        RECT 262.095 40.260 263.220 40.430 ;
        RECT 262.095 40.150 262.545 40.260 ;
        RECT 261.990 39.820 262.545 40.150 ;
        RECT 263.410 40.090 263.810 40.890 ;
        RECT 264.210 40.600 264.480 41.060 ;
        RECT 264.650 40.430 264.935 40.890 ;
        RECT 260.300 39.140 261.255 39.360 ;
        RECT 260.530 38.510 260.800 38.970 ;
        RECT 260.970 38.680 261.255 39.140 ;
        RECT 261.540 38.680 261.925 39.650 ;
        RECT 262.095 39.360 262.545 39.820 ;
        RECT 262.715 39.530 263.810 40.090 ;
        RECT 262.095 39.140 263.220 39.360 ;
        RECT 262.095 38.510 262.420 38.970 ;
        RECT 262.940 38.680 263.220 39.140 ;
        RECT 263.410 38.680 263.810 39.530 ;
        RECT 263.980 40.260 264.935 40.430 ;
        RECT 265.220 40.335 265.510 41.060 ;
        RECT 265.680 40.290 267.350 41.060 ;
        RECT 267.525 40.510 267.780 40.800 ;
        RECT 267.950 40.680 268.280 41.060 ;
        RECT 267.525 40.340 268.275 40.510 ;
        RECT 263.980 39.360 264.190 40.260 ;
        RECT 264.360 39.530 265.050 40.090 ;
        RECT 265.680 39.770 266.430 40.290 ;
        RECT 263.980 39.140 264.935 39.360 ;
        RECT 264.210 38.510 264.480 38.970 ;
        RECT 264.650 38.680 264.935 39.140 ;
        RECT 265.220 38.510 265.510 39.675 ;
        RECT 266.600 39.600 267.350 40.120 ;
        RECT 265.680 38.510 267.350 39.600 ;
        RECT 267.525 39.520 267.875 40.170 ;
        RECT 268.045 39.350 268.275 40.340 ;
        RECT 267.525 39.180 268.275 39.350 ;
        RECT 267.525 38.680 267.780 39.180 ;
        RECT 267.950 38.510 268.280 39.010 ;
        RECT 268.450 38.680 268.620 40.800 ;
        RECT 268.980 40.700 269.310 41.060 ;
        RECT 269.480 40.670 269.975 40.840 ;
        RECT 270.180 40.670 271.035 40.840 ;
        RECT 268.850 39.480 269.310 40.530 ;
        RECT 268.790 38.695 269.115 39.480 ;
        RECT 269.480 39.310 269.650 40.670 ;
        RECT 269.820 39.760 270.170 40.380 ;
        RECT 270.340 40.160 270.695 40.380 ;
        RECT 270.340 39.570 270.510 40.160 ;
        RECT 270.865 39.960 271.035 40.670 ;
        RECT 271.910 40.600 272.240 41.060 ;
        RECT 272.450 40.700 272.800 40.870 ;
        RECT 271.240 40.130 272.030 40.380 ;
        RECT 272.450 40.310 272.710 40.700 ;
        RECT 273.020 40.610 273.970 40.890 ;
        RECT 274.140 40.620 274.330 41.060 ;
        RECT 274.500 40.680 275.570 40.850 ;
        RECT 272.200 39.960 272.370 40.140 ;
        RECT 269.480 39.140 269.875 39.310 ;
        RECT 270.045 39.180 270.510 39.570 ;
        RECT 270.680 39.790 272.370 39.960 ;
        RECT 269.705 39.010 269.875 39.140 ;
        RECT 270.680 39.010 270.850 39.790 ;
        RECT 272.540 39.620 272.710 40.310 ;
        RECT 271.210 39.450 272.710 39.620 ;
        RECT 272.900 39.650 273.110 40.440 ;
        RECT 273.280 39.820 273.630 40.440 ;
        RECT 273.800 39.830 273.970 40.610 ;
        RECT 274.500 40.450 274.670 40.680 ;
        RECT 274.140 40.280 274.670 40.450 ;
        RECT 274.140 40.000 274.360 40.280 ;
        RECT 274.840 40.110 275.080 40.510 ;
        RECT 273.800 39.660 274.205 39.830 ;
        RECT 274.540 39.740 275.080 40.110 ;
        RECT 275.250 40.325 275.570 40.680 ;
        RECT 275.815 40.600 276.120 41.060 ;
        RECT 276.290 40.350 276.545 40.880 ;
        RECT 275.250 40.150 275.575 40.325 ;
        RECT 275.250 39.850 276.165 40.150 ;
        RECT 275.425 39.820 276.165 39.850 ;
        RECT 272.900 39.490 273.575 39.650 ;
        RECT 274.035 39.570 274.205 39.660 ;
        RECT 272.900 39.480 273.865 39.490 ;
        RECT 272.540 39.310 272.710 39.450 ;
        RECT 269.285 38.510 269.535 38.970 ;
        RECT 269.705 38.680 269.955 39.010 ;
        RECT 270.170 38.680 270.850 39.010 ;
        RECT 271.020 39.110 272.095 39.280 ;
        RECT 272.540 39.140 273.100 39.310 ;
        RECT 273.405 39.190 273.865 39.480 ;
        RECT 274.035 39.400 275.255 39.570 ;
        RECT 271.020 38.770 271.190 39.110 ;
        RECT 271.425 38.510 271.755 38.940 ;
        RECT 271.925 38.770 272.095 39.110 ;
        RECT 272.390 38.510 272.760 38.970 ;
        RECT 272.930 38.680 273.100 39.140 ;
        RECT 274.035 39.020 274.205 39.400 ;
        RECT 275.425 39.230 275.595 39.820 ;
        RECT 276.335 39.700 276.545 40.350 ;
        RECT 276.720 40.290 278.390 41.060 ;
        RECT 278.650 40.410 278.820 40.890 ;
        RECT 278.990 40.580 279.320 41.060 ;
        RECT 279.545 40.640 281.080 40.890 ;
        RECT 279.545 40.410 279.715 40.640 ;
        RECT 276.720 39.770 277.470 40.290 ;
        RECT 278.650 40.240 279.715 40.410 ;
        RECT 273.335 38.680 274.205 39.020 ;
        RECT 274.795 39.060 275.595 39.230 ;
        RECT 274.375 38.510 274.625 38.970 ;
        RECT 274.795 38.770 274.965 39.060 ;
        RECT 275.145 38.510 275.475 38.890 ;
        RECT 275.815 38.510 276.120 39.650 ;
        RECT 276.290 38.820 276.545 39.700 ;
        RECT 277.640 39.600 278.390 40.120 ;
        RECT 279.895 40.070 280.175 40.470 ;
        RECT 278.565 39.860 278.915 40.070 ;
        RECT 279.085 39.870 279.530 40.070 ;
        RECT 279.700 39.870 280.175 40.070 ;
        RECT 280.445 40.070 280.730 40.470 ;
        RECT 280.910 40.410 281.080 40.640 ;
        RECT 281.250 40.580 281.580 41.060 ;
        RECT 281.795 40.560 282.050 40.890 ;
        RECT 281.840 40.550 282.050 40.560 ;
        RECT 281.865 40.480 282.050 40.550 ;
        RECT 282.240 40.515 287.585 41.060 ;
        RECT 280.910 40.240 281.710 40.410 ;
        RECT 280.445 39.870 280.775 40.070 ;
        RECT 280.945 40.040 281.310 40.070 ;
        RECT 280.945 39.870 281.320 40.040 ;
        RECT 281.540 39.690 281.710 40.240 ;
        RECT 276.720 38.510 278.390 39.600 ;
        RECT 278.650 39.520 281.710 39.690 ;
        RECT 278.650 38.680 278.820 39.520 ;
        RECT 281.880 39.350 282.050 40.480 ;
        RECT 283.825 39.685 284.165 40.515 ;
        RECT 287.760 40.310 288.970 41.060 ;
        RECT 278.990 38.850 279.320 39.350 ;
        RECT 279.490 39.110 281.125 39.350 ;
        RECT 279.490 39.020 279.720 39.110 ;
        RECT 279.830 38.850 280.160 38.890 ;
        RECT 278.990 38.680 280.160 38.850 ;
        RECT 280.350 38.510 280.705 38.930 ;
        RECT 280.875 38.680 281.125 39.110 ;
        RECT 281.295 38.510 281.625 39.270 ;
        RECT 281.795 38.680 282.050 39.350 ;
        RECT 285.645 38.945 285.995 40.195 ;
        RECT 287.760 39.770 288.280 40.310 ;
        RECT 289.145 40.220 289.405 41.060 ;
        RECT 289.580 40.315 289.835 40.890 ;
        RECT 290.005 40.680 290.335 41.060 ;
        RECT 290.550 40.510 290.720 40.890 ;
        RECT 290.005 40.340 290.720 40.510 ;
        RECT 288.450 39.600 288.970 40.140 ;
        RECT 282.240 38.510 287.585 38.945 ;
        RECT 287.760 38.510 288.970 39.600 ;
        RECT 289.145 38.510 289.405 39.660 ;
        RECT 289.580 39.585 289.750 40.315 ;
        RECT 290.005 40.150 290.175 40.340 ;
        RECT 290.980 40.335 291.270 41.060 ;
        RECT 291.445 40.340 291.780 41.060 ;
        RECT 291.950 40.530 292.140 40.775 ;
        RECT 292.310 40.700 292.640 41.060 ;
        RECT 292.810 40.530 293.000 40.890 ;
        RECT 293.190 40.620 293.470 41.060 ;
        RECT 293.640 40.640 295.690 40.890 ;
        RECT 291.950 40.450 293.000 40.530 ;
        RECT 293.630 40.450 295.260 40.470 ;
        RECT 291.950 40.280 295.260 40.450 ;
        RECT 292.955 40.250 295.260 40.280 ;
        RECT 295.430 40.410 295.690 40.640 ;
        RECT 295.860 40.580 296.050 41.060 ;
        RECT 296.220 40.410 296.550 40.890 ;
        RECT 289.920 39.820 290.175 40.150 ;
        RECT 290.005 39.610 290.175 39.820 ;
        RECT 290.455 39.790 290.810 40.160 ;
        RECT 291.445 40.110 291.755 40.150 ;
        RECT 291.445 39.730 292.785 40.110 ;
        RECT 289.580 38.680 289.835 39.585 ;
        RECT 290.005 39.440 290.720 39.610 ;
        RECT 290.005 38.510 290.335 39.270 ;
        RECT 290.550 38.680 290.720 39.440 ;
        RECT 290.980 38.510 291.270 39.675 ;
        RECT 292.955 39.560 293.235 40.250 ;
        RECT 295.430 40.240 296.550 40.410 ;
        RECT 296.720 40.260 296.980 41.060 ;
        RECT 297.420 40.290 299.090 41.060 ;
        RECT 299.725 40.350 299.980 40.880 ;
        RECT 300.150 40.600 300.455 41.060 ;
        RECT 300.700 40.680 301.770 40.850 ;
        RECT 291.935 39.440 293.235 39.560 ;
        RECT 293.405 39.665 293.750 40.080 ;
        RECT 293.920 39.835 295.355 40.080 ;
        RECT 295.580 39.665 296.825 40.070 ;
        RECT 297.420 39.770 298.170 40.290 ;
        RECT 293.405 39.440 296.825 39.665 ;
        RECT 298.340 39.600 299.090 40.120 ;
        RECT 291.535 38.930 291.730 39.350 ;
        RECT 291.935 39.110 293.100 39.440 ;
        RECT 293.270 39.040 296.980 39.270 ;
        RECT 293.270 38.940 293.470 39.040 ;
        RECT 292.310 38.930 293.470 38.940 ;
        RECT 291.535 38.680 293.470 38.930 ;
        RECT 293.640 38.510 293.970 38.870 ;
        RECT 294.140 38.680 294.330 39.040 ;
        RECT 294.500 38.510 294.830 38.870 ;
        RECT 295.000 38.680 295.190 39.040 ;
        RECT 295.360 38.510 295.690 38.870 ;
        RECT 295.860 38.680 296.040 39.040 ;
        RECT 296.220 38.510 296.550 38.870 ;
        RECT 296.720 38.680 296.980 39.040 ;
        RECT 297.420 38.510 299.090 39.600 ;
        RECT 299.725 39.700 299.935 40.350 ;
        RECT 300.700 40.325 301.020 40.680 ;
        RECT 300.695 40.150 301.020 40.325 ;
        RECT 300.105 39.850 301.020 40.150 ;
        RECT 301.190 40.110 301.430 40.510 ;
        RECT 301.600 40.450 301.770 40.680 ;
        RECT 301.940 40.620 302.130 41.060 ;
        RECT 302.300 40.610 303.250 40.890 ;
        RECT 303.470 40.700 303.820 40.870 ;
        RECT 301.600 40.280 302.130 40.450 ;
        RECT 300.105 39.820 300.845 39.850 ;
        RECT 299.725 38.820 299.980 39.700 ;
        RECT 300.150 38.510 300.455 39.650 ;
        RECT 300.675 39.230 300.845 39.820 ;
        RECT 301.190 39.740 301.730 40.110 ;
        RECT 301.910 40.000 302.130 40.280 ;
        RECT 302.300 39.830 302.470 40.610 ;
        RECT 302.065 39.660 302.470 39.830 ;
        RECT 302.640 39.820 302.990 40.440 ;
        RECT 302.065 39.570 302.235 39.660 ;
        RECT 303.160 39.650 303.370 40.440 ;
        RECT 301.015 39.400 302.235 39.570 ;
        RECT 302.695 39.490 303.370 39.650 ;
        RECT 300.675 39.060 301.475 39.230 ;
        RECT 300.795 38.510 301.125 38.890 ;
        RECT 301.305 38.770 301.475 39.060 ;
        RECT 302.065 39.020 302.235 39.400 ;
        RECT 302.405 39.480 303.370 39.490 ;
        RECT 303.560 40.310 303.820 40.700 ;
        RECT 304.030 40.600 304.360 41.060 ;
        RECT 305.235 40.670 306.090 40.840 ;
        RECT 306.295 40.670 306.790 40.840 ;
        RECT 306.960 40.700 307.290 41.060 ;
        RECT 303.560 39.620 303.730 40.310 ;
        RECT 303.900 39.960 304.070 40.140 ;
        RECT 304.240 40.130 305.030 40.380 ;
        RECT 305.235 39.960 305.405 40.670 ;
        RECT 305.575 40.160 305.930 40.380 ;
        RECT 303.900 39.790 305.590 39.960 ;
        RECT 302.405 39.190 302.865 39.480 ;
        RECT 303.560 39.450 305.060 39.620 ;
        RECT 303.560 39.310 303.730 39.450 ;
        RECT 303.170 39.140 303.730 39.310 ;
        RECT 301.645 38.510 301.895 38.970 ;
        RECT 302.065 38.680 302.935 39.020 ;
        RECT 303.170 38.680 303.340 39.140 ;
        RECT 304.175 39.110 305.250 39.280 ;
        RECT 303.510 38.510 303.880 38.970 ;
        RECT 304.175 38.770 304.345 39.110 ;
        RECT 304.515 38.510 304.845 38.940 ;
        RECT 305.080 38.770 305.250 39.110 ;
        RECT 305.420 39.010 305.590 39.790 ;
        RECT 305.760 39.570 305.930 40.160 ;
        RECT 306.100 39.760 306.450 40.380 ;
        RECT 305.760 39.180 306.225 39.570 ;
        RECT 306.620 39.310 306.790 40.670 ;
        RECT 306.960 39.480 307.420 40.530 ;
        RECT 306.395 39.140 306.790 39.310 ;
        RECT 306.395 39.010 306.565 39.140 ;
        RECT 305.420 38.680 306.100 39.010 ;
        RECT 306.315 38.680 306.565 39.010 ;
        RECT 306.735 38.510 306.985 38.970 ;
        RECT 307.155 38.695 307.480 39.480 ;
        RECT 307.650 38.680 307.820 40.800 ;
        RECT 307.990 40.680 308.320 41.060 ;
        RECT 308.490 40.510 308.745 40.800 ;
        RECT 307.995 40.340 308.745 40.510 ;
        RECT 307.995 39.350 308.225 40.340 ;
        RECT 309.840 40.310 311.050 41.060 ;
        RECT 308.395 39.520 308.745 40.170 ;
        RECT 309.840 39.600 310.360 40.140 ;
        RECT 310.530 39.770 311.050 40.310 ;
        RECT 307.995 39.180 308.745 39.350 ;
        RECT 307.990 38.510 308.320 39.010 ;
        RECT 308.490 38.680 308.745 39.180 ;
        RECT 309.840 38.510 311.050 39.600 ;
        RECT 162.095 38.340 311.135 38.510 ;
        RECT 162.180 37.250 163.390 38.340 ;
        RECT 163.560 37.250 165.230 38.340 ;
        RECT 165.865 37.670 166.120 38.170 ;
        RECT 166.290 37.840 166.620 38.340 ;
        RECT 165.865 37.500 166.615 37.670 ;
        RECT 162.180 36.540 162.700 37.080 ;
        RECT 162.870 36.710 163.390 37.250 ;
        RECT 163.560 36.560 164.310 37.080 ;
        RECT 164.480 36.730 165.230 37.250 ;
        RECT 165.865 36.680 166.215 37.330 ;
        RECT 162.180 35.790 163.390 36.540 ;
        RECT 163.560 35.790 165.230 36.560 ;
        RECT 166.385 36.510 166.615 37.500 ;
        RECT 165.865 36.340 166.615 36.510 ;
        RECT 165.865 36.050 166.120 36.340 ;
        RECT 166.290 35.790 166.620 36.170 ;
        RECT 166.790 36.050 166.960 38.170 ;
        RECT 167.130 37.370 167.455 38.155 ;
        RECT 167.625 37.880 167.875 38.340 ;
        RECT 168.045 37.840 168.295 38.170 ;
        RECT 168.510 37.840 169.190 38.170 ;
        RECT 168.045 37.710 168.215 37.840 ;
        RECT 167.820 37.540 168.215 37.710 ;
        RECT 167.190 36.320 167.650 37.370 ;
        RECT 167.820 36.180 167.990 37.540 ;
        RECT 168.385 37.280 168.850 37.670 ;
        RECT 168.160 36.470 168.510 37.090 ;
        RECT 168.680 36.690 168.850 37.280 ;
        RECT 169.020 37.060 169.190 37.840 ;
        RECT 169.360 37.740 169.530 38.080 ;
        RECT 169.765 37.910 170.095 38.340 ;
        RECT 170.265 37.740 170.435 38.080 ;
        RECT 170.730 37.880 171.100 38.340 ;
        RECT 169.360 37.570 170.435 37.740 ;
        RECT 171.270 37.710 171.440 38.170 ;
        RECT 171.675 37.830 172.545 38.170 ;
        RECT 172.715 37.880 172.965 38.340 ;
        RECT 170.880 37.540 171.440 37.710 ;
        RECT 170.880 37.400 171.050 37.540 ;
        RECT 169.550 37.230 171.050 37.400 ;
        RECT 171.745 37.370 172.205 37.660 ;
        RECT 169.020 36.890 170.710 37.060 ;
        RECT 168.680 36.470 169.035 36.690 ;
        RECT 169.205 36.180 169.375 36.890 ;
        RECT 169.580 36.470 170.370 36.720 ;
        RECT 170.540 36.710 170.710 36.890 ;
        RECT 170.880 36.540 171.050 37.230 ;
        RECT 167.320 35.790 167.650 36.150 ;
        RECT 167.820 36.010 168.315 36.180 ;
        RECT 168.520 36.010 169.375 36.180 ;
        RECT 170.250 35.790 170.580 36.250 ;
        RECT 170.790 36.150 171.050 36.540 ;
        RECT 171.240 37.360 172.205 37.370 ;
        RECT 172.375 37.450 172.545 37.830 ;
        RECT 173.135 37.790 173.305 38.080 ;
        RECT 173.485 37.960 173.815 38.340 ;
        RECT 173.135 37.620 173.935 37.790 ;
        RECT 171.240 37.200 171.915 37.360 ;
        RECT 172.375 37.280 173.595 37.450 ;
        RECT 171.240 36.410 171.450 37.200 ;
        RECT 172.375 37.190 172.545 37.280 ;
        RECT 171.620 36.410 171.970 37.030 ;
        RECT 172.140 37.020 172.545 37.190 ;
        RECT 172.140 36.240 172.310 37.020 ;
        RECT 172.480 36.570 172.700 36.850 ;
        RECT 172.880 36.740 173.420 37.110 ;
        RECT 173.765 37.030 173.935 37.620 ;
        RECT 174.155 37.200 174.460 38.340 ;
        RECT 174.630 37.150 174.885 38.030 ;
        RECT 175.060 37.175 175.350 38.340 ;
        RECT 176.440 37.580 176.955 37.990 ;
        RECT 177.190 37.580 177.360 38.340 ;
        RECT 177.530 38.000 179.560 38.170 ;
        RECT 173.765 37.000 174.505 37.030 ;
        RECT 172.480 36.400 173.010 36.570 ;
        RECT 170.790 35.980 171.140 36.150 ;
        RECT 171.360 35.960 172.310 36.240 ;
        RECT 172.480 35.790 172.670 36.230 ;
        RECT 172.840 36.170 173.010 36.400 ;
        RECT 173.180 36.340 173.420 36.740 ;
        RECT 173.590 36.700 174.505 37.000 ;
        RECT 173.590 36.525 173.915 36.700 ;
        RECT 173.590 36.170 173.910 36.525 ;
        RECT 174.675 36.500 174.885 37.150 ;
        RECT 176.440 36.770 176.780 37.580 ;
        RECT 177.530 37.335 177.700 38.000 ;
        RECT 178.095 37.660 179.220 37.830 ;
        RECT 176.950 37.145 177.700 37.335 ;
        RECT 177.870 37.320 178.880 37.490 ;
        RECT 176.440 36.600 177.670 36.770 ;
        RECT 172.840 36.000 173.910 36.170 ;
        RECT 174.155 35.790 174.460 36.250 ;
        RECT 174.630 35.970 174.885 36.500 ;
        RECT 175.060 35.790 175.350 36.515 ;
        RECT 176.715 35.995 176.960 36.600 ;
        RECT 177.180 35.790 177.690 36.325 ;
        RECT 177.870 35.960 178.060 37.320 ;
        RECT 178.230 36.640 178.505 37.120 ;
        RECT 178.230 36.470 178.510 36.640 ;
        RECT 178.710 36.520 178.880 37.320 ;
        RECT 179.050 36.530 179.220 37.660 ;
        RECT 179.390 37.030 179.560 38.000 ;
        RECT 179.730 37.200 179.900 38.340 ;
        RECT 180.070 37.200 180.405 38.170 ;
        RECT 179.390 36.700 179.585 37.030 ;
        RECT 179.810 36.700 180.065 37.030 ;
        RECT 179.810 36.530 179.980 36.700 ;
        RECT 180.235 36.530 180.405 37.200 ;
        RECT 178.230 35.960 178.505 36.470 ;
        RECT 179.050 36.360 179.980 36.530 ;
        RECT 179.050 36.325 179.225 36.360 ;
        RECT 178.695 35.960 179.225 36.325 ;
        RECT 179.650 35.790 179.980 36.190 ;
        RECT 180.150 35.960 180.405 36.530 ;
        RECT 180.580 37.200 180.965 38.170 ;
        RECT 181.135 37.880 181.460 38.340 ;
        RECT 181.980 37.710 182.260 38.170 ;
        RECT 181.135 37.490 182.260 37.710 ;
        RECT 180.580 36.530 180.860 37.200 ;
        RECT 181.135 37.030 181.585 37.490 ;
        RECT 182.450 37.320 182.850 38.170 ;
        RECT 183.250 37.880 183.520 38.340 ;
        RECT 183.690 37.710 183.975 38.170 ;
        RECT 181.030 36.700 181.585 37.030 ;
        RECT 181.755 36.760 182.850 37.320 ;
        RECT 181.135 36.590 181.585 36.700 ;
        RECT 180.580 35.960 180.965 36.530 ;
        RECT 181.135 36.420 182.260 36.590 ;
        RECT 181.135 35.790 181.460 36.250 ;
        RECT 181.980 35.960 182.260 36.420 ;
        RECT 182.450 35.960 182.850 36.760 ;
        RECT 183.020 37.490 183.975 37.710 ;
        RECT 183.020 36.590 183.230 37.490 ;
        RECT 183.400 36.760 184.090 37.320 ;
        RECT 184.260 37.250 186.850 38.340 ;
        RECT 187.025 37.670 187.280 38.170 ;
        RECT 187.450 37.840 187.780 38.340 ;
        RECT 187.025 37.500 187.775 37.670 ;
        RECT 183.020 36.420 183.975 36.590 ;
        RECT 183.250 35.790 183.520 36.250 ;
        RECT 183.690 35.960 183.975 36.420 ;
        RECT 184.260 36.560 185.470 37.080 ;
        RECT 185.640 36.730 186.850 37.250 ;
        RECT 187.025 36.680 187.375 37.330 ;
        RECT 184.260 35.790 186.850 36.560 ;
        RECT 187.545 36.510 187.775 37.500 ;
        RECT 187.025 36.340 187.775 36.510 ;
        RECT 187.025 36.050 187.280 36.340 ;
        RECT 187.450 35.790 187.780 36.170 ;
        RECT 187.950 36.050 188.120 38.170 ;
        RECT 188.290 37.370 188.615 38.155 ;
        RECT 188.785 37.880 189.035 38.340 ;
        RECT 189.205 37.840 189.455 38.170 ;
        RECT 189.670 37.840 190.350 38.170 ;
        RECT 189.205 37.710 189.375 37.840 ;
        RECT 188.980 37.540 189.375 37.710 ;
        RECT 188.350 36.320 188.810 37.370 ;
        RECT 188.980 36.180 189.150 37.540 ;
        RECT 189.545 37.280 190.010 37.670 ;
        RECT 189.320 36.470 189.670 37.090 ;
        RECT 189.840 36.690 190.010 37.280 ;
        RECT 190.180 37.060 190.350 37.840 ;
        RECT 190.520 37.740 190.690 38.080 ;
        RECT 190.925 37.910 191.255 38.340 ;
        RECT 191.425 37.740 191.595 38.080 ;
        RECT 191.890 37.880 192.260 38.340 ;
        RECT 190.520 37.570 191.595 37.740 ;
        RECT 192.430 37.710 192.600 38.170 ;
        RECT 192.835 37.830 193.705 38.170 ;
        RECT 193.875 37.880 194.125 38.340 ;
        RECT 192.040 37.540 192.600 37.710 ;
        RECT 192.040 37.400 192.210 37.540 ;
        RECT 190.710 37.230 192.210 37.400 ;
        RECT 192.905 37.370 193.365 37.660 ;
        RECT 190.180 36.890 191.870 37.060 ;
        RECT 189.840 36.470 190.195 36.690 ;
        RECT 190.365 36.180 190.535 36.890 ;
        RECT 190.740 36.470 191.530 36.720 ;
        RECT 191.700 36.710 191.870 36.890 ;
        RECT 192.040 36.540 192.210 37.230 ;
        RECT 188.480 35.790 188.810 36.150 ;
        RECT 188.980 36.010 189.475 36.180 ;
        RECT 189.680 36.010 190.535 36.180 ;
        RECT 191.410 35.790 191.740 36.250 ;
        RECT 191.950 36.150 192.210 36.540 ;
        RECT 192.400 37.360 193.365 37.370 ;
        RECT 193.535 37.450 193.705 37.830 ;
        RECT 194.295 37.790 194.465 38.080 ;
        RECT 194.645 37.960 194.975 38.340 ;
        RECT 194.295 37.620 195.095 37.790 ;
        RECT 192.400 37.200 193.075 37.360 ;
        RECT 193.535 37.280 194.755 37.450 ;
        RECT 192.400 36.410 192.610 37.200 ;
        RECT 193.535 37.190 193.705 37.280 ;
        RECT 192.780 36.410 193.130 37.030 ;
        RECT 193.300 37.020 193.705 37.190 ;
        RECT 193.300 36.240 193.470 37.020 ;
        RECT 193.640 36.570 193.860 36.850 ;
        RECT 194.040 36.740 194.580 37.110 ;
        RECT 194.925 37.030 195.095 37.620 ;
        RECT 195.315 37.200 195.620 38.340 ;
        RECT 195.790 37.150 196.045 38.030 ;
        RECT 194.925 37.000 195.665 37.030 ;
        RECT 193.640 36.400 194.170 36.570 ;
        RECT 191.950 35.980 192.300 36.150 ;
        RECT 192.520 35.960 193.470 36.240 ;
        RECT 193.640 35.790 193.830 36.230 ;
        RECT 194.000 36.170 194.170 36.400 ;
        RECT 194.340 36.340 194.580 36.740 ;
        RECT 194.750 36.700 195.665 37.000 ;
        RECT 194.750 36.525 195.075 36.700 ;
        RECT 194.750 36.170 195.070 36.525 ;
        RECT 195.835 36.500 196.045 37.150 ;
        RECT 194.000 36.000 195.070 36.170 ;
        RECT 195.315 35.790 195.620 36.250 ;
        RECT 195.790 35.970 196.045 36.500 ;
        RECT 197.140 37.200 197.525 38.170 ;
        RECT 197.695 37.880 198.020 38.340 ;
        RECT 198.540 37.710 198.820 38.170 ;
        RECT 197.695 37.490 198.820 37.710 ;
        RECT 197.140 36.530 197.420 37.200 ;
        RECT 197.695 37.030 198.145 37.490 ;
        RECT 199.010 37.320 199.410 38.170 ;
        RECT 199.810 37.880 200.080 38.340 ;
        RECT 200.250 37.710 200.535 38.170 ;
        RECT 197.590 36.700 198.145 37.030 ;
        RECT 198.315 36.760 199.410 37.320 ;
        RECT 197.695 36.590 198.145 36.700 ;
        RECT 197.140 35.960 197.525 36.530 ;
        RECT 197.695 36.420 198.820 36.590 ;
        RECT 197.695 35.790 198.020 36.250 ;
        RECT 198.540 35.960 198.820 36.420 ;
        RECT 199.010 35.960 199.410 36.760 ;
        RECT 199.580 37.490 200.535 37.710 ;
        RECT 199.580 36.590 199.790 37.490 ;
        RECT 199.960 36.760 200.650 37.320 ;
        RECT 200.820 37.175 201.110 38.340 ;
        RECT 201.280 37.250 204.790 38.340 ;
        RECT 205.885 37.670 206.140 38.170 ;
        RECT 206.310 37.840 206.640 38.340 ;
        RECT 205.885 37.500 206.635 37.670 ;
        RECT 199.580 36.420 200.535 36.590 ;
        RECT 201.280 36.560 202.930 37.080 ;
        RECT 203.100 36.730 204.790 37.250 ;
        RECT 205.885 36.680 206.235 37.330 ;
        RECT 199.810 35.790 200.080 36.250 ;
        RECT 200.250 35.960 200.535 36.420 ;
        RECT 200.820 35.790 201.110 36.515 ;
        RECT 201.280 35.790 204.790 36.560 ;
        RECT 206.405 36.510 206.635 37.500 ;
        RECT 205.885 36.340 206.635 36.510 ;
        RECT 205.885 36.050 206.140 36.340 ;
        RECT 206.310 35.790 206.640 36.170 ;
        RECT 206.810 36.050 206.980 38.170 ;
        RECT 207.150 37.370 207.475 38.155 ;
        RECT 207.645 37.880 207.895 38.340 ;
        RECT 208.065 37.840 208.315 38.170 ;
        RECT 208.530 37.840 209.210 38.170 ;
        RECT 208.065 37.710 208.235 37.840 ;
        RECT 207.840 37.540 208.235 37.710 ;
        RECT 207.210 36.320 207.670 37.370 ;
        RECT 207.840 36.180 208.010 37.540 ;
        RECT 208.405 37.280 208.870 37.670 ;
        RECT 208.180 36.470 208.530 37.090 ;
        RECT 208.700 36.690 208.870 37.280 ;
        RECT 209.040 37.060 209.210 37.840 ;
        RECT 209.380 37.740 209.550 38.080 ;
        RECT 209.785 37.910 210.115 38.340 ;
        RECT 210.285 37.740 210.455 38.080 ;
        RECT 210.750 37.880 211.120 38.340 ;
        RECT 209.380 37.570 210.455 37.740 ;
        RECT 211.290 37.710 211.460 38.170 ;
        RECT 211.695 37.830 212.565 38.170 ;
        RECT 212.735 37.880 212.985 38.340 ;
        RECT 210.900 37.540 211.460 37.710 ;
        RECT 210.900 37.400 211.070 37.540 ;
        RECT 209.570 37.230 211.070 37.400 ;
        RECT 211.765 37.370 212.225 37.660 ;
        RECT 209.040 36.890 210.730 37.060 ;
        RECT 208.700 36.470 209.055 36.690 ;
        RECT 209.225 36.180 209.395 36.890 ;
        RECT 209.600 36.470 210.390 36.720 ;
        RECT 210.560 36.710 210.730 36.890 ;
        RECT 210.900 36.540 211.070 37.230 ;
        RECT 207.340 35.790 207.670 36.150 ;
        RECT 207.840 36.010 208.335 36.180 ;
        RECT 208.540 36.010 209.395 36.180 ;
        RECT 210.270 35.790 210.600 36.250 ;
        RECT 210.810 36.150 211.070 36.540 ;
        RECT 211.260 37.360 212.225 37.370 ;
        RECT 212.395 37.450 212.565 37.830 ;
        RECT 213.155 37.790 213.325 38.080 ;
        RECT 213.505 37.960 213.835 38.340 ;
        RECT 213.155 37.620 213.955 37.790 ;
        RECT 211.260 37.200 211.935 37.360 ;
        RECT 212.395 37.280 213.615 37.450 ;
        RECT 211.260 36.410 211.470 37.200 ;
        RECT 212.395 37.190 212.565 37.280 ;
        RECT 211.640 36.410 211.990 37.030 ;
        RECT 212.160 37.020 212.565 37.190 ;
        RECT 212.160 36.240 212.330 37.020 ;
        RECT 212.500 36.570 212.720 36.850 ;
        RECT 212.900 36.740 213.440 37.110 ;
        RECT 213.785 37.030 213.955 37.620 ;
        RECT 214.175 37.200 214.480 38.340 ;
        RECT 214.650 37.150 214.905 38.030 ;
        RECT 215.080 37.905 220.425 38.340 ;
        RECT 213.785 37.000 214.525 37.030 ;
        RECT 212.500 36.400 213.030 36.570 ;
        RECT 210.810 35.980 211.160 36.150 ;
        RECT 211.380 35.960 212.330 36.240 ;
        RECT 212.500 35.790 212.690 36.230 ;
        RECT 212.860 36.170 213.030 36.400 ;
        RECT 213.200 36.340 213.440 36.740 ;
        RECT 213.610 36.700 214.525 37.000 ;
        RECT 213.610 36.525 213.935 36.700 ;
        RECT 213.610 36.170 213.930 36.525 ;
        RECT 214.695 36.500 214.905 37.150 ;
        RECT 212.860 36.000 213.930 36.170 ;
        RECT 214.175 35.790 214.480 36.250 ;
        RECT 214.650 35.970 214.905 36.500 ;
        RECT 216.665 36.335 217.005 37.165 ;
        RECT 218.485 36.655 218.835 37.905 ;
        RECT 220.600 37.265 220.870 38.170 ;
        RECT 221.040 37.580 221.370 38.340 ;
        RECT 221.550 37.410 221.720 38.170 ;
        RECT 220.600 36.465 220.770 37.265 ;
        RECT 221.055 37.240 221.720 37.410 ;
        RECT 221.055 37.095 221.225 37.240 ;
        RECT 220.940 36.765 221.225 37.095 ;
        RECT 221.980 37.200 222.365 38.170 ;
        RECT 222.535 37.880 222.860 38.340 ;
        RECT 223.380 37.710 223.660 38.170 ;
        RECT 222.535 37.490 223.660 37.710 ;
        RECT 221.055 36.510 221.225 36.765 ;
        RECT 221.460 36.690 221.790 37.060 ;
        RECT 221.980 36.530 222.260 37.200 ;
        RECT 222.535 37.030 222.985 37.490 ;
        RECT 223.850 37.320 224.250 38.170 ;
        RECT 224.650 37.880 224.920 38.340 ;
        RECT 225.090 37.710 225.375 38.170 ;
        RECT 222.430 36.700 222.985 37.030 ;
        RECT 223.155 36.760 224.250 37.320 ;
        RECT 222.535 36.590 222.985 36.700 ;
        RECT 215.080 35.790 220.425 36.335 ;
        RECT 220.600 35.960 220.860 36.465 ;
        RECT 221.055 36.340 221.720 36.510 ;
        RECT 221.040 35.790 221.370 36.170 ;
        RECT 221.550 35.960 221.720 36.340 ;
        RECT 221.980 35.960 222.365 36.530 ;
        RECT 222.535 36.420 223.660 36.590 ;
        RECT 222.535 35.790 222.860 36.250 ;
        RECT 223.380 35.960 223.660 36.420 ;
        RECT 223.850 35.960 224.250 36.760 ;
        RECT 224.420 37.490 225.375 37.710 ;
        RECT 224.420 36.590 224.630 37.490 ;
        RECT 224.800 36.760 225.490 37.320 ;
        RECT 226.580 37.175 226.870 38.340 ;
        RECT 227.040 37.200 227.425 38.170 ;
        RECT 227.595 37.880 227.920 38.340 ;
        RECT 228.440 37.710 228.720 38.170 ;
        RECT 227.595 37.490 228.720 37.710 ;
        RECT 224.420 36.420 225.375 36.590 ;
        RECT 227.040 36.530 227.320 37.200 ;
        RECT 227.595 37.030 228.045 37.490 ;
        RECT 228.910 37.320 229.310 38.170 ;
        RECT 229.710 37.880 229.980 38.340 ;
        RECT 230.150 37.710 230.435 38.170 ;
        RECT 227.490 36.700 228.045 37.030 ;
        RECT 228.215 36.760 229.310 37.320 ;
        RECT 227.595 36.590 228.045 36.700 ;
        RECT 224.650 35.790 224.920 36.250 ;
        RECT 225.090 35.960 225.375 36.420 ;
        RECT 226.580 35.790 226.870 36.515 ;
        RECT 227.040 35.960 227.425 36.530 ;
        RECT 227.595 36.420 228.720 36.590 ;
        RECT 227.595 35.790 227.920 36.250 ;
        RECT 228.440 35.960 228.720 36.420 ;
        RECT 228.910 35.960 229.310 36.760 ;
        RECT 229.480 37.490 230.435 37.710 ;
        RECT 229.480 36.590 229.690 37.490 ;
        RECT 229.860 36.760 230.550 37.320 ;
        RECT 230.725 37.200 231.060 38.170 ;
        RECT 231.230 37.200 231.400 38.340 ;
        RECT 231.570 38.000 233.600 38.170 ;
        RECT 229.480 36.420 230.435 36.590 ;
        RECT 229.710 35.790 229.980 36.250 ;
        RECT 230.150 35.960 230.435 36.420 ;
        RECT 230.725 36.530 230.895 37.200 ;
        RECT 231.570 37.030 231.740 38.000 ;
        RECT 231.065 36.700 231.320 37.030 ;
        RECT 231.545 36.700 231.740 37.030 ;
        RECT 231.910 37.660 233.035 37.830 ;
        RECT 231.150 36.530 231.320 36.700 ;
        RECT 231.910 36.530 232.080 37.660 ;
        RECT 230.725 35.960 230.980 36.530 ;
        RECT 231.150 36.360 232.080 36.530 ;
        RECT 232.250 37.320 233.260 37.490 ;
        RECT 232.250 36.520 232.420 37.320 ;
        RECT 232.625 36.980 232.900 37.120 ;
        RECT 232.620 36.810 232.900 36.980 ;
        RECT 231.905 36.325 232.080 36.360 ;
        RECT 231.150 35.790 231.480 36.190 ;
        RECT 231.905 35.960 232.435 36.325 ;
        RECT 232.625 35.960 232.900 36.810 ;
        RECT 233.070 35.960 233.260 37.320 ;
        RECT 233.430 37.335 233.600 38.000 ;
        RECT 233.770 37.580 233.940 38.340 ;
        RECT 234.175 37.580 234.690 37.990 ;
        RECT 233.430 37.145 234.180 37.335 ;
        RECT 234.350 36.770 234.690 37.580 ;
        RECT 233.460 36.600 234.690 36.770 ;
        RECT 233.440 35.790 233.950 36.325 ;
        RECT 234.170 35.995 234.415 36.600 ;
        RECT 235.780 35.960 236.530 38.170 ;
        RECT 237.625 37.915 237.960 38.340 ;
        RECT 238.130 37.735 238.315 38.140 ;
        RECT 237.650 37.560 238.315 37.735 ;
        RECT 238.520 37.560 238.850 38.340 ;
        RECT 237.650 36.530 237.990 37.560 ;
        RECT 239.020 37.370 239.290 38.140 ;
        RECT 238.160 37.200 239.290 37.370 ;
        RECT 238.160 36.700 238.410 37.200 ;
        RECT 237.650 36.360 238.335 36.530 ;
        RECT 238.590 36.450 238.950 37.030 ;
        RECT 237.625 35.790 237.960 36.190 ;
        RECT 238.130 35.960 238.335 36.360 ;
        RECT 239.120 36.290 239.290 37.200 ;
        RECT 238.545 35.790 238.820 36.270 ;
        RECT 239.030 35.960 239.290 36.290 ;
        RECT 240.380 35.960 241.130 38.170 ;
        RECT 241.305 37.150 241.560 38.030 ;
        RECT 241.730 37.200 242.035 38.340 ;
        RECT 242.375 37.960 242.705 38.340 ;
        RECT 242.885 37.790 243.055 38.080 ;
        RECT 243.225 37.880 243.475 38.340 ;
        RECT 242.255 37.620 243.055 37.790 ;
        RECT 243.645 37.830 244.515 38.170 ;
        RECT 241.305 36.500 241.515 37.150 ;
        RECT 242.255 37.030 242.425 37.620 ;
        RECT 243.645 37.450 243.815 37.830 ;
        RECT 244.750 37.710 244.920 38.170 ;
        RECT 245.090 37.880 245.460 38.340 ;
        RECT 245.755 37.740 245.925 38.080 ;
        RECT 246.095 37.910 246.425 38.340 ;
        RECT 246.660 37.740 246.830 38.080 ;
        RECT 242.595 37.280 243.815 37.450 ;
        RECT 243.985 37.370 244.445 37.660 ;
        RECT 244.750 37.540 245.310 37.710 ;
        RECT 245.755 37.570 246.830 37.740 ;
        RECT 247.000 37.840 247.680 38.170 ;
        RECT 247.895 37.840 248.145 38.170 ;
        RECT 248.315 37.880 248.565 38.340 ;
        RECT 245.140 37.400 245.310 37.540 ;
        RECT 243.985 37.360 244.950 37.370 ;
        RECT 243.645 37.190 243.815 37.280 ;
        RECT 244.275 37.200 244.950 37.360 ;
        RECT 241.685 37.000 242.425 37.030 ;
        RECT 241.685 36.700 242.600 37.000 ;
        RECT 242.275 36.525 242.600 36.700 ;
        RECT 241.305 35.970 241.560 36.500 ;
        RECT 241.730 35.790 242.035 36.250 ;
        RECT 242.280 36.170 242.600 36.525 ;
        RECT 242.770 36.740 243.310 37.110 ;
        RECT 243.645 37.020 244.050 37.190 ;
        RECT 242.770 36.340 243.010 36.740 ;
        RECT 243.490 36.570 243.710 36.850 ;
        RECT 243.180 36.400 243.710 36.570 ;
        RECT 243.180 36.170 243.350 36.400 ;
        RECT 243.880 36.240 244.050 37.020 ;
        RECT 244.220 36.410 244.570 37.030 ;
        RECT 244.740 36.410 244.950 37.200 ;
        RECT 245.140 37.230 246.640 37.400 ;
        RECT 245.140 36.540 245.310 37.230 ;
        RECT 247.000 37.060 247.170 37.840 ;
        RECT 247.975 37.710 248.145 37.840 ;
        RECT 245.480 36.890 247.170 37.060 ;
        RECT 247.340 37.280 247.805 37.670 ;
        RECT 247.975 37.540 248.370 37.710 ;
        RECT 245.480 36.710 245.650 36.890 ;
        RECT 242.280 36.000 243.350 36.170 ;
        RECT 243.520 35.790 243.710 36.230 ;
        RECT 243.880 35.960 244.830 36.240 ;
        RECT 245.140 36.150 245.400 36.540 ;
        RECT 245.820 36.470 246.610 36.720 ;
        RECT 245.050 35.980 245.400 36.150 ;
        RECT 245.610 35.790 245.940 36.250 ;
        RECT 246.815 36.180 246.985 36.890 ;
        RECT 247.340 36.690 247.510 37.280 ;
        RECT 247.155 36.470 247.510 36.690 ;
        RECT 247.680 36.470 248.030 37.090 ;
        RECT 248.200 36.180 248.370 37.540 ;
        RECT 248.735 37.370 249.060 38.155 ;
        RECT 248.540 36.320 249.000 37.370 ;
        RECT 246.815 36.010 247.670 36.180 ;
        RECT 247.875 36.010 248.370 36.180 ;
        RECT 248.540 35.790 248.870 36.150 ;
        RECT 249.230 36.050 249.400 38.170 ;
        RECT 249.570 37.840 249.900 38.340 ;
        RECT 250.070 37.670 250.325 38.170 ;
        RECT 249.575 37.500 250.325 37.670 ;
        RECT 249.575 36.510 249.805 37.500 ;
        RECT 249.975 36.680 250.325 37.330 ;
        RECT 250.500 37.250 252.170 38.340 ;
        RECT 250.500 36.560 251.250 37.080 ;
        RECT 251.420 36.730 252.170 37.250 ;
        RECT 252.340 37.175 252.630 38.340 ;
        RECT 252.800 37.250 254.010 38.340 ;
        RECT 249.575 36.340 250.325 36.510 ;
        RECT 249.570 35.790 249.900 36.170 ;
        RECT 250.070 36.050 250.325 36.340 ;
        RECT 250.500 35.790 252.170 36.560 ;
        RECT 252.800 36.540 253.320 37.080 ;
        RECT 253.490 36.710 254.010 37.250 ;
        RECT 254.185 37.150 254.440 38.030 ;
        RECT 254.610 37.200 254.915 38.340 ;
        RECT 255.255 37.960 255.585 38.340 ;
        RECT 255.765 37.790 255.935 38.080 ;
        RECT 256.105 37.880 256.355 38.340 ;
        RECT 255.135 37.620 255.935 37.790 ;
        RECT 256.525 37.830 257.395 38.170 ;
        RECT 252.340 35.790 252.630 36.515 ;
        RECT 252.800 35.790 254.010 36.540 ;
        RECT 254.185 36.500 254.395 37.150 ;
        RECT 255.135 37.030 255.305 37.620 ;
        RECT 256.525 37.450 256.695 37.830 ;
        RECT 257.630 37.710 257.800 38.170 ;
        RECT 257.970 37.880 258.340 38.340 ;
        RECT 258.635 37.740 258.805 38.080 ;
        RECT 258.975 37.910 259.305 38.340 ;
        RECT 259.540 37.740 259.710 38.080 ;
        RECT 255.475 37.280 256.695 37.450 ;
        RECT 256.865 37.370 257.325 37.660 ;
        RECT 257.630 37.540 258.190 37.710 ;
        RECT 258.635 37.570 259.710 37.740 ;
        RECT 259.880 37.840 260.560 38.170 ;
        RECT 260.775 37.840 261.025 38.170 ;
        RECT 261.195 37.880 261.445 38.340 ;
        RECT 258.020 37.400 258.190 37.540 ;
        RECT 256.865 37.360 257.830 37.370 ;
        RECT 256.525 37.190 256.695 37.280 ;
        RECT 257.155 37.200 257.830 37.360 ;
        RECT 254.565 37.000 255.305 37.030 ;
        RECT 254.565 36.700 255.480 37.000 ;
        RECT 255.155 36.525 255.480 36.700 ;
        RECT 254.185 35.970 254.440 36.500 ;
        RECT 254.610 35.790 254.915 36.250 ;
        RECT 255.160 36.170 255.480 36.525 ;
        RECT 255.650 36.740 256.190 37.110 ;
        RECT 256.525 37.020 256.930 37.190 ;
        RECT 255.650 36.340 255.890 36.740 ;
        RECT 256.370 36.570 256.590 36.850 ;
        RECT 256.060 36.400 256.590 36.570 ;
        RECT 256.060 36.170 256.230 36.400 ;
        RECT 256.760 36.240 256.930 37.020 ;
        RECT 257.100 36.410 257.450 37.030 ;
        RECT 257.620 36.410 257.830 37.200 ;
        RECT 258.020 37.230 259.520 37.400 ;
        RECT 258.020 36.540 258.190 37.230 ;
        RECT 259.880 37.060 260.050 37.840 ;
        RECT 260.855 37.710 261.025 37.840 ;
        RECT 258.360 36.890 260.050 37.060 ;
        RECT 260.220 37.280 260.685 37.670 ;
        RECT 260.855 37.540 261.250 37.710 ;
        RECT 258.360 36.710 258.530 36.890 ;
        RECT 255.160 36.000 256.230 36.170 ;
        RECT 256.400 35.790 256.590 36.230 ;
        RECT 256.760 35.960 257.710 36.240 ;
        RECT 258.020 36.150 258.280 36.540 ;
        RECT 258.700 36.470 259.490 36.720 ;
        RECT 257.930 35.980 258.280 36.150 ;
        RECT 258.490 35.790 258.820 36.250 ;
        RECT 259.695 36.180 259.865 36.890 ;
        RECT 260.220 36.690 260.390 37.280 ;
        RECT 260.035 36.470 260.390 36.690 ;
        RECT 260.560 36.470 260.910 37.090 ;
        RECT 261.080 36.180 261.250 37.540 ;
        RECT 261.615 37.370 261.940 38.155 ;
        RECT 261.420 36.320 261.880 37.370 ;
        RECT 259.695 36.010 260.550 36.180 ;
        RECT 260.755 36.010 261.250 36.180 ;
        RECT 261.420 35.790 261.750 36.150 ;
        RECT 262.110 36.050 262.280 38.170 ;
        RECT 262.450 37.840 262.780 38.340 ;
        RECT 262.950 37.670 263.205 38.170 ;
        RECT 262.455 37.500 263.205 37.670 ;
        RECT 262.455 36.510 262.685 37.500 ;
        RECT 262.855 36.680 263.205 37.330 ;
        RECT 263.380 37.250 265.970 38.340 ;
        RECT 263.380 36.560 264.590 37.080 ;
        RECT 264.760 36.730 265.970 37.250 ;
        RECT 266.230 37.410 266.400 38.170 ;
        RECT 266.580 37.580 266.910 38.340 ;
        RECT 266.230 37.240 266.895 37.410 ;
        RECT 267.080 37.265 267.350 38.170 ;
        RECT 266.725 37.095 266.895 37.240 ;
        RECT 266.160 36.690 266.490 37.060 ;
        RECT 266.725 36.765 267.010 37.095 ;
        RECT 262.455 36.340 263.205 36.510 ;
        RECT 262.450 35.790 262.780 36.170 ;
        RECT 262.950 36.050 263.205 36.340 ;
        RECT 263.380 35.790 265.970 36.560 ;
        RECT 266.725 36.510 266.895 36.765 ;
        RECT 266.230 36.340 266.895 36.510 ;
        RECT 267.180 36.465 267.350 37.265 ;
        RECT 266.230 35.960 266.400 36.340 ;
        RECT 266.580 35.790 266.910 36.170 ;
        RECT 267.090 35.960 267.350 36.465 ;
        RECT 267.520 37.200 267.905 38.170 ;
        RECT 268.075 37.880 268.400 38.340 ;
        RECT 268.920 37.710 269.200 38.170 ;
        RECT 268.075 37.490 269.200 37.710 ;
        RECT 267.520 36.530 267.800 37.200 ;
        RECT 268.075 37.030 268.525 37.490 ;
        RECT 269.390 37.320 269.790 38.170 ;
        RECT 270.190 37.880 270.460 38.340 ;
        RECT 270.630 37.710 270.915 38.170 ;
        RECT 267.970 36.700 268.525 37.030 ;
        RECT 268.695 36.760 269.790 37.320 ;
        RECT 268.075 36.590 268.525 36.700 ;
        RECT 267.520 35.960 267.905 36.530 ;
        RECT 268.075 36.420 269.200 36.590 ;
        RECT 268.075 35.790 268.400 36.250 ;
        RECT 268.920 35.960 269.200 36.420 ;
        RECT 269.390 35.960 269.790 36.760 ;
        RECT 269.960 37.490 270.915 37.710 ;
        RECT 269.960 36.590 270.170 37.490 ;
        RECT 270.340 36.760 271.030 37.320 ;
        RECT 271.200 37.200 271.585 38.170 ;
        RECT 271.755 37.880 272.080 38.340 ;
        RECT 272.600 37.710 272.880 38.170 ;
        RECT 271.755 37.490 272.880 37.710 ;
        RECT 269.960 36.420 270.915 36.590 ;
        RECT 270.190 35.790 270.460 36.250 ;
        RECT 270.630 35.960 270.915 36.420 ;
        RECT 271.200 36.530 271.480 37.200 ;
        RECT 271.755 37.030 272.205 37.490 ;
        RECT 273.070 37.320 273.470 38.170 ;
        RECT 273.870 37.880 274.140 38.340 ;
        RECT 274.310 37.710 274.595 38.170 ;
        RECT 271.650 36.700 272.205 37.030 ;
        RECT 272.375 36.760 273.470 37.320 ;
        RECT 271.755 36.590 272.205 36.700 ;
        RECT 271.200 35.960 271.585 36.530 ;
        RECT 271.755 36.420 272.880 36.590 ;
        RECT 271.755 35.790 272.080 36.250 ;
        RECT 272.600 35.960 272.880 36.420 ;
        RECT 273.070 35.960 273.470 36.760 ;
        RECT 273.640 37.490 274.595 37.710 ;
        RECT 273.640 36.590 273.850 37.490 ;
        RECT 274.900 37.450 275.160 38.160 ;
        RECT 275.330 37.630 275.660 38.340 ;
        RECT 275.830 37.450 276.060 38.160 ;
        RECT 274.020 36.760 274.710 37.320 ;
        RECT 274.900 37.210 276.060 37.450 ;
        RECT 276.240 37.430 276.510 38.160 ;
        RECT 276.690 37.610 277.030 38.340 ;
        RECT 276.240 37.210 277.010 37.430 ;
        RECT 274.890 36.700 275.190 37.030 ;
        RECT 275.370 36.720 275.895 37.030 ;
        RECT 276.075 36.720 276.540 37.030 ;
        RECT 273.640 36.420 274.595 36.590 ;
        RECT 273.870 35.790 274.140 36.250 ;
        RECT 274.310 35.960 274.595 36.420 ;
        RECT 274.900 35.790 275.190 36.520 ;
        RECT 275.370 36.080 275.600 36.720 ;
        RECT 276.720 36.540 277.010 37.210 ;
        RECT 275.780 36.340 277.010 36.540 ;
        RECT 275.780 35.970 276.090 36.340 ;
        RECT 276.270 35.790 276.940 36.160 ;
        RECT 277.200 35.970 277.460 38.160 ;
        RECT 278.100 37.175 278.390 38.340 ;
        RECT 279.665 37.370 280.055 37.545 ;
        RECT 280.540 37.540 280.870 38.340 ;
        RECT 281.040 37.550 281.575 38.170 ;
        RECT 279.665 37.200 281.090 37.370 ;
        RECT 278.100 35.790 278.390 36.515 ;
        RECT 279.540 36.470 279.895 37.030 ;
        RECT 280.065 36.300 280.235 37.200 ;
        RECT 280.405 36.470 280.670 37.030 ;
        RECT 280.920 36.700 281.090 37.200 ;
        RECT 281.260 36.530 281.575 37.550 ;
        RECT 282.250 37.390 282.525 38.160 ;
        RECT 282.695 37.730 283.025 38.160 ;
        RECT 283.195 37.900 283.390 38.340 ;
        RECT 283.570 37.730 283.900 38.160 ;
        RECT 282.695 37.560 283.900 37.730 ;
        RECT 282.250 37.200 282.835 37.390 ;
        RECT 283.005 37.230 283.900 37.560 ;
        RECT 284.080 37.470 284.355 38.170 ;
        RECT 284.525 37.795 284.780 38.340 ;
        RECT 284.950 37.830 285.430 38.170 ;
        RECT 285.605 37.785 286.210 38.340 ;
        RECT 285.595 37.685 286.210 37.785 ;
        RECT 285.595 37.660 285.780 37.685 ;
        RECT 279.645 35.790 279.885 36.300 ;
        RECT 280.065 35.970 280.345 36.300 ;
        RECT 280.575 35.790 280.790 36.300 ;
        RECT 280.960 35.960 281.575 36.530 ;
        RECT 282.250 36.380 282.490 37.030 ;
        RECT 282.660 36.530 282.835 37.200 ;
        RECT 283.005 36.700 283.420 37.030 ;
        RECT 283.600 36.700 283.895 37.030 ;
        RECT 282.660 36.350 282.990 36.530 ;
        RECT 282.265 35.790 282.595 36.180 ;
        RECT 282.765 35.970 282.990 36.350 ;
        RECT 283.190 36.080 283.420 36.700 ;
        RECT 283.600 35.790 283.900 36.520 ;
        RECT 284.080 36.440 284.250 37.470 ;
        RECT 284.525 37.340 285.280 37.590 ;
        RECT 285.450 37.415 285.780 37.660 ;
        RECT 286.385 37.670 286.640 38.170 ;
        RECT 286.810 37.840 287.140 38.340 ;
        RECT 284.525 37.305 285.295 37.340 ;
        RECT 284.525 37.295 285.310 37.305 ;
        RECT 284.420 37.280 285.315 37.295 ;
        RECT 284.420 37.265 285.335 37.280 ;
        RECT 284.420 37.255 285.355 37.265 ;
        RECT 284.420 37.245 285.380 37.255 ;
        RECT 284.420 37.215 285.450 37.245 ;
        RECT 284.420 37.185 285.470 37.215 ;
        RECT 284.420 37.155 285.490 37.185 ;
        RECT 284.420 37.130 285.520 37.155 ;
        RECT 284.420 37.095 285.555 37.130 ;
        RECT 284.420 37.090 285.585 37.095 ;
        RECT 284.420 36.695 284.650 37.090 ;
        RECT 285.195 37.085 285.585 37.090 ;
        RECT 285.220 37.075 285.585 37.085 ;
        RECT 285.235 37.070 285.585 37.075 ;
        RECT 285.250 37.065 285.585 37.070 ;
        RECT 285.950 37.065 286.210 37.515 ;
        RECT 286.385 37.500 287.135 37.670 ;
        RECT 285.250 37.060 286.210 37.065 ;
        RECT 285.260 37.050 286.210 37.060 ;
        RECT 285.270 37.045 286.210 37.050 ;
        RECT 285.280 37.035 286.210 37.045 ;
        RECT 285.285 37.025 286.210 37.035 ;
        RECT 285.290 37.020 286.210 37.025 ;
        RECT 285.300 37.005 286.210 37.020 ;
        RECT 285.305 36.990 286.210 37.005 ;
        RECT 285.315 36.965 286.210 36.990 ;
        RECT 284.820 36.495 285.150 36.920 ;
        RECT 284.080 35.960 284.340 36.440 ;
        RECT 284.510 35.790 284.760 36.330 ;
        RECT 284.930 36.010 285.150 36.495 ;
        RECT 285.320 36.895 286.210 36.965 ;
        RECT 285.320 36.170 285.490 36.895 ;
        RECT 285.660 36.340 286.210 36.725 ;
        RECT 286.385 36.680 286.735 37.330 ;
        RECT 286.905 36.510 287.135 37.500 ;
        RECT 286.385 36.340 287.135 36.510 ;
        RECT 285.320 36.000 286.210 36.170 ;
        RECT 286.385 36.050 286.640 36.340 ;
        RECT 286.810 35.790 287.140 36.170 ;
        RECT 287.310 36.050 287.480 38.170 ;
        RECT 287.650 37.370 287.975 38.155 ;
        RECT 288.145 37.880 288.395 38.340 ;
        RECT 288.565 37.840 288.815 38.170 ;
        RECT 289.030 37.840 289.710 38.170 ;
        RECT 288.565 37.710 288.735 37.840 ;
        RECT 288.340 37.540 288.735 37.710 ;
        RECT 287.710 36.320 288.170 37.370 ;
        RECT 288.340 36.180 288.510 37.540 ;
        RECT 288.905 37.280 289.370 37.670 ;
        RECT 288.680 36.470 289.030 37.090 ;
        RECT 289.200 36.690 289.370 37.280 ;
        RECT 289.540 37.060 289.710 37.840 ;
        RECT 289.880 37.740 290.050 38.080 ;
        RECT 290.285 37.910 290.615 38.340 ;
        RECT 290.785 37.740 290.955 38.080 ;
        RECT 291.250 37.880 291.620 38.340 ;
        RECT 289.880 37.570 290.955 37.740 ;
        RECT 291.790 37.710 291.960 38.170 ;
        RECT 292.195 37.830 293.065 38.170 ;
        RECT 293.235 37.880 293.485 38.340 ;
        RECT 291.400 37.540 291.960 37.710 ;
        RECT 291.400 37.400 291.570 37.540 ;
        RECT 290.070 37.230 291.570 37.400 ;
        RECT 292.265 37.370 292.725 37.660 ;
        RECT 289.540 36.890 291.230 37.060 ;
        RECT 289.200 36.470 289.555 36.690 ;
        RECT 289.725 36.180 289.895 36.890 ;
        RECT 290.100 36.470 290.890 36.720 ;
        RECT 291.060 36.710 291.230 36.890 ;
        RECT 291.400 36.540 291.570 37.230 ;
        RECT 287.840 35.790 288.170 36.150 ;
        RECT 288.340 36.010 288.835 36.180 ;
        RECT 289.040 36.010 289.895 36.180 ;
        RECT 290.770 35.790 291.100 36.250 ;
        RECT 291.310 36.150 291.570 36.540 ;
        RECT 291.760 37.360 292.725 37.370 ;
        RECT 292.895 37.450 293.065 37.830 ;
        RECT 293.655 37.790 293.825 38.080 ;
        RECT 294.005 37.960 294.335 38.340 ;
        RECT 293.655 37.620 294.455 37.790 ;
        RECT 291.760 37.200 292.435 37.360 ;
        RECT 292.895 37.280 294.115 37.450 ;
        RECT 291.760 36.410 291.970 37.200 ;
        RECT 292.895 37.190 293.065 37.280 ;
        RECT 292.140 36.410 292.490 37.030 ;
        RECT 292.660 37.020 293.065 37.190 ;
        RECT 292.660 36.240 292.830 37.020 ;
        RECT 293.000 36.570 293.220 36.850 ;
        RECT 293.400 36.740 293.940 37.110 ;
        RECT 294.285 37.030 294.455 37.620 ;
        RECT 294.675 37.200 294.980 38.340 ;
        RECT 295.150 37.150 295.405 38.030 ;
        RECT 294.285 37.000 295.025 37.030 ;
        RECT 293.000 36.400 293.530 36.570 ;
        RECT 291.310 35.980 291.660 36.150 ;
        RECT 291.880 35.960 292.830 36.240 ;
        RECT 293.000 35.790 293.190 36.230 ;
        RECT 293.360 36.170 293.530 36.400 ;
        RECT 293.700 36.340 293.940 36.740 ;
        RECT 294.110 36.700 295.025 37.000 ;
        RECT 294.110 36.525 294.435 36.700 ;
        RECT 294.110 36.170 294.430 36.525 ;
        RECT 295.195 36.500 295.405 37.150 ;
        RECT 293.360 36.000 294.430 36.170 ;
        RECT 294.675 35.790 294.980 36.250 ;
        RECT 295.150 35.970 295.405 36.500 ;
        RECT 295.580 37.470 295.855 38.170 ;
        RECT 296.025 37.795 296.280 38.340 ;
        RECT 296.450 37.830 296.930 38.170 ;
        RECT 297.105 37.785 297.710 38.340 ;
        RECT 297.095 37.685 297.710 37.785 ;
        RECT 297.095 37.660 297.280 37.685 ;
        RECT 295.580 36.440 295.750 37.470 ;
        RECT 296.025 37.340 296.780 37.590 ;
        RECT 296.950 37.415 297.280 37.660 ;
        RECT 296.025 37.305 296.795 37.340 ;
        RECT 296.025 37.295 296.810 37.305 ;
        RECT 295.920 37.280 296.815 37.295 ;
        RECT 295.920 37.265 296.835 37.280 ;
        RECT 295.920 37.255 296.855 37.265 ;
        RECT 295.920 37.245 296.880 37.255 ;
        RECT 295.920 37.215 296.950 37.245 ;
        RECT 295.920 37.185 296.970 37.215 ;
        RECT 295.920 37.155 296.990 37.185 ;
        RECT 295.920 37.130 297.020 37.155 ;
        RECT 295.920 37.095 297.055 37.130 ;
        RECT 295.920 37.090 297.085 37.095 ;
        RECT 295.920 36.695 296.150 37.090 ;
        RECT 296.695 37.085 297.085 37.090 ;
        RECT 296.720 37.075 297.085 37.085 ;
        RECT 296.735 37.070 297.085 37.075 ;
        RECT 296.750 37.065 297.085 37.070 ;
        RECT 297.450 37.065 297.710 37.515 ;
        RECT 298.065 37.370 298.455 37.545 ;
        RECT 298.940 37.540 299.270 38.340 ;
        RECT 299.440 37.550 299.975 38.170 ;
        RECT 298.065 37.200 299.490 37.370 ;
        RECT 296.750 37.060 297.710 37.065 ;
        RECT 296.760 37.050 297.710 37.060 ;
        RECT 296.770 37.045 297.710 37.050 ;
        RECT 296.780 37.035 297.710 37.045 ;
        RECT 296.785 37.025 297.710 37.035 ;
        RECT 296.790 37.020 297.710 37.025 ;
        RECT 296.800 37.005 297.710 37.020 ;
        RECT 296.805 36.990 297.710 37.005 ;
        RECT 296.815 36.965 297.710 36.990 ;
        RECT 296.320 36.495 296.650 36.920 ;
        RECT 295.580 35.960 295.840 36.440 ;
        RECT 296.010 35.790 296.260 36.330 ;
        RECT 296.430 36.010 296.650 36.495 ;
        RECT 296.820 36.895 297.710 36.965 ;
        RECT 296.820 36.170 296.990 36.895 ;
        RECT 297.160 36.340 297.710 36.725 ;
        RECT 297.940 36.470 298.295 37.030 ;
        RECT 298.465 36.300 298.635 37.200 ;
        RECT 298.805 36.470 299.070 37.030 ;
        RECT 299.320 36.700 299.490 37.200 ;
        RECT 299.660 36.530 299.975 37.550 ;
        RECT 300.295 37.710 300.580 38.170 ;
        RECT 300.750 37.880 301.020 38.340 ;
        RECT 300.295 37.490 301.250 37.710 ;
        RECT 300.180 36.760 300.870 37.320 ;
        RECT 301.040 36.590 301.250 37.490 ;
        RECT 296.820 36.000 297.710 36.170 ;
        RECT 298.045 35.790 298.285 36.300 ;
        RECT 298.465 35.970 298.745 36.300 ;
        RECT 298.975 35.790 299.190 36.300 ;
        RECT 299.360 35.960 299.975 36.530 ;
        RECT 300.295 36.420 301.250 36.590 ;
        RECT 301.420 37.320 301.820 38.170 ;
        RECT 302.010 37.710 302.290 38.170 ;
        RECT 302.810 37.880 303.135 38.340 ;
        RECT 302.010 37.490 303.135 37.710 ;
        RECT 301.420 36.760 302.515 37.320 ;
        RECT 302.685 37.030 303.135 37.490 ;
        RECT 303.305 37.200 303.690 38.170 ;
        RECT 300.295 35.960 300.580 36.420 ;
        RECT 300.750 35.790 301.020 36.250 ;
        RECT 301.420 35.960 301.820 36.760 ;
        RECT 302.685 36.700 303.240 37.030 ;
        RECT 302.685 36.590 303.135 36.700 ;
        RECT 302.010 36.420 303.135 36.590 ;
        RECT 303.410 36.530 303.690 37.200 ;
        RECT 303.860 37.175 304.150 38.340 ;
        RECT 305.245 37.915 305.580 38.340 ;
        RECT 305.750 37.735 305.935 38.140 ;
        RECT 305.270 37.560 305.935 37.735 ;
        RECT 306.140 37.560 306.470 38.340 ;
        RECT 302.010 35.960 302.290 36.420 ;
        RECT 302.810 35.790 303.135 36.250 ;
        RECT 303.305 35.960 303.690 36.530 ;
        RECT 305.270 36.530 305.610 37.560 ;
        RECT 306.640 37.370 306.910 38.140 ;
        RECT 305.780 37.200 306.910 37.370 ;
        RECT 307.080 37.250 309.670 38.340 ;
        RECT 305.780 36.700 306.030 37.200 ;
        RECT 303.860 35.790 304.150 36.515 ;
        RECT 305.270 36.360 305.955 36.530 ;
        RECT 306.210 36.450 306.570 37.030 ;
        RECT 305.245 35.790 305.580 36.190 ;
        RECT 305.750 35.960 305.955 36.360 ;
        RECT 306.740 36.290 306.910 37.200 ;
        RECT 306.165 35.790 306.440 36.270 ;
        RECT 306.650 35.960 306.910 36.290 ;
        RECT 307.080 36.560 308.290 37.080 ;
        RECT 308.460 36.730 309.670 37.250 ;
        RECT 309.840 37.250 311.050 38.340 ;
        RECT 309.840 36.710 310.360 37.250 ;
        RECT 307.080 35.790 309.670 36.560 ;
        RECT 310.530 36.540 311.050 37.080 ;
        RECT 309.840 35.790 311.050 36.540 ;
        RECT 162.095 35.620 311.135 35.790 ;
        RECT 162.180 34.870 163.390 35.620 ;
        RECT 162.180 34.330 162.700 34.870 ;
        RECT 163.560 34.850 167.070 35.620 ;
        RECT 167.245 35.070 167.500 35.360 ;
        RECT 167.670 35.240 168.000 35.620 ;
        RECT 167.245 34.900 167.995 35.070 ;
        RECT 162.870 34.160 163.390 34.700 ;
        RECT 163.560 34.330 165.210 34.850 ;
        RECT 165.380 34.160 167.070 34.680 ;
        RECT 162.180 33.070 163.390 34.160 ;
        RECT 163.560 33.070 167.070 34.160 ;
        RECT 167.245 34.080 167.595 34.730 ;
        RECT 167.765 33.910 167.995 34.900 ;
        RECT 167.245 33.740 167.995 33.910 ;
        RECT 167.245 33.240 167.500 33.740 ;
        RECT 167.670 33.070 168.000 33.570 ;
        RECT 168.170 33.240 168.340 35.360 ;
        RECT 168.700 35.260 169.030 35.620 ;
        RECT 169.200 35.230 169.695 35.400 ;
        RECT 169.900 35.230 170.755 35.400 ;
        RECT 168.570 34.040 169.030 35.090 ;
        RECT 168.510 33.255 168.835 34.040 ;
        RECT 169.200 33.870 169.370 35.230 ;
        RECT 169.540 34.320 169.890 34.940 ;
        RECT 170.060 34.720 170.415 34.940 ;
        RECT 170.060 34.130 170.230 34.720 ;
        RECT 170.585 34.520 170.755 35.230 ;
        RECT 171.630 35.160 171.960 35.620 ;
        RECT 172.170 35.260 172.520 35.430 ;
        RECT 170.960 34.690 171.750 34.940 ;
        RECT 172.170 34.870 172.430 35.260 ;
        RECT 172.740 35.170 173.690 35.450 ;
        RECT 173.860 35.180 174.050 35.620 ;
        RECT 174.220 35.240 175.290 35.410 ;
        RECT 171.920 34.520 172.090 34.700 ;
        RECT 169.200 33.700 169.595 33.870 ;
        RECT 169.765 33.740 170.230 34.130 ;
        RECT 170.400 34.350 172.090 34.520 ;
        RECT 169.425 33.570 169.595 33.700 ;
        RECT 170.400 33.570 170.570 34.350 ;
        RECT 172.260 34.180 172.430 34.870 ;
        RECT 170.930 34.010 172.430 34.180 ;
        RECT 172.620 34.210 172.830 35.000 ;
        RECT 173.000 34.380 173.350 35.000 ;
        RECT 173.520 34.390 173.690 35.170 ;
        RECT 174.220 35.010 174.390 35.240 ;
        RECT 173.860 34.840 174.390 35.010 ;
        RECT 173.860 34.560 174.080 34.840 ;
        RECT 174.560 34.670 174.800 35.070 ;
        RECT 173.520 34.220 173.925 34.390 ;
        RECT 174.260 34.300 174.800 34.670 ;
        RECT 174.970 34.885 175.290 35.240 ;
        RECT 175.535 35.160 175.840 35.620 ;
        RECT 176.010 34.910 176.265 35.440 ;
        RECT 174.970 34.710 175.295 34.885 ;
        RECT 174.970 34.410 175.885 34.710 ;
        RECT 175.145 34.380 175.885 34.410 ;
        RECT 172.620 34.050 173.295 34.210 ;
        RECT 173.755 34.130 173.925 34.220 ;
        RECT 172.620 34.040 173.585 34.050 ;
        RECT 172.260 33.870 172.430 34.010 ;
        RECT 169.005 33.070 169.255 33.530 ;
        RECT 169.425 33.240 169.675 33.570 ;
        RECT 169.890 33.240 170.570 33.570 ;
        RECT 170.740 33.670 171.815 33.840 ;
        RECT 172.260 33.700 172.820 33.870 ;
        RECT 173.125 33.750 173.585 34.040 ;
        RECT 173.755 33.960 174.975 34.130 ;
        RECT 170.740 33.330 170.910 33.670 ;
        RECT 171.145 33.070 171.475 33.500 ;
        RECT 171.645 33.330 171.815 33.670 ;
        RECT 172.110 33.070 172.480 33.530 ;
        RECT 172.650 33.240 172.820 33.700 ;
        RECT 173.755 33.580 173.925 33.960 ;
        RECT 175.145 33.790 175.315 34.380 ;
        RECT 176.055 34.260 176.265 34.910 ;
        RECT 173.055 33.240 173.925 33.580 ;
        RECT 174.515 33.620 175.315 33.790 ;
        RECT 174.095 33.070 174.345 33.530 ;
        RECT 174.515 33.330 174.685 33.620 ;
        RECT 174.865 33.070 175.195 33.450 ;
        RECT 175.535 33.070 175.840 34.210 ;
        RECT 176.010 33.380 176.265 34.260 ;
        RECT 176.445 34.880 176.700 35.450 ;
        RECT 176.870 35.220 177.200 35.620 ;
        RECT 177.625 35.085 178.155 35.450 ;
        RECT 178.345 35.280 178.620 35.450 ;
        RECT 178.340 35.110 178.620 35.280 ;
        RECT 177.625 35.050 177.800 35.085 ;
        RECT 176.870 34.880 177.800 35.050 ;
        RECT 176.445 34.210 176.615 34.880 ;
        RECT 176.870 34.710 177.040 34.880 ;
        RECT 176.785 34.380 177.040 34.710 ;
        RECT 177.265 34.380 177.460 34.710 ;
        RECT 176.445 33.240 176.780 34.210 ;
        RECT 176.950 33.070 177.120 34.210 ;
        RECT 177.290 33.410 177.460 34.380 ;
        RECT 177.630 33.750 177.800 34.880 ;
        RECT 177.970 34.090 178.140 34.890 ;
        RECT 178.345 34.290 178.620 35.110 ;
        RECT 178.790 34.090 178.980 35.450 ;
        RECT 179.160 35.085 179.670 35.620 ;
        RECT 179.890 34.810 180.135 35.415 ;
        RECT 180.580 35.075 185.925 35.620 ;
        RECT 179.180 34.640 180.410 34.810 ;
        RECT 177.970 33.920 178.980 34.090 ;
        RECT 179.150 34.075 179.900 34.265 ;
        RECT 177.630 33.580 178.755 33.750 ;
        RECT 179.150 33.410 179.320 34.075 ;
        RECT 180.070 33.830 180.410 34.640 ;
        RECT 182.165 34.245 182.505 35.075 ;
        RECT 186.100 34.850 187.770 35.620 ;
        RECT 187.940 34.895 188.230 35.620 ;
        RECT 188.400 34.870 189.610 35.620 ;
        RECT 177.290 33.240 179.320 33.410 ;
        RECT 179.490 33.070 179.660 33.830 ;
        RECT 179.895 33.420 180.410 33.830 ;
        RECT 183.985 33.505 184.335 34.755 ;
        RECT 186.100 34.330 186.850 34.850 ;
        RECT 187.020 34.160 187.770 34.680 ;
        RECT 188.400 34.330 188.920 34.870 ;
        RECT 190.055 34.810 190.300 35.415 ;
        RECT 190.520 35.085 191.030 35.620 ;
        RECT 180.580 33.070 185.925 33.505 ;
        RECT 186.100 33.070 187.770 34.160 ;
        RECT 187.940 33.070 188.230 34.235 ;
        RECT 189.090 34.160 189.610 34.700 ;
        RECT 188.400 33.070 189.610 34.160 ;
        RECT 189.780 34.640 191.010 34.810 ;
        RECT 189.780 33.830 190.120 34.640 ;
        RECT 190.290 34.075 191.040 34.265 ;
        RECT 189.780 33.420 190.295 33.830 ;
        RECT 190.530 33.070 190.700 33.830 ;
        RECT 190.870 33.410 191.040 34.075 ;
        RECT 191.210 34.090 191.400 35.450 ;
        RECT 191.570 34.600 191.845 35.450 ;
        RECT 192.035 35.085 192.565 35.450 ;
        RECT 192.990 35.220 193.320 35.620 ;
        RECT 192.390 35.050 192.565 35.085 ;
        RECT 191.570 34.430 191.850 34.600 ;
        RECT 191.570 34.290 191.845 34.430 ;
        RECT 192.050 34.090 192.220 34.890 ;
        RECT 191.210 33.920 192.220 34.090 ;
        RECT 192.390 34.880 193.320 35.050 ;
        RECT 193.490 34.880 193.745 35.450 ;
        RECT 192.390 33.750 192.560 34.880 ;
        RECT 193.150 34.710 193.320 34.880 ;
        RECT 191.435 33.580 192.560 33.750 ;
        RECT 192.730 34.380 192.925 34.710 ;
        RECT 193.150 34.380 193.405 34.710 ;
        RECT 192.730 33.410 192.900 34.380 ;
        RECT 193.575 34.210 193.745 34.880 ;
        RECT 190.870 33.240 192.900 33.410 ;
        RECT 193.070 33.070 193.240 34.210 ;
        RECT 193.410 33.240 193.745 34.210 ;
        RECT 193.920 34.945 194.180 35.450 ;
        RECT 194.360 35.240 194.690 35.620 ;
        RECT 194.870 35.070 195.040 35.450 ;
        RECT 193.920 34.145 194.090 34.945 ;
        RECT 194.375 34.900 195.040 35.070 ;
        RECT 194.375 34.645 194.545 34.900 ;
        RECT 195.300 34.850 198.810 35.620 ;
        RECT 198.980 34.870 200.190 35.620 ;
        RECT 200.475 34.990 200.760 35.450 ;
        RECT 200.930 35.160 201.200 35.620 ;
        RECT 194.260 34.315 194.545 34.645 ;
        RECT 194.780 34.350 195.110 34.720 ;
        RECT 195.300 34.330 196.950 34.850 ;
        RECT 194.375 34.170 194.545 34.315 ;
        RECT 193.920 33.240 194.190 34.145 ;
        RECT 194.375 34.000 195.040 34.170 ;
        RECT 197.120 34.160 198.810 34.680 ;
        RECT 198.980 34.330 199.500 34.870 ;
        RECT 200.475 34.820 201.430 34.990 ;
        RECT 199.670 34.160 200.190 34.700 ;
        RECT 194.360 33.070 194.690 33.830 ;
        RECT 194.870 33.240 195.040 34.000 ;
        RECT 195.300 33.070 198.810 34.160 ;
        RECT 198.980 33.070 200.190 34.160 ;
        RECT 200.360 34.090 201.050 34.650 ;
        RECT 201.220 33.920 201.430 34.820 ;
        RECT 200.475 33.700 201.430 33.920 ;
        RECT 201.600 34.650 202.000 35.450 ;
        RECT 202.190 34.990 202.470 35.450 ;
        RECT 202.990 35.160 203.315 35.620 ;
        RECT 202.190 34.820 203.315 34.990 ;
        RECT 203.485 34.880 203.870 35.450 ;
        RECT 202.865 34.710 203.315 34.820 ;
        RECT 201.600 34.090 202.695 34.650 ;
        RECT 202.865 34.380 203.420 34.710 ;
        RECT 200.475 33.240 200.760 33.700 ;
        RECT 200.930 33.070 201.200 33.530 ;
        RECT 201.600 33.240 202.000 34.090 ;
        RECT 202.865 33.920 203.315 34.380 ;
        RECT 203.590 34.210 203.870 34.880 ;
        RECT 202.190 33.700 203.315 33.920 ;
        RECT 202.190 33.240 202.470 33.700 ;
        RECT 202.990 33.070 203.315 33.530 ;
        RECT 203.485 33.240 203.870 34.210 ;
        RECT 204.045 34.880 204.300 35.450 ;
        RECT 204.470 35.220 204.800 35.620 ;
        RECT 205.225 35.085 205.755 35.450 ;
        RECT 205.225 35.050 205.400 35.085 ;
        RECT 204.470 34.880 205.400 35.050 ;
        RECT 204.045 34.210 204.215 34.880 ;
        RECT 204.470 34.710 204.640 34.880 ;
        RECT 204.385 34.380 204.640 34.710 ;
        RECT 204.865 34.380 205.060 34.710 ;
        RECT 204.045 33.240 204.380 34.210 ;
        RECT 204.550 33.070 204.720 34.210 ;
        RECT 204.890 33.410 205.060 34.380 ;
        RECT 205.230 33.750 205.400 34.880 ;
        RECT 205.570 34.090 205.740 34.890 ;
        RECT 205.945 34.600 206.220 35.450 ;
        RECT 205.940 34.430 206.220 34.600 ;
        RECT 205.945 34.290 206.220 34.430 ;
        RECT 206.390 34.090 206.580 35.450 ;
        RECT 206.760 35.085 207.270 35.620 ;
        RECT 207.490 34.810 207.735 35.415 ;
        RECT 208.180 34.945 208.440 35.450 ;
        RECT 208.620 35.240 208.950 35.620 ;
        RECT 209.130 35.070 209.300 35.450 ;
        RECT 206.780 34.640 208.010 34.810 ;
        RECT 205.570 33.920 206.580 34.090 ;
        RECT 206.750 34.075 207.500 34.265 ;
        RECT 205.230 33.580 206.355 33.750 ;
        RECT 206.750 33.410 206.920 34.075 ;
        RECT 207.670 33.830 208.010 34.640 ;
        RECT 204.890 33.240 206.920 33.410 ;
        RECT 207.090 33.070 207.260 33.830 ;
        RECT 207.495 33.420 208.010 33.830 ;
        RECT 208.180 34.145 208.350 34.945 ;
        RECT 208.635 34.900 209.300 35.070 ;
        RECT 208.635 34.645 208.805 34.900 ;
        RECT 209.565 34.880 209.820 35.450 ;
        RECT 209.990 35.220 210.320 35.620 ;
        RECT 210.745 35.085 211.275 35.450 ;
        RECT 211.465 35.280 211.740 35.450 ;
        RECT 211.460 35.110 211.740 35.280 ;
        RECT 210.745 35.050 210.920 35.085 ;
        RECT 209.990 34.880 210.920 35.050 ;
        RECT 208.520 34.315 208.805 34.645 ;
        RECT 209.040 34.350 209.370 34.720 ;
        RECT 208.635 34.170 208.805 34.315 ;
        RECT 209.565 34.210 209.735 34.880 ;
        RECT 209.990 34.710 210.160 34.880 ;
        RECT 209.905 34.380 210.160 34.710 ;
        RECT 210.385 34.380 210.580 34.710 ;
        RECT 208.180 33.240 208.450 34.145 ;
        RECT 208.635 34.000 209.300 34.170 ;
        RECT 208.620 33.070 208.950 33.830 ;
        RECT 209.130 33.240 209.300 34.000 ;
        RECT 209.565 33.240 209.900 34.210 ;
        RECT 210.070 33.070 210.240 34.210 ;
        RECT 210.410 33.410 210.580 34.380 ;
        RECT 210.750 33.750 210.920 34.880 ;
        RECT 211.090 34.090 211.260 34.890 ;
        RECT 211.465 34.290 211.740 35.110 ;
        RECT 211.910 34.090 212.100 35.450 ;
        RECT 212.280 35.085 212.790 35.620 ;
        RECT 213.010 34.810 213.255 35.415 ;
        RECT 213.700 34.895 213.990 35.620 ;
        RECT 214.620 34.880 215.005 35.450 ;
        RECT 215.175 35.160 215.500 35.620 ;
        RECT 216.020 34.990 216.300 35.450 ;
        RECT 212.300 34.640 213.530 34.810 ;
        RECT 211.090 33.920 212.100 34.090 ;
        RECT 212.270 34.075 213.020 34.265 ;
        RECT 210.750 33.580 211.875 33.750 ;
        RECT 212.270 33.410 212.440 34.075 ;
        RECT 213.190 33.830 213.530 34.640 ;
        RECT 210.410 33.240 212.440 33.410 ;
        RECT 212.610 33.070 212.780 33.830 ;
        RECT 213.015 33.420 213.530 33.830 ;
        RECT 213.700 33.070 213.990 34.235 ;
        RECT 214.620 34.210 214.900 34.880 ;
        RECT 215.175 34.820 216.300 34.990 ;
        RECT 215.175 34.710 215.625 34.820 ;
        RECT 215.070 34.380 215.625 34.710 ;
        RECT 216.490 34.650 216.890 35.450 ;
        RECT 217.290 35.160 217.560 35.620 ;
        RECT 217.730 34.990 218.015 35.450 ;
        RECT 214.620 33.240 215.005 34.210 ;
        RECT 215.175 33.920 215.625 34.380 ;
        RECT 215.795 34.090 216.890 34.650 ;
        RECT 215.175 33.700 216.300 33.920 ;
        RECT 215.175 33.070 215.500 33.530 ;
        RECT 216.020 33.240 216.300 33.700 ;
        RECT 216.490 33.240 216.890 34.090 ;
        RECT 217.060 34.820 218.015 34.990 ;
        RECT 218.305 34.880 218.560 35.450 ;
        RECT 218.730 35.220 219.060 35.620 ;
        RECT 219.485 35.085 220.015 35.450 ;
        RECT 219.485 35.050 219.660 35.085 ;
        RECT 218.730 34.880 219.660 35.050 ;
        RECT 217.060 33.920 217.270 34.820 ;
        RECT 217.440 34.090 218.130 34.650 ;
        RECT 218.305 34.210 218.475 34.880 ;
        RECT 218.730 34.710 218.900 34.880 ;
        RECT 218.645 34.380 218.900 34.710 ;
        RECT 219.125 34.380 219.320 34.710 ;
        RECT 217.060 33.700 218.015 33.920 ;
        RECT 217.290 33.070 217.560 33.530 ;
        RECT 217.730 33.240 218.015 33.700 ;
        RECT 218.305 33.240 218.640 34.210 ;
        RECT 218.810 33.070 218.980 34.210 ;
        RECT 219.150 33.410 219.320 34.380 ;
        RECT 219.490 33.750 219.660 34.880 ;
        RECT 219.830 34.090 220.000 34.890 ;
        RECT 220.205 34.600 220.480 35.450 ;
        RECT 220.200 34.430 220.480 34.600 ;
        RECT 220.205 34.290 220.480 34.430 ;
        RECT 220.650 34.090 220.840 35.450 ;
        RECT 221.020 35.085 221.530 35.620 ;
        RECT 221.750 34.810 221.995 35.415 ;
        RECT 222.445 34.880 222.700 35.450 ;
        RECT 222.870 35.220 223.200 35.620 ;
        RECT 223.625 35.085 224.155 35.450 ;
        RECT 223.625 35.050 223.800 35.085 ;
        RECT 222.870 34.880 223.800 35.050 ;
        RECT 221.040 34.640 222.270 34.810 ;
        RECT 219.830 33.920 220.840 34.090 ;
        RECT 221.010 34.075 221.760 34.265 ;
        RECT 219.490 33.580 220.615 33.750 ;
        RECT 221.010 33.410 221.180 34.075 ;
        RECT 221.930 33.830 222.270 34.640 ;
        RECT 219.150 33.240 221.180 33.410 ;
        RECT 221.350 33.070 221.520 33.830 ;
        RECT 221.755 33.420 222.270 33.830 ;
        RECT 222.445 34.210 222.615 34.880 ;
        RECT 222.870 34.710 223.040 34.880 ;
        RECT 222.785 34.380 223.040 34.710 ;
        RECT 223.265 34.380 223.460 34.710 ;
        RECT 222.445 33.240 222.780 34.210 ;
        RECT 222.950 33.070 223.120 34.210 ;
        RECT 223.290 33.410 223.460 34.380 ;
        RECT 223.630 33.750 223.800 34.880 ;
        RECT 223.970 34.090 224.140 34.890 ;
        RECT 224.345 34.600 224.620 35.450 ;
        RECT 224.340 34.430 224.620 34.600 ;
        RECT 224.345 34.290 224.620 34.430 ;
        RECT 224.790 34.090 224.980 35.450 ;
        RECT 225.160 35.085 225.670 35.620 ;
        RECT 225.890 34.810 226.135 35.415 ;
        RECT 226.695 34.990 226.980 35.450 ;
        RECT 227.150 35.160 227.420 35.620 ;
        RECT 226.695 34.820 227.650 34.990 ;
        RECT 225.180 34.640 226.410 34.810 ;
        RECT 223.970 33.920 224.980 34.090 ;
        RECT 225.150 34.075 225.900 34.265 ;
        RECT 223.630 33.580 224.755 33.750 ;
        RECT 225.150 33.410 225.320 34.075 ;
        RECT 226.070 33.830 226.410 34.640 ;
        RECT 226.580 34.090 227.270 34.650 ;
        RECT 227.440 33.920 227.650 34.820 ;
        RECT 223.290 33.240 225.320 33.410 ;
        RECT 225.490 33.070 225.660 33.830 ;
        RECT 225.895 33.420 226.410 33.830 ;
        RECT 226.695 33.700 227.650 33.920 ;
        RECT 227.820 34.650 228.220 35.450 ;
        RECT 228.410 34.990 228.690 35.450 ;
        RECT 229.210 35.160 229.535 35.620 ;
        RECT 228.410 34.820 229.535 34.990 ;
        RECT 229.705 34.880 230.090 35.450 ;
        RECT 230.265 35.070 230.520 35.360 ;
        RECT 230.690 35.240 231.020 35.620 ;
        RECT 230.265 34.900 231.015 35.070 ;
        RECT 229.085 34.710 229.535 34.820 ;
        RECT 227.820 34.090 228.915 34.650 ;
        RECT 229.085 34.380 229.640 34.710 ;
        RECT 226.695 33.240 226.980 33.700 ;
        RECT 227.150 33.070 227.420 33.530 ;
        RECT 227.820 33.240 228.220 34.090 ;
        RECT 229.085 33.920 229.535 34.380 ;
        RECT 229.810 34.210 230.090 34.880 ;
        RECT 228.410 33.700 229.535 33.920 ;
        RECT 228.410 33.240 228.690 33.700 ;
        RECT 229.210 33.070 229.535 33.530 ;
        RECT 229.705 33.240 230.090 34.210 ;
        RECT 230.265 34.080 230.615 34.730 ;
        RECT 230.785 33.910 231.015 34.900 ;
        RECT 230.265 33.740 231.015 33.910 ;
        RECT 230.265 33.240 230.520 33.740 ;
        RECT 230.690 33.070 231.020 33.570 ;
        RECT 231.190 33.240 231.360 35.360 ;
        RECT 231.720 35.260 232.050 35.620 ;
        RECT 232.220 35.230 232.715 35.400 ;
        RECT 232.920 35.230 233.775 35.400 ;
        RECT 231.590 34.040 232.050 35.090 ;
        RECT 231.530 33.255 231.855 34.040 ;
        RECT 232.220 33.870 232.390 35.230 ;
        RECT 232.560 34.320 232.910 34.940 ;
        RECT 233.080 34.720 233.435 34.940 ;
        RECT 233.080 34.130 233.250 34.720 ;
        RECT 233.605 34.520 233.775 35.230 ;
        RECT 234.650 35.160 234.980 35.620 ;
        RECT 235.190 35.260 235.540 35.430 ;
        RECT 233.980 34.690 234.770 34.940 ;
        RECT 235.190 34.870 235.450 35.260 ;
        RECT 235.760 35.170 236.710 35.450 ;
        RECT 236.880 35.180 237.070 35.620 ;
        RECT 237.240 35.240 238.310 35.410 ;
        RECT 234.940 34.520 235.110 34.700 ;
        RECT 232.220 33.700 232.615 33.870 ;
        RECT 232.785 33.740 233.250 34.130 ;
        RECT 233.420 34.350 235.110 34.520 ;
        RECT 232.445 33.570 232.615 33.700 ;
        RECT 233.420 33.570 233.590 34.350 ;
        RECT 235.280 34.180 235.450 34.870 ;
        RECT 233.950 34.010 235.450 34.180 ;
        RECT 235.640 34.210 235.850 35.000 ;
        RECT 236.020 34.380 236.370 35.000 ;
        RECT 236.540 34.390 236.710 35.170 ;
        RECT 237.240 35.010 237.410 35.240 ;
        RECT 236.880 34.840 237.410 35.010 ;
        RECT 236.880 34.560 237.100 34.840 ;
        RECT 237.580 34.670 237.820 35.070 ;
        RECT 236.540 34.220 236.945 34.390 ;
        RECT 237.280 34.300 237.820 34.670 ;
        RECT 237.990 34.885 238.310 35.240 ;
        RECT 238.555 35.160 238.860 35.620 ;
        RECT 239.030 34.910 239.285 35.440 ;
        RECT 237.990 34.710 238.315 34.885 ;
        RECT 237.990 34.410 238.905 34.710 ;
        RECT 238.165 34.380 238.905 34.410 ;
        RECT 235.640 34.050 236.315 34.210 ;
        RECT 236.775 34.130 236.945 34.220 ;
        RECT 235.640 34.040 236.605 34.050 ;
        RECT 235.280 33.870 235.450 34.010 ;
        RECT 232.025 33.070 232.275 33.530 ;
        RECT 232.445 33.240 232.695 33.570 ;
        RECT 232.910 33.240 233.590 33.570 ;
        RECT 233.760 33.670 234.835 33.840 ;
        RECT 235.280 33.700 235.840 33.870 ;
        RECT 236.145 33.750 236.605 34.040 ;
        RECT 236.775 33.960 237.995 34.130 ;
        RECT 233.760 33.330 233.930 33.670 ;
        RECT 234.165 33.070 234.495 33.500 ;
        RECT 234.665 33.330 234.835 33.670 ;
        RECT 235.130 33.070 235.500 33.530 ;
        RECT 235.670 33.240 235.840 33.700 ;
        RECT 236.775 33.580 236.945 33.960 ;
        RECT 238.165 33.790 238.335 34.380 ;
        RECT 239.075 34.260 239.285 34.910 ;
        RECT 239.460 34.895 239.750 35.620 ;
        RECT 240.930 35.070 241.100 35.450 ;
        RECT 241.280 35.240 241.610 35.620 ;
        RECT 240.930 34.900 241.595 35.070 ;
        RECT 241.790 34.945 242.050 35.450 ;
        RECT 240.860 34.350 241.190 34.720 ;
        RECT 241.425 34.645 241.595 34.900 ;
        RECT 236.075 33.240 236.945 33.580 ;
        RECT 237.535 33.620 238.335 33.790 ;
        RECT 237.115 33.070 237.365 33.530 ;
        RECT 237.535 33.330 237.705 33.620 ;
        RECT 237.885 33.070 238.215 33.450 ;
        RECT 238.555 33.070 238.860 34.210 ;
        RECT 239.030 33.380 239.285 34.260 ;
        RECT 241.425 34.315 241.710 34.645 ;
        RECT 239.460 33.070 239.750 34.235 ;
        RECT 241.425 34.170 241.595 34.315 ;
        RECT 240.930 34.000 241.595 34.170 ;
        RECT 241.880 34.145 242.050 34.945 ;
        RECT 242.225 35.070 242.480 35.360 ;
        RECT 242.650 35.240 242.980 35.620 ;
        RECT 242.225 34.900 242.975 35.070 ;
        RECT 240.930 33.240 241.100 34.000 ;
        RECT 241.280 33.070 241.610 33.830 ;
        RECT 241.780 33.240 242.050 34.145 ;
        RECT 242.225 34.080 242.575 34.730 ;
        RECT 242.745 33.910 242.975 34.900 ;
        RECT 242.225 33.740 242.975 33.910 ;
        RECT 242.225 33.240 242.480 33.740 ;
        RECT 242.650 33.070 242.980 33.570 ;
        RECT 243.150 33.240 243.320 35.360 ;
        RECT 243.680 35.260 244.010 35.620 ;
        RECT 244.180 35.230 244.675 35.400 ;
        RECT 244.880 35.230 245.735 35.400 ;
        RECT 243.550 34.040 244.010 35.090 ;
        RECT 243.490 33.255 243.815 34.040 ;
        RECT 244.180 33.870 244.350 35.230 ;
        RECT 244.520 34.320 244.870 34.940 ;
        RECT 245.040 34.720 245.395 34.940 ;
        RECT 245.040 34.130 245.210 34.720 ;
        RECT 245.565 34.520 245.735 35.230 ;
        RECT 246.610 35.160 246.940 35.620 ;
        RECT 247.150 35.260 247.500 35.430 ;
        RECT 245.940 34.690 246.730 34.940 ;
        RECT 247.150 34.870 247.410 35.260 ;
        RECT 247.720 35.170 248.670 35.450 ;
        RECT 248.840 35.180 249.030 35.620 ;
        RECT 249.200 35.240 250.270 35.410 ;
        RECT 246.900 34.520 247.070 34.700 ;
        RECT 244.180 33.700 244.575 33.870 ;
        RECT 244.745 33.740 245.210 34.130 ;
        RECT 245.380 34.350 247.070 34.520 ;
        RECT 244.405 33.570 244.575 33.700 ;
        RECT 245.380 33.570 245.550 34.350 ;
        RECT 247.240 34.180 247.410 34.870 ;
        RECT 245.910 34.010 247.410 34.180 ;
        RECT 247.600 34.210 247.810 35.000 ;
        RECT 247.980 34.380 248.330 35.000 ;
        RECT 248.500 34.390 248.670 35.170 ;
        RECT 249.200 35.010 249.370 35.240 ;
        RECT 248.840 34.840 249.370 35.010 ;
        RECT 248.840 34.560 249.060 34.840 ;
        RECT 249.540 34.670 249.780 35.070 ;
        RECT 248.500 34.220 248.905 34.390 ;
        RECT 249.240 34.300 249.780 34.670 ;
        RECT 249.950 34.885 250.270 35.240 ;
        RECT 250.515 35.160 250.820 35.620 ;
        RECT 250.990 34.910 251.245 35.440 ;
        RECT 249.950 34.710 250.275 34.885 ;
        RECT 249.950 34.410 250.865 34.710 ;
        RECT 250.125 34.380 250.865 34.410 ;
        RECT 247.600 34.050 248.275 34.210 ;
        RECT 248.735 34.130 248.905 34.220 ;
        RECT 247.600 34.040 248.565 34.050 ;
        RECT 247.240 33.870 247.410 34.010 ;
        RECT 243.985 33.070 244.235 33.530 ;
        RECT 244.405 33.240 244.655 33.570 ;
        RECT 244.870 33.240 245.550 33.570 ;
        RECT 245.720 33.670 246.795 33.840 ;
        RECT 247.240 33.700 247.800 33.870 ;
        RECT 248.105 33.750 248.565 34.040 ;
        RECT 248.735 33.960 249.955 34.130 ;
        RECT 245.720 33.330 245.890 33.670 ;
        RECT 246.125 33.070 246.455 33.500 ;
        RECT 246.625 33.330 246.795 33.670 ;
        RECT 247.090 33.070 247.460 33.530 ;
        RECT 247.630 33.240 247.800 33.700 ;
        RECT 248.735 33.580 248.905 33.960 ;
        RECT 250.125 33.790 250.295 34.380 ;
        RECT 251.035 34.260 251.245 34.910 ;
        RECT 248.035 33.240 248.905 33.580 ;
        RECT 249.495 33.620 250.295 33.790 ;
        RECT 249.075 33.070 249.325 33.530 ;
        RECT 249.495 33.330 249.665 33.620 ;
        RECT 249.845 33.070 250.175 33.450 ;
        RECT 250.515 33.070 250.820 34.210 ;
        RECT 250.990 33.380 251.245 34.260 ;
        RECT 251.420 34.880 251.805 35.450 ;
        RECT 251.975 35.160 252.300 35.620 ;
        RECT 252.820 34.990 253.100 35.450 ;
        RECT 251.420 34.210 251.700 34.880 ;
        RECT 251.975 34.820 253.100 34.990 ;
        RECT 251.975 34.710 252.425 34.820 ;
        RECT 251.870 34.380 252.425 34.710 ;
        RECT 253.290 34.650 253.690 35.450 ;
        RECT 254.090 35.160 254.360 35.620 ;
        RECT 254.530 34.990 254.815 35.450 ;
        RECT 255.100 35.075 260.445 35.620 ;
        RECT 251.420 33.240 251.805 34.210 ;
        RECT 251.975 33.920 252.425 34.380 ;
        RECT 252.595 34.090 253.690 34.650 ;
        RECT 251.975 33.700 253.100 33.920 ;
        RECT 251.975 33.070 252.300 33.530 ;
        RECT 252.820 33.240 253.100 33.700 ;
        RECT 253.290 33.240 253.690 34.090 ;
        RECT 253.860 34.820 254.815 34.990 ;
        RECT 253.860 33.920 254.070 34.820 ;
        RECT 254.240 34.090 254.930 34.650 ;
        RECT 256.685 34.245 257.025 35.075 ;
        RECT 260.620 34.850 264.130 35.620 ;
        RECT 265.220 34.895 265.510 35.620 ;
        RECT 265.680 34.850 268.270 35.620 ;
        RECT 268.450 35.110 269.680 35.450 ;
        RECT 269.850 35.130 270.105 35.620 ;
        RECT 268.450 34.880 268.780 35.110 ;
        RECT 253.860 33.700 254.815 33.920 ;
        RECT 254.090 33.070 254.360 33.530 ;
        RECT 254.530 33.240 254.815 33.700 ;
        RECT 258.505 33.505 258.855 34.755 ;
        RECT 260.620 34.330 262.270 34.850 ;
        RECT 262.440 34.160 264.130 34.680 ;
        RECT 265.680 34.330 266.890 34.850 ;
        RECT 255.100 33.070 260.445 33.505 ;
        RECT 260.620 33.070 264.130 34.160 ;
        RECT 265.220 33.070 265.510 34.235 ;
        RECT 267.060 34.160 268.270 34.680 ;
        RECT 268.440 34.380 268.750 34.710 ;
        RECT 268.955 34.380 269.330 34.940 ;
        RECT 269.500 34.210 269.680 35.110 ;
        RECT 269.865 34.380 270.085 34.960 ;
        RECT 270.285 34.910 270.540 35.440 ;
        RECT 270.710 35.160 271.015 35.620 ;
        RECT 271.260 35.240 272.330 35.410 ;
        RECT 270.285 34.260 270.495 34.910 ;
        RECT 271.260 34.885 271.580 35.240 ;
        RECT 271.255 34.710 271.580 34.885 ;
        RECT 270.665 34.410 271.580 34.710 ;
        RECT 271.750 34.670 271.990 35.070 ;
        RECT 272.160 35.010 272.330 35.240 ;
        RECT 272.500 35.180 272.690 35.620 ;
        RECT 272.860 35.170 273.810 35.450 ;
        RECT 274.030 35.260 274.380 35.430 ;
        RECT 272.160 34.840 272.690 35.010 ;
        RECT 270.665 34.380 271.405 34.410 ;
        RECT 265.680 33.070 268.270 34.160 ;
        RECT 268.450 34.040 269.680 34.210 ;
        RECT 268.450 33.240 268.780 34.040 ;
        RECT 268.950 33.070 269.180 33.870 ;
        RECT 269.350 33.240 269.680 34.040 ;
        RECT 269.850 33.070 270.105 34.210 ;
        RECT 270.285 33.380 270.540 34.260 ;
        RECT 270.710 33.070 271.015 34.210 ;
        RECT 271.235 33.790 271.405 34.380 ;
        RECT 271.750 34.300 272.290 34.670 ;
        RECT 272.470 34.560 272.690 34.840 ;
        RECT 272.860 34.390 273.030 35.170 ;
        RECT 272.625 34.220 273.030 34.390 ;
        RECT 273.200 34.380 273.550 35.000 ;
        RECT 272.625 34.130 272.795 34.220 ;
        RECT 273.720 34.210 273.930 35.000 ;
        RECT 271.575 33.960 272.795 34.130 ;
        RECT 273.255 34.050 273.930 34.210 ;
        RECT 271.235 33.620 272.035 33.790 ;
        RECT 271.355 33.070 271.685 33.450 ;
        RECT 271.865 33.330 272.035 33.620 ;
        RECT 272.625 33.580 272.795 33.960 ;
        RECT 272.965 34.040 273.930 34.050 ;
        RECT 274.120 34.870 274.380 35.260 ;
        RECT 274.590 35.160 274.920 35.620 ;
        RECT 275.795 35.230 276.650 35.400 ;
        RECT 276.855 35.230 277.350 35.400 ;
        RECT 277.520 35.260 277.850 35.620 ;
        RECT 274.120 34.180 274.290 34.870 ;
        RECT 274.460 34.520 274.630 34.700 ;
        RECT 274.800 34.690 275.590 34.940 ;
        RECT 275.795 34.520 275.965 35.230 ;
        RECT 276.135 34.720 276.490 34.940 ;
        RECT 274.460 34.350 276.150 34.520 ;
        RECT 272.965 33.750 273.425 34.040 ;
        RECT 274.120 34.010 275.620 34.180 ;
        RECT 274.120 33.870 274.290 34.010 ;
        RECT 273.730 33.700 274.290 33.870 ;
        RECT 272.205 33.070 272.455 33.530 ;
        RECT 272.625 33.240 273.495 33.580 ;
        RECT 273.730 33.240 273.900 33.700 ;
        RECT 274.735 33.670 275.810 33.840 ;
        RECT 274.070 33.070 274.440 33.530 ;
        RECT 274.735 33.330 274.905 33.670 ;
        RECT 275.075 33.070 275.405 33.500 ;
        RECT 275.640 33.330 275.810 33.670 ;
        RECT 275.980 33.570 276.150 34.350 ;
        RECT 276.320 34.130 276.490 34.720 ;
        RECT 276.660 34.320 277.010 34.940 ;
        RECT 276.320 33.740 276.785 34.130 ;
        RECT 277.180 33.870 277.350 35.230 ;
        RECT 277.520 34.040 277.980 35.090 ;
        RECT 276.955 33.700 277.350 33.870 ;
        RECT 276.955 33.570 277.125 33.700 ;
        RECT 275.980 33.240 276.660 33.570 ;
        RECT 276.875 33.240 277.125 33.570 ;
        RECT 277.295 33.070 277.545 33.530 ;
        RECT 277.715 33.255 278.040 34.040 ;
        RECT 278.210 33.240 278.380 35.360 ;
        RECT 278.550 35.240 278.880 35.620 ;
        RECT 279.050 35.070 279.305 35.360 ;
        RECT 278.555 34.900 279.305 35.070 ;
        RECT 279.595 34.990 279.880 35.450 ;
        RECT 280.050 35.160 280.320 35.620 ;
        RECT 278.555 33.910 278.785 34.900 ;
        RECT 279.595 34.820 280.550 34.990 ;
        RECT 278.955 34.080 279.305 34.730 ;
        RECT 279.480 34.090 280.170 34.650 ;
        RECT 280.340 33.920 280.550 34.820 ;
        RECT 278.555 33.740 279.305 33.910 ;
        RECT 278.550 33.070 278.880 33.570 ;
        RECT 279.050 33.240 279.305 33.740 ;
        RECT 279.595 33.700 280.550 33.920 ;
        RECT 280.720 34.650 281.120 35.450 ;
        RECT 281.310 34.990 281.590 35.450 ;
        RECT 282.110 35.160 282.435 35.620 ;
        RECT 281.310 34.820 282.435 34.990 ;
        RECT 282.605 34.880 282.990 35.450 ;
        RECT 281.985 34.710 282.435 34.820 ;
        RECT 280.720 34.090 281.815 34.650 ;
        RECT 281.985 34.380 282.540 34.710 ;
        RECT 279.595 33.240 279.880 33.700 ;
        RECT 280.050 33.070 280.320 33.530 ;
        RECT 280.720 33.240 281.120 34.090 ;
        RECT 281.985 33.920 282.435 34.380 ;
        RECT 282.710 34.210 282.990 34.880 ;
        RECT 283.160 34.850 284.830 35.620 ;
        RECT 285.060 35.140 285.340 35.620 ;
        RECT 285.510 34.970 285.770 35.360 ;
        RECT 285.945 35.140 286.200 35.620 ;
        RECT 286.370 34.970 286.665 35.360 ;
        RECT 286.845 35.140 287.120 35.620 ;
        RECT 287.290 35.120 287.590 35.450 ;
        RECT 283.160 34.330 283.910 34.850 ;
        RECT 285.015 34.800 286.665 34.970 ;
        RECT 281.310 33.700 282.435 33.920 ;
        RECT 281.310 33.240 281.590 33.700 ;
        RECT 282.110 33.070 282.435 33.530 ;
        RECT 282.605 33.240 282.990 34.210 ;
        RECT 284.080 34.160 284.830 34.680 ;
        RECT 283.160 33.070 284.830 34.160 ;
        RECT 285.015 34.290 285.420 34.800 ;
        RECT 285.590 34.460 286.730 34.630 ;
        RECT 285.015 34.120 285.770 34.290 ;
        RECT 285.055 33.070 285.340 33.940 ;
        RECT 285.510 33.870 285.770 34.120 ;
        RECT 286.560 34.210 286.730 34.460 ;
        RECT 286.900 34.380 287.250 34.950 ;
        RECT 287.420 34.210 287.590 35.120 ;
        RECT 286.560 34.040 287.590 34.210 ;
        RECT 285.510 33.700 286.630 33.870 ;
        RECT 285.510 33.240 285.770 33.700 ;
        RECT 285.945 33.070 286.200 33.530 ;
        RECT 286.370 33.240 286.630 33.700 ;
        RECT 286.800 33.070 287.110 33.870 ;
        RECT 287.280 33.240 287.590 34.040 ;
        RECT 287.760 34.945 288.035 35.290 ;
        RECT 288.225 35.220 288.600 35.620 ;
        RECT 288.770 35.050 288.940 35.400 ;
        RECT 289.110 35.220 289.440 35.620 ;
        RECT 289.610 35.050 289.870 35.450 ;
        RECT 287.760 34.210 287.930 34.945 ;
        RECT 288.205 34.880 289.870 35.050 ;
        RECT 288.205 34.710 288.375 34.880 ;
        RECT 290.050 34.800 290.380 35.220 ;
        RECT 290.550 34.800 290.810 35.620 ;
        RECT 290.980 34.895 291.270 35.620 ;
        RECT 291.500 34.800 291.710 35.620 ;
        RECT 291.880 34.820 292.210 35.450 ;
        RECT 290.050 34.710 290.300 34.800 ;
        RECT 288.100 34.380 288.375 34.710 ;
        RECT 288.545 34.380 289.370 34.710 ;
        RECT 289.585 34.380 290.300 34.710 ;
        RECT 290.470 34.380 290.805 34.630 ;
        RECT 288.205 34.210 288.375 34.380 ;
        RECT 287.760 33.240 288.035 34.210 ;
        RECT 288.205 34.040 288.865 34.210 ;
        RECT 289.125 34.090 289.370 34.380 ;
        RECT 288.695 33.920 288.865 34.040 ;
        RECT 289.540 33.920 289.870 34.210 ;
        RECT 288.245 33.070 288.525 33.870 ;
        RECT 288.695 33.750 289.870 33.920 ;
        RECT 290.130 33.820 290.300 34.380 ;
        RECT 288.695 33.250 290.310 33.580 ;
        RECT 290.550 33.070 290.810 34.210 ;
        RECT 290.980 33.070 291.270 34.235 ;
        RECT 291.880 34.220 292.130 34.820 ;
        RECT 292.380 34.800 292.610 35.620 ;
        RECT 293.280 34.880 293.665 35.450 ;
        RECT 293.835 35.160 294.160 35.620 ;
        RECT 294.680 34.990 294.960 35.450 ;
        RECT 292.300 34.380 292.630 34.630 ;
        RECT 291.500 33.070 291.710 34.210 ;
        RECT 291.880 33.240 292.210 34.220 ;
        RECT 293.280 34.210 293.560 34.880 ;
        RECT 293.835 34.820 294.960 34.990 ;
        RECT 293.835 34.710 294.285 34.820 ;
        RECT 293.730 34.380 294.285 34.710 ;
        RECT 295.150 34.650 295.550 35.450 ;
        RECT 295.950 35.160 296.220 35.620 ;
        RECT 296.390 34.990 296.675 35.450 ;
        RECT 297.885 35.220 298.220 35.620 ;
        RECT 298.390 35.050 298.595 35.450 ;
        RECT 298.805 35.140 299.080 35.620 ;
        RECT 299.290 35.120 299.550 35.450 ;
        RECT 292.380 33.070 292.610 34.210 ;
        RECT 293.280 33.240 293.665 34.210 ;
        RECT 293.835 33.920 294.285 34.380 ;
        RECT 294.455 34.090 295.550 34.650 ;
        RECT 293.835 33.700 294.960 33.920 ;
        RECT 293.835 33.070 294.160 33.530 ;
        RECT 294.680 33.240 294.960 33.700 ;
        RECT 295.150 33.240 295.550 34.090 ;
        RECT 295.720 34.820 296.675 34.990 ;
        RECT 297.910 34.880 298.595 35.050 ;
        RECT 295.720 33.920 295.930 34.820 ;
        RECT 296.100 34.090 296.790 34.650 ;
        RECT 295.720 33.700 296.675 33.920 ;
        RECT 295.950 33.070 296.220 33.530 ;
        RECT 296.390 33.240 296.675 33.700 ;
        RECT 297.910 33.850 298.250 34.880 ;
        RECT 298.420 34.210 298.670 34.710 ;
        RECT 298.850 34.380 299.210 34.960 ;
        RECT 299.380 34.210 299.550 35.120 ;
        RECT 298.420 34.040 299.550 34.210 ;
        RECT 297.910 33.675 298.575 33.850 ;
        RECT 297.885 33.070 298.220 33.495 ;
        RECT 298.390 33.270 298.575 33.675 ;
        RECT 298.780 33.070 299.110 33.850 ;
        RECT 299.280 33.270 299.550 34.040 ;
        RECT 299.725 34.910 299.980 35.440 ;
        RECT 300.150 35.160 300.455 35.620 ;
        RECT 300.700 35.240 301.770 35.410 ;
        RECT 299.725 34.260 299.935 34.910 ;
        RECT 300.700 34.885 301.020 35.240 ;
        RECT 300.695 34.710 301.020 34.885 ;
        RECT 300.105 34.410 301.020 34.710 ;
        RECT 301.190 34.670 301.430 35.070 ;
        RECT 301.600 35.010 301.770 35.240 ;
        RECT 301.940 35.180 302.130 35.620 ;
        RECT 302.300 35.170 303.250 35.450 ;
        RECT 303.470 35.260 303.820 35.430 ;
        RECT 301.600 34.840 302.130 35.010 ;
        RECT 300.105 34.380 300.845 34.410 ;
        RECT 299.725 33.380 299.980 34.260 ;
        RECT 300.150 33.070 300.455 34.210 ;
        RECT 300.675 33.790 300.845 34.380 ;
        RECT 301.190 34.300 301.730 34.670 ;
        RECT 301.910 34.560 302.130 34.840 ;
        RECT 302.300 34.390 302.470 35.170 ;
        RECT 302.065 34.220 302.470 34.390 ;
        RECT 302.640 34.380 302.990 35.000 ;
        RECT 302.065 34.130 302.235 34.220 ;
        RECT 303.160 34.210 303.370 35.000 ;
        RECT 301.015 33.960 302.235 34.130 ;
        RECT 302.695 34.050 303.370 34.210 ;
        RECT 300.675 33.620 301.475 33.790 ;
        RECT 300.795 33.070 301.125 33.450 ;
        RECT 301.305 33.330 301.475 33.620 ;
        RECT 302.065 33.580 302.235 33.960 ;
        RECT 302.405 34.040 303.370 34.050 ;
        RECT 303.560 34.870 303.820 35.260 ;
        RECT 304.030 35.160 304.360 35.620 ;
        RECT 305.235 35.230 306.090 35.400 ;
        RECT 306.295 35.230 306.790 35.400 ;
        RECT 306.960 35.260 307.290 35.620 ;
        RECT 303.560 34.180 303.730 34.870 ;
        RECT 303.900 34.520 304.070 34.700 ;
        RECT 304.240 34.690 305.030 34.940 ;
        RECT 305.235 34.520 305.405 35.230 ;
        RECT 305.575 34.720 305.930 34.940 ;
        RECT 303.900 34.350 305.590 34.520 ;
        RECT 302.405 33.750 302.865 34.040 ;
        RECT 303.560 34.010 305.060 34.180 ;
        RECT 303.560 33.870 303.730 34.010 ;
        RECT 303.170 33.700 303.730 33.870 ;
        RECT 301.645 33.070 301.895 33.530 ;
        RECT 302.065 33.240 302.935 33.580 ;
        RECT 303.170 33.240 303.340 33.700 ;
        RECT 304.175 33.670 305.250 33.840 ;
        RECT 303.510 33.070 303.880 33.530 ;
        RECT 304.175 33.330 304.345 33.670 ;
        RECT 304.515 33.070 304.845 33.500 ;
        RECT 305.080 33.330 305.250 33.670 ;
        RECT 305.420 33.570 305.590 34.350 ;
        RECT 305.760 34.130 305.930 34.720 ;
        RECT 306.100 34.320 306.450 34.940 ;
        RECT 305.760 33.740 306.225 34.130 ;
        RECT 306.620 33.870 306.790 35.230 ;
        RECT 306.960 34.040 307.420 35.090 ;
        RECT 306.395 33.700 306.790 33.870 ;
        RECT 306.395 33.570 306.565 33.700 ;
        RECT 305.420 33.240 306.100 33.570 ;
        RECT 306.315 33.240 306.565 33.570 ;
        RECT 306.735 33.070 306.985 33.530 ;
        RECT 307.155 33.255 307.480 34.040 ;
        RECT 307.650 33.240 307.820 35.360 ;
        RECT 307.990 35.240 308.320 35.620 ;
        RECT 308.490 35.070 308.745 35.360 ;
        RECT 307.995 34.900 308.745 35.070 ;
        RECT 307.995 33.910 308.225 34.900 ;
        RECT 309.840 34.870 311.050 35.620 ;
        RECT 308.395 34.080 308.745 34.730 ;
        RECT 309.840 34.160 310.360 34.700 ;
        RECT 310.530 34.330 311.050 34.870 ;
        RECT 307.995 33.740 308.745 33.910 ;
        RECT 307.990 33.070 308.320 33.570 ;
        RECT 308.490 33.240 308.745 33.740 ;
        RECT 309.840 33.070 311.050 34.160 ;
        RECT 162.095 32.900 311.135 33.070 ;
        RECT 162.180 31.810 163.390 32.900 ;
        RECT 163.560 32.465 168.905 32.900 ;
        RECT 162.180 31.100 162.700 31.640 ;
        RECT 162.870 31.270 163.390 31.810 ;
        RECT 162.180 30.350 163.390 31.100 ;
        RECT 165.145 30.895 165.485 31.725 ;
        RECT 166.965 31.215 167.315 32.465 ;
        RECT 169.080 31.825 169.350 32.730 ;
        RECT 169.520 32.140 169.850 32.900 ;
        RECT 170.030 31.970 170.200 32.730 ;
        RECT 169.080 31.025 169.250 31.825 ;
        RECT 169.535 31.800 170.200 31.970 ;
        RECT 170.920 31.825 171.190 32.730 ;
        RECT 171.360 32.140 171.690 32.900 ;
        RECT 171.870 31.970 172.040 32.730 ;
        RECT 169.535 31.655 169.705 31.800 ;
        RECT 169.420 31.325 169.705 31.655 ;
        RECT 169.535 31.070 169.705 31.325 ;
        RECT 169.940 31.250 170.270 31.620 ;
        RECT 163.560 30.350 168.905 30.895 ;
        RECT 169.080 30.520 169.340 31.025 ;
        RECT 169.535 30.900 170.200 31.070 ;
        RECT 169.520 30.350 169.850 30.730 ;
        RECT 170.030 30.520 170.200 30.900 ;
        RECT 170.920 31.025 171.090 31.825 ;
        RECT 171.375 31.800 172.040 31.970 ;
        RECT 172.300 31.810 174.890 32.900 ;
        RECT 171.375 31.655 171.545 31.800 ;
        RECT 171.260 31.325 171.545 31.655 ;
        RECT 171.375 31.070 171.545 31.325 ;
        RECT 171.780 31.250 172.110 31.620 ;
        RECT 172.300 31.120 173.510 31.640 ;
        RECT 173.680 31.290 174.890 31.810 ;
        RECT 175.060 31.735 175.350 32.900 ;
        RECT 175.525 31.760 175.860 32.730 ;
        RECT 176.030 31.760 176.200 32.900 ;
        RECT 176.370 32.560 178.400 32.730 ;
        RECT 170.920 30.520 171.180 31.025 ;
        RECT 171.375 30.900 172.040 31.070 ;
        RECT 171.360 30.350 171.690 30.730 ;
        RECT 171.870 30.520 172.040 30.900 ;
        RECT 172.300 30.350 174.890 31.120 ;
        RECT 175.525 31.090 175.695 31.760 ;
        RECT 176.370 31.590 176.540 32.560 ;
        RECT 175.865 31.260 176.120 31.590 ;
        RECT 176.345 31.260 176.540 31.590 ;
        RECT 176.710 32.220 177.835 32.390 ;
        RECT 175.950 31.090 176.120 31.260 ;
        RECT 176.710 31.090 176.880 32.220 ;
        RECT 175.060 30.350 175.350 31.075 ;
        RECT 175.525 30.520 175.780 31.090 ;
        RECT 175.950 30.920 176.880 31.090 ;
        RECT 177.050 31.880 178.060 32.050 ;
        RECT 177.050 31.080 177.220 31.880 ;
        RECT 176.705 30.885 176.880 30.920 ;
        RECT 175.950 30.350 176.280 30.750 ;
        RECT 176.705 30.520 177.235 30.885 ;
        RECT 177.425 30.860 177.700 31.680 ;
        RECT 177.420 30.690 177.700 30.860 ;
        RECT 177.425 30.520 177.700 30.690 ;
        RECT 177.870 30.520 178.060 31.880 ;
        RECT 178.230 31.895 178.400 32.560 ;
        RECT 178.570 32.140 178.740 32.900 ;
        RECT 178.975 32.140 179.490 32.550 ;
        RECT 178.230 31.705 178.980 31.895 ;
        RECT 179.150 31.330 179.490 32.140 ;
        RECT 178.260 31.160 179.490 31.330 ;
        RECT 179.665 31.710 179.920 32.590 ;
        RECT 180.090 31.760 180.395 32.900 ;
        RECT 180.735 32.520 181.065 32.900 ;
        RECT 181.245 32.350 181.415 32.640 ;
        RECT 181.585 32.440 181.835 32.900 ;
        RECT 180.615 32.180 181.415 32.350 ;
        RECT 182.005 32.390 182.875 32.730 ;
        RECT 178.240 30.350 178.750 30.885 ;
        RECT 178.970 30.555 179.215 31.160 ;
        RECT 179.665 31.060 179.875 31.710 ;
        RECT 180.615 31.590 180.785 32.180 ;
        RECT 182.005 32.010 182.175 32.390 ;
        RECT 183.110 32.270 183.280 32.730 ;
        RECT 183.450 32.440 183.820 32.900 ;
        RECT 184.115 32.300 184.285 32.640 ;
        RECT 184.455 32.470 184.785 32.900 ;
        RECT 185.020 32.300 185.190 32.640 ;
        RECT 180.955 31.840 182.175 32.010 ;
        RECT 182.345 31.930 182.805 32.220 ;
        RECT 183.110 32.100 183.670 32.270 ;
        RECT 184.115 32.130 185.190 32.300 ;
        RECT 185.360 32.400 186.040 32.730 ;
        RECT 186.255 32.400 186.505 32.730 ;
        RECT 186.675 32.440 186.925 32.900 ;
        RECT 183.500 31.960 183.670 32.100 ;
        RECT 182.345 31.920 183.310 31.930 ;
        RECT 182.005 31.750 182.175 31.840 ;
        RECT 182.635 31.760 183.310 31.920 ;
        RECT 180.045 31.560 180.785 31.590 ;
        RECT 180.045 31.260 180.960 31.560 ;
        RECT 180.635 31.085 180.960 31.260 ;
        RECT 179.665 30.530 179.920 31.060 ;
        RECT 180.090 30.350 180.395 30.810 ;
        RECT 180.640 30.730 180.960 31.085 ;
        RECT 181.130 31.300 181.670 31.670 ;
        RECT 182.005 31.580 182.410 31.750 ;
        RECT 181.130 30.900 181.370 31.300 ;
        RECT 181.850 31.130 182.070 31.410 ;
        RECT 181.540 30.960 182.070 31.130 ;
        RECT 181.540 30.730 181.710 30.960 ;
        RECT 182.240 30.800 182.410 31.580 ;
        RECT 182.580 30.970 182.930 31.590 ;
        RECT 183.100 30.970 183.310 31.760 ;
        RECT 183.500 31.790 185.000 31.960 ;
        RECT 183.500 31.100 183.670 31.790 ;
        RECT 185.360 31.620 185.530 32.400 ;
        RECT 186.335 32.270 186.505 32.400 ;
        RECT 183.840 31.450 185.530 31.620 ;
        RECT 185.700 31.840 186.165 32.230 ;
        RECT 186.335 32.100 186.730 32.270 ;
        RECT 183.840 31.270 184.010 31.450 ;
        RECT 180.640 30.560 181.710 30.730 ;
        RECT 181.880 30.350 182.070 30.790 ;
        RECT 182.240 30.520 183.190 30.800 ;
        RECT 183.500 30.710 183.760 31.100 ;
        RECT 184.180 31.030 184.970 31.280 ;
        RECT 183.410 30.540 183.760 30.710 ;
        RECT 183.970 30.350 184.300 30.810 ;
        RECT 185.175 30.740 185.345 31.450 ;
        RECT 185.700 31.250 185.870 31.840 ;
        RECT 185.515 31.030 185.870 31.250 ;
        RECT 186.040 31.030 186.390 31.650 ;
        RECT 186.560 30.740 186.730 32.100 ;
        RECT 187.095 31.930 187.420 32.715 ;
        RECT 186.900 30.880 187.360 31.930 ;
        RECT 185.175 30.570 186.030 30.740 ;
        RECT 186.235 30.570 186.730 30.740 ;
        RECT 186.900 30.350 187.230 30.710 ;
        RECT 187.590 30.610 187.760 32.730 ;
        RECT 187.930 32.400 188.260 32.900 ;
        RECT 188.430 32.230 188.685 32.730 ;
        RECT 187.935 32.060 188.685 32.230 ;
        RECT 188.865 32.230 189.120 32.730 ;
        RECT 189.290 32.400 189.620 32.900 ;
        RECT 188.865 32.060 189.615 32.230 ;
        RECT 187.935 31.070 188.165 32.060 ;
        RECT 188.335 31.240 188.685 31.890 ;
        RECT 188.865 31.240 189.215 31.890 ;
        RECT 189.385 31.070 189.615 32.060 ;
        RECT 187.935 30.900 188.685 31.070 ;
        RECT 187.930 30.350 188.260 30.730 ;
        RECT 188.430 30.610 188.685 30.900 ;
        RECT 188.865 30.900 189.615 31.070 ;
        RECT 188.865 30.610 189.120 30.900 ;
        RECT 189.290 30.350 189.620 30.730 ;
        RECT 189.790 30.610 189.960 32.730 ;
        RECT 190.130 31.930 190.455 32.715 ;
        RECT 190.625 32.440 190.875 32.900 ;
        RECT 191.045 32.400 191.295 32.730 ;
        RECT 191.510 32.400 192.190 32.730 ;
        RECT 191.045 32.270 191.215 32.400 ;
        RECT 190.820 32.100 191.215 32.270 ;
        RECT 190.190 30.880 190.650 31.930 ;
        RECT 190.820 30.740 190.990 32.100 ;
        RECT 191.385 31.840 191.850 32.230 ;
        RECT 191.160 31.030 191.510 31.650 ;
        RECT 191.680 31.250 191.850 31.840 ;
        RECT 192.020 31.620 192.190 32.400 ;
        RECT 192.360 32.300 192.530 32.640 ;
        RECT 192.765 32.470 193.095 32.900 ;
        RECT 193.265 32.300 193.435 32.640 ;
        RECT 193.730 32.440 194.100 32.900 ;
        RECT 192.360 32.130 193.435 32.300 ;
        RECT 194.270 32.270 194.440 32.730 ;
        RECT 194.675 32.390 195.545 32.730 ;
        RECT 195.715 32.440 195.965 32.900 ;
        RECT 193.880 32.100 194.440 32.270 ;
        RECT 193.880 31.960 194.050 32.100 ;
        RECT 192.550 31.790 194.050 31.960 ;
        RECT 194.745 31.930 195.205 32.220 ;
        RECT 192.020 31.450 193.710 31.620 ;
        RECT 191.680 31.030 192.035 31.250 ;
        RECT 192.205 30.740 192.375 31.450 ;
        RECT 192.580 31.030 193.370 31.280 ;
        RECT 193.540 31.270 193.710 31.450 ;
        RECT 193.880 31.100 194.050 31.790 ;
        RECT 190.320 30.350 190.650 30.710 ;
        RECT 190.820 30.570 191.315 30.740 ;
        RECT 191.520 30.570 192.375 30.740 ;
        RECT 193.250 30.350 193.580 30.810 ;
        RECT 193.790 30.710 194.050 31.100 ;
        RECT 194.240 31.920 195.205 31.930 ;
        RECT 195.375 32.010 195.545 32.390 ;
        RECT 196.135 32.350 196.305 32.640 ;
        RECT 196.485 32.520 196.815 32.900 ;
        RECT 196.135 32.180 196.935 32.350 ;
        RECT 194.240 31.760 194.915 31.920 ;
        RECT 195.375 31.840 196.595 32.010 ;
        RECT 194.240 30.970 194.450 31.760 ;
        RECT 195.375 31.750 195.545 31.840 ;
        RECT 194.620 30.970 194.970 31.590 ;
        RECT 195.140 31.580 195.545 31.750 ;
        RECT 195.140 30.800 195.310 31.580 ;
        RECT 195.480 31.130 195.700 31.410 ;
        RECT 195.880 31.300 196.420 31.670 ;
        RECT 196.765 31.590 196.935 32.180 ;
        RECT 197.155 31.760 197.460 32.900 ;
        RECT 197.630 31.710 197.885 32.590 ;
        RECT 198.060 31.810 200.650 32.900 ;
        RECT 196.765 31.560 197.505 31.590 ;
        RECT 195.480 30.960 196.010 31.130 ;
        RECT 193.790 30.540 194.140 30.710 ;
        RECT 194.360 30.520 195.310 30.800 ;
        RECT 195.480 30.350 195.670 30.790 ;
        RECT 195.840 30.730 196.010 30.960 ;
        RECT 196.180 30.900 196.420 31.300 ;
        RECT 196.590 31.260 197.505 31.560 ;
        RECT 196.590 31.085 196.915 31.260 ;
        RECT 196.590 30.730 196.910 31.085 ;
        RECT 197.675 31.060 197.885 31.710 ;
        RECT 195.840 30.560 196.910 30.730 ;
        RECT 197.155 30.350 197.460 30.810 ;
        RECT 197.630 30.530 197.885 31.060 ;
        RECT 198.060 31.120 199.270 31.640 ;
        RECT 199.440 31.290 200.650 31.810 ;
        RECT 200.820 31.735 201.110 32.900 ;
        RECT 201.280 31.810 202.490 32.900 ;
        RECT 202.715 32.030 203.000 32.900 ;
        RECT 203.170 32.270 203.430 32.730 ;
        RECT 203.605 32.440 203.860 32.900 ;
        RECT 204.030 32.270 204.290 32.730 ;
        RECT 203.170 32.100 204.290 32.270 ;
        RECT 204.460 32.100 204.770 32.900 ;
        RECT 203.170 31.850 203.430 32.100 ;
        RECT 204.940 31.930 205.250 32.730 ;
        RECT 198.060 30.350 200.650 31.120 ;
        RECT 201.280 31.100 201.800 31.640 ;
        RECT 201.970 31.270 202.490 31.810 ;
        RECT 202.675 31.680 203.430 31.850 ;
        RECT 204.220 31.760 205.250 31.930 ;
        RECT 202.675 31.170 203.080 31.680 ;
        RECT 204.220 31.510 204.390 31.760 ;
        RECT 203.250 31.340 204.390 31.510 ;
        RECT 200.820 30.350 201.110 31.075 ;
        RECT 201.280 30.350 202.490 31.100 ;
        RECT 202.675 31.000 204.325 31.170 ;
        RECT 204.560 31.020 204.910 31.590 ;
        RECT 202.720 30.350 203.000 30.830 ;
        RECT 203.170 30.610 203.430 31.000 ;
        RECT 203.605 30.350 203.860 30.830 ;
        RECT 204.030 30.610 204.325 31.000 ;
        RECT 205.080 30.850 205.250 31.760 ;
        RECT 204.505 30.350 204.780 30.830 ;
        RECT 204.950 30.520 205.250 30.850 ;
        RECT 205.425 31.710 205.680 32.590 ;
        RECT 205.850 31.760 206.155 32.900 ;
        RECT 206.495 32.520 206.825 32.900 ;
        RECT 207.005 32.350 207.175 32.640 ;
        RECT 207.345 32.440 207.595 32.900 ;
        RECT 206.375 32.180 207.175 32.350 ;
        RECT 207.765 32.390 208.635 32.730 ;
        RECT 205.425 31.060 205.635 31.710 ;
        RECT 206.375 31.590 206.545 32.180 ;
        RECT 207.765 32.010 207.935 32.390 ;
        RECT 208.870 32.270 209.040 32.730 ;
        RECT 209.210 32.440 209.580 32.900 ;
        RECT 209.875 32.300 210.045 32.640 ;
        RECT 210.215 32.470 210.545 32.900 ;
        RECT 210.780 32.300 210.950 32.640 ;
        RECT 206.715 31.840 207.935 32.010 ;
        RECT 208.105 31.930 208.565 32.220 ;
        RECT 208.870 32.100 209.430 32.270 ;
        RECT 209.875 32.130 210.950 32.300 ;
        RECT 211.120 32.400 211.800 32.730 ;
        RECT 212.015 32.400 212.265 32.730 ;
        RECT 212.435 32.440 212.685 32.900 ;
        RECT 209.260 31.960 209.430 32.100 ;
        RECT 208.105 31.920 209.070 31.930 ;
        RECT 207.765 31.750 207.935 31.840 ;
        RECT 208.395 31.760 209.070 31.920 ;
        RECT 205.805 31.560 206.545 31.590 ;
        RECT 205.805 31.260 206.720 31.560 ;
        RECT 206.395 31.085 206.720 31.260 ;
        RECT 205.425 30.530 205.680 31.060 ;
        RECT 205.850 30.350 206.155 30.810 ;
        RECT 206.400 30.730 206.720 31.085 ;
        RECT 206.890 31.300 207.430 31.670 ;
        RECT 207.765 31.580 208.170 31.750 ;
        RECT 206.890 30.900 207.130 31.300 ;
        RECT 207.610 31.130 207.830 31.410 ;
        RECT 207.300 30.960 207.830 31.130 ;
        RECT 207.300 30.730 207.470 30.960 ;
        RECT 208.000 30.800 208.170 31.580 ;
        RECT 208.340 30.970 208.690 31.590 ;
        RECT 208.860 30.970 209.070 31.760 ;
        RECT 209.260 31.790 210.760 31.960 ;
        RECT 209.260 31.100 209.430 31.790 ;
        RECT 211.120 31.620 211.290 32.400 ;
        RECT 212.095 32.270 212.265 32.400 ;
        RECT 209.600 31.450 211.290 31.620 ;
        RECT 211.460 31.840 211.925 32.230 ;
        RECT 212.095 32.100 212.490 32.270 ;
        RECT 209.600 31.270 209.770 31.450 ;
        RECT 206.400 30.560 207.470 30.730 ;
        RECT 207.640 30.350 207.830 30.790 ;
        RECT 208.000 30.520 208.950 30.800 ;
        RECT 209.260 30.710 209.520 31.100 ;
        RECT 209.940 31.030 210.730 31.280 ;
        RECT 209.170 30.540 209.520 30.710 ;
        RECT 209.730 30.350 210.060 30.810 ;
        RECT 210.935 30.740 211.105 31.450 ;
        RECT 211.460 31.250 211.630 31.840 ;
        RECT 211.275 31.030 211.630 31.250 ;
        RECT 211.800 31.030 212.150 31.650 ;
        RECT 212.320 30.740 212.490 32.100 ;
        RECT 212.855 31.930 213.180 32.715 ;
        RECT 212.660 30.880 213.120 31.930 ;
        RECT 210.935 30.570 211.790 30.740 ;
        RECT 211.995 30.570 212.490 30.740 ;
        RECT 212.660 30.350 212.990 30.710 ;
        RECT 213.350 30.610 213.520 32.730 ;
        RECT 213.690 32.400 214.020 32.900 ;
        RECT 214.190 32.230 214.445 32.730 ;
        RECT 213.695 32.060 214.445 32.230 ;
        RECT 213.695 31.070 213.925 32.060 ;
        RECT 214.095 31.240 214.445 31.890 ;
        RECT 214.620 31.825 214.890 32.730 ;
        RECT 215.060 32.140 215.390 32.900 ;
        RECT 215.570 31.970 215.740 32.730 ;
        RECT 213.695 30.900 214.445 31.070 ;
        RECT 213.690 30.350 214.020 30.730 ;
        RECT 214.190 30.610 214.445 30.900 ;
        RECT 214.620 31.025 214.790 31.825 ;
        RECT 215.075 31.800 215.740 31.970 ;
        RECT 216.000 31.825 216.270 32.730 ;
        RECT 216.440 32.140 216.770 32.900 ;
        RECT 216.950 31.970 217.120 32.730 ;
        RECT 217.385 32.230 217.640 32.730 ;
        RECT 217.810 32.400 218.140 32.900 ;
        RECT 217.385 32.060 218.135 32.230 ;
        RECT 215.075 31.655 215.245 31.800 ;
        RECT 214.960 31.325 215.245 31.655 ;
        RECT 215.075 31.070 215.245 31.325 ;
        RECT 215.480 31.250 215.810 31.620 ;
        RECT 214.620 30.520 214.880 31.025 ;
        RECT 215.075 30.900 215.740 31.070 ;
        RECT 215.060 30.350 215.390 30.730 ;
        RECT 215.570 30.520 215.740 30.900 ;
        RECT 216.000 31.025 216.170 31.825 ;
        RECT 216.455 31.800 217.120 31.970 ;
        RECT 216.455 31.655 216.625 31.800 ;
        RECT 216.340 31.325 216.625 31.655 ;
        RECT 216.455 31.070 216.625 31.325 ;
        RECT 216.860 31.250 217.190 31.620 ;
        RECT 217.385 31.240 217.735 31.890 ;
        RECT 217.905 31.070 218.135 32.060 ;
        RECT 216.000 30.520 216.260 31.025 ;
        RECT 216.455 30.900 217.120 31.070 ;
        RECT 216.440 30.350 216.770 30.730 ;
        RECT 216.950 30.520 217.120 30.900 ;
        RECT 217.385 30.900 218.135 31.070 ;
        RECT 217.385 30.610 217.640 30.900 ;
        RECT 217.810 30.350 218.140 30.730 ;
        RECT 218.310 30.610 218.480 32.730 ;
        RECT 218.650 31.930 218.975 32.715 ;
        RECT 219.145 32.440 219.395 32.900 ;
        RECT 219.565 32.400 219.815 32.730 ;
        RECT 220.030 32.400 220.710 32.730 ;
        RECT 219.565 32.270 219.735 32.400 ;
        RECT 219.340 32.100 219.735 32.270 ;
        RECT 218.710 30.880 219.170 31.930 ;
        RECT 219.340 30.740 219.510 32.100 ;
        RECT 219.905 31.840 220.370 32.230 ;
        RECT 219.680 31.030 220.030 31.650 ;
        RECT 220.200 31.250 220.370 31.840 ;
        RECT 220.540 31.620 220.710 32.400 ;
        RECT 220.880 32.300 221.050 32.640 ;
        RECT 221.285 32.470 221.615 32.900 ;
        RECT 221.785 32.300 221.955 32.640 ;
        RECT 222.250 32.440 222.620 32.900 ;
        RECT 220.880 32.130 221.955 32.300 ;
        RECT 222.790 32.270 222.960 32.730 ;
        RECT 223.195 32.390 224.065 32.730 ;
        RECT 224.235 32.440 224.485 32.900 ;
        RECT 222.400 32.100 222.960 32.270 ;
        RECT 222.400 31.960 222.570 32.100 ;
        RECT 221.070 31.790 222.570 31.960 ;
        RECT 223.265 31.930 223.725 32.220 ;
        RECT 220.540 31.450 222.230 31.620 ;
        RECT 220.200 31.030 220.555 31.250 ;
        RECT 220.725 30.740 220.895 31.450 ;
        RECT 221.100 31.030 221.890 31.280 ;
        RECT 222.060 31.270 222.230 31.450 ;
        RECT 222.400 31.100 222.570 31.790 ;
        RECT 218.840 30.350 219.170 30.710 ;
        RECT 219.340 30.570 219.835 30.740 ;
        RECT 220.040 30.570 220.895 30.740 ;
        RECT 221.770 30.350 222.100 30.810 ;
        RECT 222.310 30.710 222.570 31.100 ;
        RECT 222.760 31.920 223.725 31.930 ;
        RECT 223.895 32.010 224.065 32.390 ;
        RECT 224.655 32.350 224.825 32.640 ;
        RECT 225.005 32.520 225.335 32.900 ;
        RECT 224.655 32.180 225.455 32.350 ;
        RECT 222.760 31.760 223.435 31.920 ;
        RECT 223.895 31.840 225.115 32.010 ;
        RECT 222.760 30.970 222.970 31.760 ;
        RECT 223.895 31.750 224.065 31.840 ;
        RECT 223.140 30.970 223.490 31.590 ;
        RECT 223.660 31.580 224.065 31.750 ;
        RECT 223.660 30.800 223.830 31.580 ;
        RECT 224.000 31.130 224.220 31.410 ;
        RECT 224.400 31.300 224.940 31.670 ;
        RECT 225.285 31.590 225.455 32.180 ;
        RECT 225.675 31.760 225.980 32.900 ;
        RECT 226.150 31.710 226.405 32.590 ;
        RECT 226.580 31.735 226.870 32.900 ;
        RECT 225.285 31.560 226.025 31.590 ;
        RECT 224.000 30.960 224.530 31.130 ;
        RECT 222.310 30.540 222.660 30.710 ;
        RECT 222.880 30.520 223.830 30.800 ;
        RECT 224.000 30.350 224.190 30.790 ;
        RECT 224.360 30.730 224.530 30.960 ;
        RECT 224.700 30.900 224.940 31.300 ;
        RECT 225.110 31.260 226.025 31.560 ;
        RECT 225.110 31.085 225.435 31.260 ;
        RECT 225.110 30.730 225.430 31.085 ;
        RECT 226.195 31.060 226.405 31.710 ;
        RECT 227.045 31.710 227.300 32.590 ;
        RECT 227.470 31.760 227.775 32.900 ;
        RECT 228.115 32.520 228.445 32.900 ;
        RECT 228.625 32.350 228.795 32.640 ;
        RECT 228.965 32.440 229.215 32.900 ;
        RECT 227.995 32.180 228.795 32.350 ;
        RECT 229.385 32.390 230.255 32.730 ;
        RECT 224.360 30.560 225.430 30.730 ;
        RECT 225.675 30.350 225.980 30.810 ;
        RECT 226.150 30.530 226.405 31.060 ;
        RECT 226.580 30.350 226.870 31.075 ;
        RECT 227.045 31.060 227.255 31.710 ;
        RECT 227.995 31.590 228.165 32.180 ;
        RECT 229.385 32.010 229.555 32.390 ;
        RECT 230.490 32.270 230.660 32.730 ;
        RECT 230.830 32.440 231.200 32.900 ;
        RECT 231.495 32.300 231.665 32.640 ;
        RECT 231.835 32.470 232.165 32.900 ;
        RECT 232.400 32.300 232.570 32.640 ;
        RECT 228.335 31.840 229.555 32.010 ;
        RECT 229.725 31.930 230.185 32.220 ;
        RECT 230.490 32.100 231.050 32.270 ;
        RECT 231.495 32.130 232.570 32.300 ;
        RECT 232.740 32.400 233.420 32.730 ;
        RECT 233.635 32.400 233.885 32.730 ;
        RECT 234.055 32.440 234.305 32.900 ;
        RECT 230.880 31.960 231.050 32.100 ;
        RECT 229.725 31.920 230.690 31.930 ;
        RECT 229.385 31.750 229.555 31.840 ;
        RECT 230.015 31.760 230.690 31.920 ;
        RECT 227.425 31.560 228.165 31.590 ;
        RECT 227.425 31.260 228.340 31.560 ;
        RECT 228.015 31.085 228.340 31.260 ;
        RECT 227.045 30.530 227.300 31.060 ;
        RECT 227.470 30.350 227.775 30.810 ;
        RECT 228.020 30.730 228.340 31.085 ;
        RECT 228.510 31.300 229.050 31.670 ;
        RECT 229.385 31.580 229.790 31.750 ;
        RECT 228.510 30.900 228.750 31.300 ;
        RECT 229.230 31.130 229.450 31.410 ;
        RECT 228.920 30.960 229.450 31.130 ;
        RECT 228.920 30.730 229.090 30.960 ;
        RECT 229.620 30.800 229.790 31.580 ;
        RECT 229.960 30.970 230.310 31.590 ;
        RECT 230.480 30.970 230.690 31.760 ;
        RECT 230.880 31.790 232.380 31.960 ;
        RECT 230.880 31.100 231.050 31.790 ;
        RECT 232.740 31.620 232.910 32.400 ;
        RECT 233.715 32.270 233.885 32.400 ;
        RECT 231.220 31.450 232.910 31.620 ;
        RECT 233.080 31.840 233.545 32.230 ;
        RECT 233.715 32.100 234.110 32.270 ;
        RECT 231.220 31.270 231.390 31.450 ;
        RECT 228.020 30.560 229.090 30.730 ;
        RECT 229.260 30.350 229.450 30.790 ;
        RECT 229.620 30.520 230.570 30.800 ;
        RECT 230.880 30.710 231.140 31.100 ;
        RECT 231.560 31.030 232.350 31.280 ;
        RECT 230.790 30.540 231.140 30.710 ;
        RECT 231.350 30.350 231.680 30.810 ;
        RECT 232.555 30.740 232.725 31.450 ;
        RECT 233.080 31.250 233.250 31.840 ;
        RECT 232.895 31.030 233.250 31.250 ;
        RECT 233.420 31.030 233.770 31.650 ;
        RECT 233.940 30.740 234.110 32.100 ;
        RECT 234.475 31.930 234.800 32.715 ;
        RECT 234.280 30.880 234.740 31.930 ;
        RECT 232.555 30.570 233.410 30.740 ;
        RECT 233.615 30.570 234.110 30.740 ;
        RECT 234.280 30.350 234.610 30.710 ;
        RECT 234.970 30.610 235.140 32.730 ;
        RECT 235.310 32.400 235.640 32.900 ;
        RECT 235.810 32.230 236.065 32.730 ;
        RECT 235.315 32.060 236.065 32.230 ;
        RECT 235.315 31.070 235.545 32.060 ;
        RECT 236.295 32.030 236.580 32.900 ;
        RECT 236.750 32.270 237.010 32.730 ;
        RECT 237.185 32.440 237.440 32.900 ;
        RECT 237.610 32.270 237.870 32.730 ;
        RECT 236.750 32.100 237.870 32.270 ;
        RECT 238.040 32.100 238.350 32.900 ;
        RECT 235.715 31.240 236.065 31.890 ;
        RECT 236.750 31.850 237.010 32.100 ;
        RECT 238.520 31.930 238.830 32.730 ;
        RECT 236.255 31.680 237.010 31.850 ;
        RECT 237.800 31.760 238.830 31.930 ;
        RECT 239.000 31.810 242.510 32.900 ;
        RECT 242.680 31.810 243.890 32.900 ;
        RECT 236.255 31.170 236.660 31.680 ;
        RECT 237.800 31.510 237.970 31.760 ;
        RECT 236.830 31.340 237.970 31.510 ;
        RECT 235.315 30.900 236.065 31.070 ;
        RECT 236.255 31.000 237.905 31.170 ;
        RECT 238.140 31.020 238.490 31.590 ;
        RECT 235.310 30.350 235.640 30.730 ;
        RECT 235.810 30.610 236.065 30.900 ;
        RECT 236.300 30.350 236.580 30.830 ;
        RECT 236.750 30.610 237.010 31.000 ;
        RECT 237.185 30.350 237.440 30.830 ;
        RECT 237.610 30.610 237.905 31.000 ;
        RECT 238.660 30.850 238.830 31.760 ;
        RECT 238.085 30.350 238.360 30.830 ;
        RECT 238.530 30.520 238.830 30.850 ;
        RECT 239.000 31.120 240.650 31.640 ;
        RECT 240.820 31.290 242.510 31.810 ;
        RECT 239.000 30.350 242.510 31.120 ;
        RECT 242.680 31.100 243.200 31.640 ;
        RECT 243.370 31.270 243.890 31.810 ;
        RECT 244.060 31.825 244.330 32.730 ;
        RECT 244.500 32.140 244.830 32.900 ;
        RECT 245.010 31.970 245.180 32.730 ;
        RECT 242.680 30.350 243.890 31.100 ;
        RECT 244.060 31.025 244.230 31.825 ;
        RECT 244.515 31.800 245.180 31.970 ;
        RECT 244.515 31.655 244.685 31.800 ;
        RECT 244.400 31.325 244.685 31.655 ;
        RECT 245.445 31.760 245.780 32.730 ;
        RECT 245.950 31.760 246.120 32.900 ;
        RECT 246.290 32.560 248.320 32.730 ;
        RECT 244.515 31.070 244.685 31.325 ;
        RECT 244.920 31.250 245.250 31.620 ;
        RECT 245.445 31.090 245.615 31.760 ;
        RECT 246.290 31.590 246.460 32.560 ;
        RECT 245.785 31.260 246.040 31.590 ;
        RECT 246.265 31.260 246.460 31.590 ;
        RECT 246.630 32.220 247.755 32.390 ;
        RECT 245.870 31.090 246.040 31.260 ;
        RECT 246.630 31.090 246.800 32.220 ;
        RECT 244.060 30.520 244.320 31.025 ;
        RECT 244.515 30.900 245.180 31.070 ;
        RECT 244.500 30.350 244.830 30.730 ;
        RECT 245.010 30.520 245.180 30.900 ;
        RECT 245.445 30.520 245.700 31.090 ;
        RECT 245.870 30.920 246.800 31.090 ;
        RECT 246.970 31.880 247.980 32.050 ;
        RECT 246.970 31.080 247.140 31.880 ;
        RECT 247.345 31.200 247.620 31.680 ;
        RECT 247.340 31.030 247.620 31.200 ;
        RECT 246.625 30.885 246.800 30.920 ;
        RECT 245.870 30.350 246.200 30.750 ;
        RECT 246.625 30.520 247.155 30.885 ;
        RECT 247.345 30.520 247.620 31.030 ;
        RECT 247.790 30.520 247.980 31.880 ;
        RECT 248.150 31.895 248.320 32.560 ;
        RECT 248.490 32.140 248.660 32.900 ;
        RECT 248.895 32.140 249.410 32.550 ;
        RECT 248.150 31.705 248.900 31.895 ;
        RECT 249.070 31.330 249.410 32.140 ;
        RECT 249.580 31.810 252.170 32.900 ;
        RECT 248.180 31.160 249.410 31.330 ;
        RECT 248.160 30.350 248.670 30.885 ;
        RECT 248.890 30.555 249.135 31.160 ;
        RECT 249.580 31.120 250.790 31.640 ;
        RECT 250.960 31.290 252.170 31.810 ;
        RECT 252.340 31.735 252.630 32.900 ;
        RECT 252.800 31.810 255.390 32.900 ;
        RECT 256.075 32.030 256.360 32.900 ;
        RECT 256.530 32.270 256.790 32.730 ;
        RECT 256.965 32.440 257.220 32.900 ;
        RECT 257.390 32.270 257.650 32.730 ;
        RECT 256.530 32.100 257.650 32.270 ;
        RECT 257.820 32.100 258.130 32.900 ;
        RECT 256.530 31.850 256.790 32.100 ;
        RECT 258.300 31.930 258.610 32.730 ;
        RECT 252.800 31.120 254.010 31.640 ;
        RECT 254.180 31.290 255.390 31.810 ;
        RECT 256.035 31.680 256.790 31.850 ;
        RECT 257.580 31.760 258.610 31.930 ;
        RECT 256.035 31.170 256.440 31.680 ;
        RECT 257.580 31.510 257.750 31.760 ;
        RECT 256.610 31.340 257.750 31.510 ;
        RECT 249.580 30.350 252.170 31.120 ;
        RECT 252.340 30.350 252.630 31.075 ;
        RECT 252.800 30.350 255.390 31.120 ;
        RECT 256.035 31.000 257.685 31.170 ;
        RECT 257.920 31.020 258.270 31.590 ;
        RECT 256.080 30.350 256.360 30.830 ;
        RECT 256.530 30.610 256.790 31.000 ;
        RECT 256.965 30.350 257.220 30.830 ;
        RECT 257.390 30.610 257.685 31.000 ;
        RECT 258.440 30.850 258.610 31.760 ;
        RECT 257.865 30.350 258.140 30.830 ;
        RECT 258.310 30.520 258.610 30.850 ;
        RECT 258.815 32.110 259.350 32.730 ;
        RECT 258.815 31.090 259.130 32.110 ;
        RECT 259.520 32.100 259.850 32.900 ;
        RECT 260.335 31.930 260.725 32.105 ;
        RECT 259.300 31.760 260.725 31.930 ;
        RECT 261.080 31.810 264.590 32.900 ;
        RECT 259.300 31.260 259.470 31.760 ;
        RECT 258.815 30.520 259.430 31.090 ;
        RECT 259.720 31.030 259.985 31.590 ;
        RECT 260.155 30.860 260.325 31.760 ;
        RECT 260.495 31.030 260.850 31.590 ;
        RECT 261.080 31.120 262.730 31.640 ;
        RECT 262.900 31.290 264.590 31.810 ;
        RECT 265.225 31.710 265.480 32.590 ;
        RECT 265.650 31.760 265.955 32.900 ;
        RECT 266.295 32.520 266.625 32.900 ;
        RECT 266.805 32.350 266.975 32.640 ;
        RECT 267.145 32.440 267.395 32.900 ;
        RECT 266.175 32.180 266.975 32.350 ;
        RECT 267.565 32.390 268.435 32.730 ;
        RECT 259.600 30.350 259.815 30.860 ;
        RECT 260.045 30.530 260.325 30.860 ;
        RECT 260.505 30.350 260.745 30.860 ;
        RECT 261.080 30.350 264.590 31.120 ;
        RECT 265.225 31.060 265.435 31.710 ;
        RECT 266.175 31.590 266.345 32.180 ;
        RECT 267.565 32.010 267.735 32.390 ;
        RECT 268.670 32.270 268.840 32.730 ;
        RECT 269.010 32.440 269.380 32.900 ;
        RECT 269.675 32.300 269.845 32.640 ;
        RECT 270.015 32.470 270.345 32.900 ;
        RECT 270.580 32.300 270.750 32.640 ;
        RECT 266.515 31.840 267.735 32.010 ;
        RECT 267.905 31.930 268.365 32.220 ;
        RECT 268.670 32.100 269.230 32.270 ;
        RECT 269.675 32.130 270.750 32.300 ;
        RECT 270.920 32.400 271.600 32.730 ;
        RECT 271.815 32.400 272.065 32.730 ;
        RECT 272.235 32.440 272.485 32.900 ;
        RECT 269.060 31.960 269.230 32.100 ;
        RECT 267.905 31.920 268.870 31.930 ;
        RECT 267.565 31.750 267.735 31.840 ;
        RECT 268.195 31.760 268.870 31.920 ;
        RECT 265.605 31.560 266.345 31.590 ;
        RECT 265.605 31.260 266.520 31.560 ;
        RECT 266.195 31.085 266.520 31.260 ;
        RECT 265.225 30.530 265.480 31.060 ;
        RECT 265.650 30.350 265.955 30.810 ;
        RECT 266.200 30.730 266.520 31.085 ;
        RECT 266.690 31.300 267.230 31.670 ;
        RECT 267.565 31.580 267.970 31.750 ;
        RECT 266.690 30.900 266.930 31.300 ;
        RECT 267.410 31.130 267.630 31.410 ;
        RECT 267.100 30.960 267.630 31.130 ;
        RECT 267.100 30.730 267.270 30.960 ;
        RECT 267.800 30.800 267.970 31.580 ;
        RECT 268.140 30.970 268.490 31.590 ;
        RECT 268.660 30.970 268.870 31.760 ;
        RECT 269.060 31.790 270.560 31.960 ;
        RECT 269.060 31.100 269.230 31.790 ;
        RECT 270.920 31.620 271.090 32.400 ;
        RECT 271.895 32.270 272.065 32.400 ;
        RECT 269.400 31.450 271.090 31.620 ;
        RECT 271.260 31.840 271.725 32.230 ;
        RECT 271.895 32.100 272.290 32.270 ;
        RECT 269.400 31.270 269.570 31.450 ;
        RECT 266.200 30.560 267.270 30.730 ;
        RECT 267.440 30.350 267.630 30.790 ;
        RECT 267.800 30.520 268.750 30.800 ;
        RECT 269.060 30.710 269.320 31.100 ;
        RECT 269.740 31.030 270.530 31.280 ;
        RECT 268.970 30.540 269.320 30.710 ;
        RECT 269.530 30.350 269.860 30.810 ;
        RECT 270.735 30.740 270.905 31.450 ;
        RECT 271.260 31.250 271.430 31.840 ;
        RECT 271.075 31.030 271.430 31.250 ;
        RECT 271.600 31.030 271.950 31.650 ;
        RECT 272.120 30.740 272.290 32.100 ;
        RECT 272.655 31.930 272.980 32.715 ;
        RECT 272.460 30.880 272.920 31.930 ;
        RECT 270.735 30.570 271.590 30.740 ;
        RECT 271.795 30.570 272.290 30.740 ;
        RECT 272.460 30.350 272.790 30.710 ;
        RECT 273.150 30.610 273.320 32.730 ;
        RECT 273.490 32.400 273.820 32.900 ;
        RECT 273.990 32.230 274.245 32.730 ;
        RECT 273.495 32.060 274.245 32.230 ;
        RECT 274.535 32.270 274.820 32.730 ;
        RECT 274.990 32.440 275.260 32.900 ;
        RECT 273.495 31.070 273.725 32.060 ;
        RECT 274.535 32.050 275.490 32.270 ;
        RECT 273.895 31.240 274.245 31.890 ;
        RECT 274.420 31.320 275.110 31.880 ;
        RECT 275.280 31.150 275.490 32.050 ;
        RECT 273.495 30.900 274.245 31.070 ;
        RECT 273.490 30.350 273.820 30.730 ;
        RECT 273.990 30.610 274.245 30.900 ;
        RECT 274.535 30.980 275.490 31.150 ;
        RECT 275.660 31.880 276.060 32.730 ;
        RECT 276.250 32.270 276.530 32.730 ;
        RECT 277.050 32.440 277.375 32.900 ;
        RECT 276.250 32.050 277.375 32.270 ;
        RECT 275.660 31.320 276.755 31.880 ;
        RECT 276.925 31.590 277.375 32.050 ;
        RECT 277.545 31.760 277.930 32.730 ;
        RECT 274.535 30.520 274.820 30.980 ;
        RECT 274.990 30.350 275.260 30.810 ;
        RECT 275.660 30.520 276.060 31.320 ;
        RECT 276.925 31.260 277.480 31.590 ;
        RECT 276.925 31.150 277.375 31.260 ;
        RECT 276.250 30.980 277.375 31.150 ;
        RECT 277.650 31.090 277.930 31.760 ;
        RECT 278.100 31.735 278.390 32.900 ;
        RECT 278.565 31.760 278.900 32.730 ;
        RECT 279.070 31.760 279.240 32.900 ;
        RECT 279.410 32.560 281.440 32.730 ;
        RECT 276.250 30.520 276.530 30.980 ;
        RECT 277.050 30.350 277.375 30.810 ;
        RECT 277.545 30.520 277.930 31.090 ;
        RECT 278.565 31.090 278.735 31.760 ;
        RECT 279.410 31.590 279.580 32.560 ;
        RECT 278.905 31.260 279.160 31.590 ;
        RECT 279.385 31.260 279.580 31.590 ;
        RECT 279.750 32.220 280.875 32.390 ;
        RECT 278.990 31.090 279.160 31.260 ;
        RECT 279.750 31.090 279.920 32.220 ;
        RECT 278.100 30.350 278.390 31.075 ;
        RECT 278.565 30.520 278.820 31.090 ;
        RECT 278.990 30.920 279.920 31.090 ;
        RECT 280.090 31.880 281.100 32.050 ;
        RECT 280.090 31.080 280.260 31.880 ;
        RECT 280.465 31.200 280.740 31.680 ;
        RECT 280.460 31.030 280.740 31.200 ;
        RECT 279.745 30.885 279.920 30.920 ;
        RECT 278.990 30.350 279.320 30.750 ;
        RECT 279.745 30.520 280.275 30.885 ;
        RECT 280.465 30.520 280.740 31.030 ;
        RECT 280.910 30.520 281.100 31.880 ;
        RECT 281.270 31.895 281.440 32.560 ;
        RECT 281.610 32.140 281.780 32.900 ;
        RECT 282.015 32.140 282.530 32.550 ;
        RECT 281.270 31.705 282.020 31.895 ;
        RECT 282.190 31.330 282.530 32.140 ;
        RECT 282.700 31.760 282.960 32.900 ;
        RECT 283.130 31.750 283.460 32.730 ;
        RECT 283.630 31.760 283.910 32.900 ;
        RECT 284.080 31.810 285.290 32.900 ;
        RECT 282.720 31.340 283.055 31.590 ;
        RECT 281.300 31.160 282.530 31.330 ;
        RECT 281.280 30.350 281.790 30.885 ;
        RECT 282.010 30.555 282.255 31.160 ;
        RECT 283.225 31.150 283.395 31.750 ;
        RECT 283.565 31.320 283.900 31.590 ;
        RECT 282.700 30.520 283.395 31.150 ;
        RECT 283.600 30.350 283.910 31.150 ;
        RECT 284.080 31.100 284.600 31.640 ;
        RECT 284.770 31.270 285.290 31.810 ;
        RECT 285.465 31.710 285.720 32.590 ;
        RECT 285.890 31.760 286.195 32.900 ;
        RECT 286.535 32.520 286.865 32.900 ;
        RECT 287.045 32.350 287.215 32.640 ;
        RECT 287.385 32.440 287.635 32.900 ;
        RECT 286.415 32.180 287.215 32.350 ;
        RECT 287.805 32.390 288.675 32.730 ;
        RECT 284.080 30.350 285.290 31.100 ;
        RECT 285.465 31.060 285.675 31.710 ;
        RECT 286.415 31.590 286.585 32.180 ;
        RECT 287.805 32.010 287.975 32.390 ;
        RECT 288.910 32.270 289.080 32.730 ;
        RECT 289.250 32.440 289.620 32.900 ;
        RECT 289.915 32.300 290.085 32.640 ;
        RECT 290.255 32.470 290.585 32.900 ;
        RECT 290.820 32.300 290.990 32.640 ;
        RECT 286.755 31.840 287.975 32.010 ;
        RECT 288.145 31.930 288.605 32.220 ;
        RECT 288.910 32.100 289.470 32.270 ;
        RECT 289.915 32.130 290.990 32.300 ;
        RECT 291.160 32.400 291.840 32.730 ;
        RECT 292.055 32.400 292.305 32.730 ;
        RECT 292.475 32.440 292.725 32.900 ;
        RECT 289.300 31.960 289.470 32.100 ;
        RECT 288.145 31.920 289.110 31.930 ;
        RECT 287.805 31.750 287.975 31.840 ;
        RECT 288.435 31.760 289.110 31.920 ;
        RECT 285.845 31.560 286.585 31.590 ;
        RECT 285.845 31.260 286.760 31.560 ;
        RECT 286.435 31.085 286.760 31.260 ;
        RECT 285.465 30.530 285.720 31.060 ;
        RECT 285.890 30.350 286.195 30.810 ;
        RECT 286.440 30.730 286.760 31.085 ;
        RECT 286.930 31.300 287.470 31.670 ;
        RECT 287.805 31.580 288.210 31.750 ;
        RECT 286.930 30.900 287.170 31.300 ;
        RECT 287.650 31.130 287.870 31.410 ;
        RECT 287.340 30.960 287.870 31.130 ;
        RECT 287.340 30.730 287.510 30.960 ;
        RECT 288.040 30.800 288.210 31.580 ;
        RECT 288.380 30.970 288.730 31.590 ;
        RECT 288.900 30.970 289.110 31.760 ;
        RECT 289.300 31.790 290.800 31.960 ;
        RECT 289.300 31.100 289.470 31.790 ;
        RECT 291.160 31.620 291.330 32.400 ;
        RECT 292.135 32.270 292.305 32.400 ;
        RECT 289.640 31.450 291.330 31.620 ;
        RECT 291.500 31.840 291.965 32.230 ;
        RECT 292.135 32.100 292.530 32.270 ;
        RECT 289.640 31.270 289.810 31.450 ;
        RECT 286.440 30.560 287.510 30.730 ;
        RECT 287.680 30.350 287.870 30.790 ;
        RECT 288.040 30.520 288.990 30.800 ;
        RECT 289.300 30.710 289.560 31.100 ;
        RECT 289.980 31.030 290.770 31.280 ;
        RECT 289.210 30.540 289.560 30.710 ;
        RECT 289.770 30.350 290.100 30.810 ;
        RECT 290.975 30.740 291.145 31.450 ;
        RECT 291.500 31.250 291.670 31.840 ;
        RECT 291.315 31.030 291.670 31.250 ;
        RECT 291.840 31.030 292.190 31.650 ;
        RECT 292.360 30.740 292.530 32.100 ;
        RECT 292.895 31.930 293.220 32.715 ;
        RECT 292.700 30.880 293.160 31.930 ;
        RECT 290.975 30.570 291.830 30.740 ;
        RECT 292.035 30.570 292.530 30.740 ;
        RECT 292.700 30.350 293.030 30.710 ;
        RECT 293.390 30.610 293.560 32.730 ;
        RECT 293.730 32.400 294.060 32.900 ;
        RECT 294.230 32.230 294.485 32.730 ;
        RECT 293.735 32.060 294.485 32.230 ;
        RECT 293.735 31.070 293.965 32.060 ;
        RECT 294.135 31.240 294.485 31.890 ;
        RECT 294.665 31.710 294.920 32.590 ;
        RECT 295.090 31.760 295.395 32.900 ;
        RECT 295.735 32.520 296.065 32.900 ;
        RECT 296.245 32.350 296.415 32.640 ;
        RECT 296.585 32.440 296.835 32.900 ;
        RECT 295.615 32.180 296.415 32.350 ;
        RECT 297.005 32.390 297.875 32.730 ;
        RECT 293.735 30.900 294.485 31.070 ;
        RECT 293.730 30.350 294.060 30.730 ;
        RECT 294.230 30.610 294.485 30.900 ;
        RECT 294.665 31.060 294.875 31.710 ;
        RECT 295.615 31.590 295.785 32.180 ;
        RECT 297.005 32.010 297.175 32.390 ;
        RECT 298.110 32.270 298.280 32.730 ;
        RECT 298.450 32.440 298.820 32.900 ;
        RECT 299.115 32.300 299.285 32.640 ;
        RECT 299.455 32.470 299.785 32.900 ;
        RECT 300.020 32.300 300.190 32.640 ;
        RECT 295.955 31.840 297.175 32.010 ;
        RECT 297.345 31.930 297.805 32.220 ;
        RECT 298.110 32.100 298.670 32.270 ;
        RECT 299.115 32.130 300.190 32.300 ;
        RECT 300.360 32.400 301.040 32.730 ;
        RECT 301.255 32.400 301.505 32.730 ;
        RECT 301.675 32.440 301.925 32.900 ;
        RECT 298.500 31.960 298.670 32.100 ;
        RECT 297.345 31.920 298.310 31.930 ;
        RECT 297.005 31.750 297.175 31.840 ;
        RECT 297.635 31.760 298.310 31.920 ;
        RECT 295.045 31.560 295.785 31.590 ;
        RECT 295.045 31.260 295.960 31.560 ;
        RECT 295.635 31.085 295.960 31.260 ;
        RECT 294.665 30.530 294.920 31.060 ;
        RECT 295.090 30.350 295.395 30.810 ;
        RECT 295.640 30.730 295.960 31.085 ;
        RECT 296.130 31.300 296.670 31.670 ;
        RECT 297.005 31.580 297.410 31.750 ;
        RECT 296.130 30.900 296.370 31.300 ;
        RECT 296.850 31.130 297.070 31.410 ;
        RECT 296.540 30.960 297.070 31.130 ;
        RECT 296.540 30.730 296.710 30.960 ;
        RECT 297.240 30.800 297.410 31.580 ;
        RECT 297.580 30.970 297.930 31.590 ;
        RECT 298.100 30.970 298.310 31.760 ;
        RECT 298.500 31.790 300.000 31.960 ;
        RECT 298.500 31.100 298.670 31.790 ;
        RECT 300.360 31.620 300.530 32.400 ;
        RECT 301.335 32.270 301.505 32.400 ;
        RECT 298.840 31.450 300.530 31.620 ;
        RECT 300.700 31.840 301.165 32.230 ;
        RECT 301.335 32.100 301.730 32.270 ;
        RECT 298.840 31.270 299.010 31.450 ;
        RECT 295.640 30.560 296.710 30.730 ;
        RECT 296.880 30.350 297.070 30.790 ;
        RECT 297.240 30.520 298.190 30.800 ;
        RECT 298.500 30.710 298.760 31.100 ;
        RECT 299.180 31.030 299.970 31.280 ;
        RECT 298.410 30.540 298.760 30.710 ;
        RECT 298.970 30.350 299.300 30.810 ;
        RECT 300.175 30.740 300.345 31.450 ;
        RECT 300.700 31.250 300.870 31.840 ;
        RECT 300.515 31.030 300.870 31.250 ;
        RECT 301.040 31.030 301.390 31.650 ;
        RECT 301.560 30.740 301.730 32.100 ;
        RECT 302.095 31.930 302.420 32.715 ;
        RECT 301.900 30.880 302.360 31.930 ;
        RECT 300.175 30.570 301.030 30.740 ;
        RECT 301.235 30.570 301.730 30.740 ;
        RECT 301.900 30.350 302.230 30.710 ;
        RECT 302.590 30.610 302.760 32.730 ;
        RECT 302.930 32.400 303.260 32.900 ;
        RECT 303.430 32.230 303.685 32.730 ;
        RECT 302.935 32.060 303.685 32.230 ;
        RECT 302.935 31.070 303.165 32.060 ;
        RECT 303.335 31.240 303.685 31.890 ;
        RECT 303.860 31.735 304.150 32.900 ;
        RECT 304.320 31.760 304.705 32.730 ;
        RECT 304.875 32.440 305.200 32.900 ;
        RECT 305.720 32.270 306.000 32.730 ;
        RECT 304.875 32.050 306.000 32.270 ;
        RECT 304.320 31.090 304.600 31.760 ;
        RECT 304.875 31.590 305.325 32.050 ;
        RECT 306.190 31.880 306.590 32.730 ;
        RECT 306.990 32.440 307.260 32.900 ;
        RECT 307.430 32.270 307.715 32.730 ;
        RECT 304.770 31.260 305.325 31.590 ;
        RECT 305.495 31.320 306.590 31.880 ;
        RECT 304.875 31.150 305.325 31.260 ;
        RECT 302.935 30.900 303.685 31.070 ;
        RECT 302.930 30.350 303.260 30.730 ;
        RECT 303.430 30.610 303.685 30.900 ;
        RECT 303.860 30.350 304.150 31.075 ;
        RECT 304.320 30.520 304.705 31.090 ;
        RECT 304.875 30.980 306.000 31.150 ;
        RECT 304.875 30.350 305.200 30.810 ;
        RECT 305.720 30.520 306.000 30.980 ;
        RECT 306.190 30.520 306.590 31.320 ;
        RECT 306.760 32.050 307.715 32.270 ;
        RECT 306.760 31.150 306.970 32.050 ;
        RECT 307.140 31.320 307.830 31.880 ;
        RECT 308.000 31.810 309.670 32.900 ;
        RECT 306.760 30.980 307.715 31.150 ;
        RECT 306.990 30.350 307.260 30.810 ;
        RECT 307.430 30.520 307.715 30.980 ;
        RECT 308.000 31.120 308.750 31.640 ;
        RECT 308.920 31.290 309.670 31.810 ;
        RECT 309.840 31.810 311.050 32.900 ;
        RECT 309.840 31.270 310.360 31.810 ;
        RECT 308.000 30.350 309.670 31.120 ;
        RECT 310.530 31.100 311.050 31.640 ;
        RECT 309.840 30.350 311.050 31.100 ;
        RECT 162.095 30.180 311.135 30.350 ;
        RECT 162.180 29.430 163.390 30.180 ;
        RECT 162.180 28.890 162.700 29.430 ;
        RECT 163.565 29.340 163.825 30.180 ;
        RECT 164.000 29.435 164.255 30.010 ;
        RECT 164.425 29.800 164.755 30.180 ;
        RECT 164.970 29.630 165.140 30.010 ;
        RECT 165.400 29.635 170.745 30.180 ;
        RECT 170.920 29.635 176.265 30.180 ;
        RECT 176.440 29.635 181.785 30.180 ;
        RECT 164.425 29.460 165.140 29.630 ;
        RECT 162.870 28.720 163.390 29.260 ;
        RECT 162.180 27.630 163.390 28.720 ;
        RECT 163.565 27.630 163.825 28.780 ;
        RECT 164.000 28.705 164.170 29.435 ;
        RECT 164.425 29.270 164.595 29.460 ;
        RECT 164.340 28.940 164.595 29.270 ;
        RECT 164.425 28.730 164.595 28.940 ;
        RECT 164.875 28.910 165.230 29.280 ;
        RECT 166.985 28.805 167.325 29.635 ;
        RECT 164.000 27.800 164.255 28.705 ;
        RECT 164.425 28.560 165.140 28.730 ;
        RECT 164.425 27.630 164.755 28.390 ;
        RECT 164.970 27.800 165.140 28.560 ;
        RECT 168.805 28.065 169.155 29.315 ;
        RECT 172.505 28.805 172.845 29.635 ;
        RECT 174.325 28.065 174.675 29.315 ;
        RECT 178.025 28.805 178.365 29.635 ;
        RECT 181.960 29.410 185.470 30.180 ;
        RECT 186.190 29.630 186.360 30.010 ;
        RECT 186.540 29.800 186.870 30.180 ;
        RECT 186.190 29.460 186.855 29.630 ;
        RECT 187.050 29.505 187.310 30.010 ;
        RECT 179.845 28.065 180.195 29.315 ;
        RECT 181.960 28.890 183.610 29.410 ;
        RECT 183.780 28.720 185.470 29.240 ;
        RECT 186.120 28.910 186.450 29.280 ;
        RECT 186.685 29.205 186.855 29.460 ;
        RECT 186.685 28.875 186.970 29.205 ;
        RECT 186.685 28.730 186.855 28.875 ;
        RECT 165.400 27.630 170.745 28.065 ;
        RECT 170.920 27.630 176.265 28.065 ;
        RECT 176.440 27.630 181.785 28.065 ;
        RECT 181.960 27.630 185.470 28.720 ;
        RECT 186.190 28.560 186.855 28.730 ;
        RECT 187.140 28.705 187.310 29.505 ;
        RECT 187.940 29.455 188.230 30.180 ;
        RECT 188.400 29.410 191.910 30.180 ;
        RECT 188.400 28.890 190.050 29.410 ;
        RECT 192.355 29.370 192.600 29.975 ;
        RECT 192.820 29.645 193.330 30.180 ;
        RECT 186.190 27.800 186.360 28.560 ;
        RECT 186.540 27.630 186.870 28.390 ;
        RECT 187.040 27.800 187.310 28.705 ;
        RECT 187.940 27.630 188.230 28.795 ;
        RECT 190.220 28.720 191.910 29.240 ;
        RECT 188.400 27.630 191.910 28.720 ;
        RECT 192.080 29.200 193.310 29.370 ;
        RECT 192.080 28.390 192.420 29.200 ;
        RECT 192.590 28.635 193.340 28.825 ;
        RECT 192.080 27.980 192.595 28.390 ;
        RECT 192.830 27.630 193.000 28.390 ;
        RECT 193.170 27.970 193.340 28.635 ;
        RECT 193.510 28.650 193.700 30.010 ;
        RECT 193.870 29.160 194.145 30.010 ;
        RECT 194.335 29.645 194.865 30.010 ;
        RECT 195.290 29.780 195.620 30.180 ;
        RECT 194.690 29.610 194.865 29.645 ;
        RECT 193.870 28.990 194.150 29.160 ;
        RECT 193.870 28.850 194.145 28.990 ;
        RECT 194.350 28.650 194.520 29.450 ;
        RECT 193.510 28.480 194.520 28.650 ;
        RECT 194.690 29.440 195.620 29.610 ;
        RECT 195.790 29.440 196.045 30.010 ;
        RECT 194.690 28.310 194.860 29.440 ;
        RECT 195.450 29.270 195.620 29.440 ;
        RECT 193.735 28.140 194.860 28.310 ;
        RECT 195.030 28.940 195.225 29.270 ;
        RECT 195.450 28.940 195.705 29.270 ;
        RECT 195.030 27.970 195.200 28.940 ;
        RECT 195.875 28.770 196.045 29.440 ;
        RECT 196.220 29.410 198.810 30.180 ;
        RECT 198.985 29.630 199.240 29.920 ;
        RECT 199.410 29.800 199.740 30.180 ;
        RECT 198.985 29.460 199.735 29.630 ;
        RECT 196.220 28.890 197.430 29.410 ;
        RECT 193.170 27.800 195.200 27.970 ;
        RECT 195.370 27.630 195.540 28.770 ;
        RECT 195.710 27.800 196.045 28.770 ;
        RECT 197.600 28.720 198.810 29.240 ;
        RECT 196.220 27.630 198.810 28.720 ;
        RECT 198.985 28.640 199.335 29.290 ;
        RECT 199.505 28.470 199.735 29.460 ;
        RECT 198.985 28.300 199.735 28.470 ;
        RECT 198.985 27.800 199.240 28.300 ;
        RECT 199.410 27.630 199.740 28.130 ;
        RECT 199.910 27.800 200.080 29.920 ;
        RECT 200.440 29.820 200.770 30.180 ;
        RECT 200.940 29.790 201.435 29.960 ;
        RECT 201.640 29.790 202.495 29.960 ;
        RECT 200.310 28.600 200.770 29.650 ;
        RECT 200.250 27.815 200.575 28.600 ;
        RECT 200.940 28.430 201.110 29.790 ;
        RECT 201.280 28.880 201.630 29.500 ;
        RECT 201.800 29.280 202.155 29.500 ;
        RECT 201.800 28.690 201.970 29.280 ;
        RECT 202.325 29.080 202.495 29.790 ;
        RECT 203.370 29.720 203.700 30.180 ;
        RECT 203.910 29.820 204.260 29.990 ;
        RECT 202.700 29.250 203.490 29.500 ;
        RECT 203.910 29.430 204.170 29.820 ;
        RECT 204.480 29.730 205.430 30.010 ;
        RECT 205.600 29.740 205.790 30.180 ;
        RECT 205.960 29.800 207.030 29.970 ;
        RECT 203.660 29.080 203.830 29.260 ;
        RECT 200.940 28.260 201.335 28.430 ;
        RECT 201.505 28.300 201.970 28.690 ;
        RECT 202.140 28.910 203.830 29.080 ;
        RECT 201.165 28.130 201.335 28.260 ;
        RECT 202.140 28.130 202.310 28.910 ;
        RECT 204.000 28.740 204.170 29.430 ;
        RECT 202.670 28.570 204.170 28.740 ;
        RECT 204.360 28.770 204.570 29.560 ;
        RECT 204.740 28.940 205.090 29.560 ;
        RECT 205.260 28.950 205.430 29.730 ;
        RECT 205.960 29.570 206.130 29.800 ;
        RECT 205.600 29.400 206.130 29.570 ;
        RECT 205.600 29.120 205.820 29.400 ;
        RECT 206.300 29.230 206.540 29.630 ;
        RECT 205.260 28.780 205.665 28.950 ;
        RECT 206.000 28.860 206.540 29.230 ;
        RECT 206.710 29.445 207.030 29.800 ;
        RECT 207.275 29.720 207.580 30.180 ;
        RECT 207.750 29.470 208.005 30.000 ;
        RECT 206.710 29.270 207.035 29.445 ;
        RECT 206.710 28.970 207.625 29.270 ;
        RECT 206.885 28.940 207.625 28.970 ;
        RECT 204.360 28.610 205.035 28.770 ;
        RECT 205.495 28.690 205.665 28.780 ;
        RECT 204.360 28.600 205.325 28.610 ;
        RECT 204.000 28.430 204.170 28.570 ;
        RECT 200.745 27.630 200.995 28.090 ;
        RECT 201.165 27.800 201.415 28.130 ;
        RECT 201.630 27.800 202.310 28.130 ;
        RECT 202.480 28.230 203.555 28.400 ;
        RECT 204.000 28.260 204.560 28.430 ;
        RECT 204.865 28.310 205.325 28.600 ;
        RECT 205.495 28.520 206.715 28.690 ;
        RECT 202.480 27.890 202.650 28.230 ;
        RECT 202.885 27.630 203.215 28.060 ;
        RECT 203.385 27.890 203.555 28.230 ;
        RECT 203.850 27.630 204.220 28.090 ;
        RECT 204.390 27.800 204.560 28.260 ;
        RECT 205.495 28.140 205.665 28.520 ;
        RECT 206.885 28.350 207.055 28.940 ;
        RECT 207.795 28.820 208.005 29.470 ;
        RECT 209.375 29.370 209.620 29.975 ;
        RECT 209.840 29.645 210.350 30.180 ;
        RECT 204.795 27.800 205.665 28.140 ;
        RECT 206.255 28.180 207.055 28.350 ;
        RECT 205.835 27.630 206.085 28.090 ;
        RECT 206.255 27.890 206.425 28.180 ;
        RECT 206.605 27.630 206.935 28.010 ;
        RECT 207.275 27.630 207.580 28.770 ;
        RECT 207.750 27.940 208.005 28.820 ;
        RECT 209.100 29.200 210.330 29.370 ;
        RECT 209.100 28.390 209.440 29.200 ;
        RECT 209.610 28.635 210.360 28.825 ;
        RECT 209.100 27.980 209.615 28.390 ;
        RECT 209.850 27.630 210.020 28.390 ;
        RECT 210.190 27.970 210.360 28.635 ;
        RECT 210.530 28.650 210.720 30.010 ;
        RECT 210.890 29.500 211.165 30.010 ;
        RECT 211.355 29.645 211.885 30.010 ;
        RECT 212.310 29.780 212.640 30.180 ;
        RECT 211.710 29.610 211.885 29.645 ;
        RECT 210.890 29.330 211.170 29.500 ;
        RECT 210.890 28.850 211.165 29.330 ;
        RECT 211.370 28.650 211.540 29.450 ;
        RECT 210.530 28.480 211.540 28.650 ;
        RECT 211.710 29.440 212.640 29.610 ;
        RECT 212.810 29.440 213.065 30.010 ;
        RECT 213.700 29.455 213.990 30.180 ;
        RECT 214.165 29.630 214.420 29.920 ;
        RECT 214.590 29.800 214.920 30.180 ;
        RECT 214.165 29.460 214.915 29.630 ;
        RECT 211.710 28.310 211.880 29.440 ;
        RECT 212.470 29.270 212.640 29.440 ;
        RECT 210.755 28.140 211.880 28.310 ;
        RECT 212.050 28.940 212.245 29.270 ;
        RECT 212.470 28.940 212.725 29.270 ;
        RECT 212.050 27.970 212.220 28.940 ;
        RECT 212.895 28.770 213.065 29.440 ;
        RECT 210.190 27.800 212.220 27.970 ;
        RECT 212.390 27.630 212.560 28.770 ;
        RECT 212.730 27.800 213.065 28.770 ;
        RECT 213.700 27.630 213.990 28.795 ;
        RECT 214.165 28.640 214.515 29.290 ;
        RECT 214.685 28.470 214.915 29.460 ;
        RECT 214.165 28.300 214.915 28.470 ;
        RECT 214.165 27.800 214.420 28.300 ;
        RECT 214.590 27.630 214.920 28.130 ;
        RECT 215.090 27.800 215.260 29.920 ;
        RECT 215.620 29.820 215.950 30.180 ;
        RECT 216.120 29.790 216.615 29.960 ;
        RECT 216.820 29.790 217.675 29.960 ;
        RECT 215.490 28.600 215.950 29.650 ;
        RECT 215.430 27.815 215.755 28.600 ;
        RECT 216.120 28.430 216.290 29.790 ;
        RECT 216.460 28.880 216.810 29.500 ;
        RECT 216.980 29.280 217.335 29.500 ;
        RECT 216.980 28.690 217.150 29.280 ;
        RECT 217.505 29.080 217.675 29.790 ;
        RECT 218.550 29.720 218.880 30.180 ;
        RECT 219.090 29.820 219.440 29.990 ;
        RECT 217.880 29.250 218.670 29.500 ;
        RECT 219.090 29.430 219.350 29.820 ;
        RECT 219.660 29.730 220.610 30.010 ;
        RECT 220.780 29.740 220.970 30.180 ;
        RECT 221.140 29.800 222.210 29.970 ;
        RECT 218.840 29.080 219.010 29.260 ;
        RECT 216.120 28.260 216.515 28.430 ;
        RECT 216.685 28.300 217.150 28.690 ;
        RECT 217.320 28.910 219.010 29.080 ;
        RECT 216.345 28.130 216.515 28.260 ;
        RECT 217.320 28.130 217.490 28.910 ;
        RECT 219.180 28.740 219.350 29.430 ;
        RECT 217.850 28.570 219.350 28.740 ;
        RECT 219.540 28.770 219.750 29.560 ;
        RECT 219.920 28.940 220.270 29.560 ;
        RECT 220.440 28.950 220.610 29.730 ;
        RECT 221.140 29.570 221.310 29.800 ;
        RECT 220.780 29.400 221.310 29.570 ;
        RECT 220.780 29.120 221.000 29.400 ;
        RECT 221.480 29.230 221.720 29.630 ;
        RECT 220.440 28.780 220.845 28.950 ;
        RECT 221.180 28.860 221.720 29.230 ;
        RECT 221.890 29.445 222.210 29.800 ;
        RECT 222.455 29.720 222.760 30.180 ;
        RECT 222.930 29.470 223.185 30.000 ;
        RECT 223.360 29.635 228.705 30.180 ;
        RECT 221.890 29.270 222.215 29.445 ;
        RECT 221.890 28.970 222.805 29.270 ;
        RECT 222.065 28.940 222.805 28.970 ;
        RECT 219.540 28.610 220.215 28.770 ;
        RECT 220.675 28.690 220.845 28.780 ;
        RECT 219.540 28.600 220.505 28.610 ;
        RECT 219.180 28.430 219.350 28.570 ;
        RECT 215.925 27.630 216.175 28.090 ;
        RECT 216.345 27.800 216.595 28.130 ;
        RECT 216.810 27.800 217.490 28.130 ;
        RECT 217.660 28.230 218.735 28.400 ;
        RECT 219.180 28.260 219.740 28.430 ;
        RECT 220.045 28.310 220.505 28.600 ;
        RECT 220.675 28.520 221.895 28.690 ;
        RECT 217.660 27.890 217.830 28.230 ;
        RECT 218.065 27.630 218.395 28.060 ;
        RECT 218.565 27.890 218.735 28.230 ;
        RECT 219.030 27.630 219.400 28.090 ;
        RECT 219.570 27.800 219.740 28.260 ;
        RECT 220.675 28.140 220.845 28.520 ;
        RECT 222.065 28.350 222.235 28.940 ;
        RECT 222.975 28.820 223.185 29.470 ;
        RECT 219.975 27.800 220.845 28.140 ;
        RECT 221.435 28.180 222.235 28.350 ;
        RECT 221.015 27.630 221.265 28.090 ;
        RECT 221.435 27.890 221.605 28.180 ;
        RECT 221.785 27.630 222.115 28.010 ;
        RECT 222.455 27.630 222.760 28.770 ;
        RECT 222.930 27.940 223.185 28.820 ;
        RECT 224.945 28.805 225.285 29.635 ;
        RECT 229.890 29.630 230.060 30.010 ;
        RECT 230.240 29.800 230.570 30.180 ;
        RECT 229.890 29.460 230.555 29.630 ;
        RECT 230.750 29.505 231.010 30.010 ;
        RECT 226.765 28.065 227.115 29.315 ;
        RECT 229.820 28.910 230.150 29.280 ;
        RECT 230.385 29.205 230.555 29.460 ;
        RECT 230.385 28.875 230.670 29.205 ;
        RECT 230.385 28.730 230.555 28.875 ;
        RECT 229.890 28.560 230.555 28.730 ;
        RECT 230.840 28.705 231.010 29.505 ;
        RECT 223.360 27.630 228.705 28.065 ;
        RECT 229.890 27.800 230.060 28.560 ;
        RECT 230.240 27.630 230.570 28.390 ;
        RECT 230.740 27.800 231.010 28.705 ;
        RECT 231.645 29.440 231.900 30.010 ;
        RECT 232.070 29.780 232.400 30.180 ;
        RECT 232.825 29.645 233.355 30.010 ;
        RECT 233.545 29.840 233.820 30.010 ;
        RECT 233.540 29.670 233.820 29.840 ;
        RECT 232.825 29.610 233.000 29.645 ;
        RECT 232.070 29.440 233.000 29.610 ;
        RECT 231.645 28.770 231.815 29.440 ;
        RECT 232.070 29.270 232.240 29.440 ;
        RECT 231.985 28.940 232.240 29.270 ;
        RECT 232.465 28.940 232.660 29.270 ;
        RECT 231.645 27.800 231.980 28.770 ;
        RECT 232.150 27.630 232.320 28.770 ;
        RECT 232.490 27.970 232.660 28.940 ;
        RECT 232.830 28.310 233.000 29.440 ;
        RECT 233.170 28.650 233.340 29.450 ;
        RECT 233.545 28.850 233.820 29.670 ;
        RECT 233.990 28.650 234.180 30.010 ;
        RECT 234.360 29.645 234.870 30.180 ;
        RECT 235.090 29.370 235.335 29.975 ;
        RECT 235.780 29.410 239.290 30.180 ;
        RECT 239.460 29.455 239.750 30.180 ;
        RECT 239.920 29.635 245.265 30.180 ;
        RECT 245.440 29.635 250.785 30.180 ;
        RECT 250.960 29.635 256.305 30.180 ;
        RECT 256.480 29.635 261.825 30.180 ;
        RECT 234.380 29.200 235.610 29.370 ;
        RECT 233.170 28.480 234.180 28.650 ;
        RECT 234.350 28.635 235.100 28.825 ;
        RECT 232.830 28.140 233.955 28.310 ;
        RECT 234.350 27.970 234.520 28.635 ;
        RECT 235.270 28.390 235.610 29.200 ;
        RECT 235.780 28.890 237.430 29.410 ;
        RECT 237.600 28.720 239.290 29.240 ;
        RECT 241.505 28.805 241.845 29.635 ;
        RECT 232.490 27.800 234.520 27.970 ;
        RECT 234.690 27.630 234.860 28.390 ;
        RECT 235.095 27.980 235.610 28.390 ;
        RECT 235.780 27.630 239.290 28.720 ;
        RECT 239.460 27.630 239.750 28.795 ;
        RECT 243.325 28.065 243.675 29.315 ;
        RECT 247.025 28.805 247.365 29.635 ;
        RECT 248.845 28.065 249.195 29.315 ;
        RECT 252.545 28.805 252.885 29.635 ;
        RECT 254.365 28.065 254.715 29.315 ;
        RECT 258.065 28.805 258.405 29.635 ;
        RECT 262.000 29.410 264.590 30.180 ;
        RECT 265.220 29.455 265.510 30.180 ;
        RECT 265.680 29.410 267.350 30.180 ;
        RECT 267.985 29.630 268.240 29.920 ;
        RECT 268.410 29.800 268.740 30.180 ;
        RECT 267.985 29.460 268.735 29.630 ;
        RECT 259.885 28.065 260.235 29.315 ;
        RECT 262.000 28.890 263.210 29.410 ;
        RECT 263.380 28.720 264.590 29.240 ;
        RECT 265.680 28.890 266.430 29.410 ;
        RECT 239.920 27.630 245.265 28.065 ;
        RECT 245.440 27.630 250.785 28.065 ;
        RECT 250.960 27.630 256.305 28.065 ;
        RECT 256.480 27.630 261.825 28.065 ;
        RECT 262.000 27.630 264.590 28.720 ;
        RECT 265.220 27.630 265.510 28.795 ;
        RECT 266.600 28.720 267.350 29.240 ;
        RECT 265.680 27.630 267.350 28.720 ;
        RECT 267.985 28.640 268.335 29.290 ;
        RECT 268.505 28.470 268.735 29.460 ;
        RECT 267.985 28.300 268.735 28.470 ;
        RECT 267.985 27.800 268.240 28.300 ;
        RECT 268.410 27.630 268.740 28.130 ;
        RECT 268.910 27.800 269.080 29.920 ;
        RECT 269.440 29.820 269.770 30.180 ;
        RECT 269.940 29.790 270.435 29.960 ;
        RECT 270.640 29.790 271.495 29.960 ;
        RECT 269.310 28.600 269.770 29.650 ;
        RECT 269.250 27.815 269.575 28.600 ;
        RECT 269.940 28.430 270.110 29.790 ;
        RECT 270.280 28.880 270.630 29.500 ;
        RECT 270.800 29.280 271.155 29.500 ;
        RECT 270.800 28.690 270.970 29.280 ;
        RECT 271.325 29.080 271.495 29.790 ;
        RECT 272.370 29.720 272.700 30.180 ;
        RECT 272.910 29.820 273.260 29.990 ;
        RECT 271.700 29.250 272.490 29.500 ;
        RECT 272.910 29.430 273.170 29.820 ;
        RECT 273.480 29.730 274.430 30.010 ;
        RECT 274.600 29.740 274.790 30.180 ;
        RECT 274.960 29.800 276.030 29.970 ;
        RECT 272.660 29.080 272.830 29.260 ;
        RECT 269.940 28.260 270.335 28.430 ;
        RECT 270.505 28.300 270.970 28.690 ;
        RECT 271.140 28.910 272.830 29.080 ;
        RECT 270.165 28.130 270.335 28.260 ;
        RECT 271.140 28.130 271.310 28.910 ;
        RECT 273.000 28.740 273.170 29.430 ;
        RECT 271.670 28.570 273.170 28.740 ;
        RECT 273.360 28.770 273.570 29.560 ;
        RECT 273.740 28.940 274.090 29.560 ;
        RECT 274.260 28.950 274.430 29.730 ;
        RECT 274.960 29.570 275.130 29.800 ;
        RECT 274.600 29.400 275.130 29.570 ;
        RECT 274.600 29.120 274.820 29.400 ;
        RECT 275.300 29.230 275.540 29.630 ;
        RECT 274.260 28.780 274.665 28.950 ;
        RECT 275.000 28.860 275.540 29.230 ;
        RECT 275.710 29.445 276.030 29.800 ;
        RECT 276.275 29.720 276.580 30.180 ;
        RECT 276.750 29.470 277.005 30.000 ;
        RECT 275.710 29.270 276.035 29.445 ;
        RECT 275.710 28.970 276.625 29.270 ;
        RECT 275.885 28.940 276.625 28.970 ;
        RECT 273.360 28.610 274.035 28.770 ;
        RECT 274.495 28.690 274.665 28.780 ;
        RECT 273.360 28.600 274.325 28.610 ;
        RECT 273.000 28.430 273.170 28.570 ;
        RECT 269.745 27.630 269.995 28.090 ;
        RECT 270.165 27.800 270.415 28.130 ;
        RECT 270.630 27.800 271.310 28.130 ;
        RECT 271.480 28.230 272.555 28.400 ;
        RECT 273.000 28.260 273.560 28.430 ;
        RECT 273.865 28.310 274.325 28.600 ;
        RECT 274.495 28.520 275.715 28.690 ;
        RECT 271.480 27.890 271.650 28.230 ;
        RECT 271.885 27.630 272.215 28.060 ;
        RECT 272.385 27.890 272.555 28.230 ;
        RECT 272.850 27.630 273.220 28.090 ;
        RECT 273.390 27.800 273.560 28.260 ;
        RECT 274.495 28.140 274.665 28.520 ;
        RECT 275.885 28.350 276.055 28.940 ;
        RECT 276.795 28.820 277.005 29.470 ;
        RECT 273.795 27.800 274.665 28.140 ;
        RECT 275.255 28.180 276.055 28.350 ;
        RECT 274.835 27.630 275.085 28.090 ;
        RECT 275.255 27.890 275.425 28.180 ;
        RECT 275.605 27.630 275.935 28.010 ;
        RECT 276.275 27.630 276.580 28.770 ;
        RECT 276.750 27.940 277.005 28.820 ;
        RECT 277.185 29.705 277.520 29.965 ;
        RECT 277.690 29.780 278.020 30.180 ;
        RECT 278.190 29.780 279.805 29.950 ;
        RECT 277.185 28.350 277.440 29.705 ;
        RECT 278.190 29.610 278.360 29.780 ;
        RECT 277.800 29.440 278.360 29.610 ;
        RECT 277.800 29.270 277.970 29.440 ;
        RECT 277.665 28.940 277.970 29.270 ;
        RECT 278.165 29.160 278.415 29.270 ;
        RECT 278.625 29.160 278.895 29.600 ;
        RECT 279.085 29.160 279.375 29.600 ;
        RECT 278.160 28.990 278.415 29.160 ;
        RECT 278.620 28.990 278.895 29.160 ;
        RECT 279.080 28.990 279.375 29.160 ;
        RECT 278.165 28.940 278.415 28.990 ;
        RECT 278.625 28.940 278.895 28.990 ;
        RECT 279.085 28.940 279.375 28.990 ;
        RECT 279.545 28.940 279.965 29.605 ;
        RECT 280.350 29.460 280.680 30.180 ;
        RECT 280.865 29.705 281.200 29.965 ;
        RECT 281.370 29.780 281.700 30.180 ;
        RECT 281.870 29.780 283.485 29.950 ;
        RECT 280.275 29.160 280.625 29.270 ;
        RECT 280.275 28.990 280.630 29.160 ;
        RECT 280.275 28.940 280.625 28.990 ;
        RECT 277.800 28.770 277.970 28.940 ;
        RECT 277.800 28.600 280.170 28.770 ;
        RECT 280.420 28.650 280.625 28.940 ;
        RECT 277.185 27.840 277.520 28.350 ;
        RECT 277.770 27.630 278.100 28.430 ;
        RECT 278.345 28.220 279.770 28.390 ;
        RECT 278.345 27.800 278.630 28.220 ;
        RECT 278.885 27.630 279.215 28.050 ;
        RECT 279.440 27.970 279.770 28.220 ;
        RECT 280.000 28.140 280.170 28.600 ;
        RECT 280.430 27.970 280.600 28.470 ;
        RECT 279.440 27.800 280.600 27.970 ;
        RECT 280.865 28.350 281.120 29.705 ;
        RECT 281.870 29.610 282.040 29.780 ;
        RECT 281.480 29.440 282.040 29.610 ;
        RECT 281.480 29.270 281.650 29.440 ;
        RECT 281.345 28.940 281.650 29.270 ;
        RECT 281.845 29.160 282.095 29.270 ;
        RECT 282.305 29.160 282.575 29.600 ;
        RECT 282.765 29.160 283.055 29.600 ;
        RECT 281.840 28.990 282.095 29.160 ;
        RECT 282.300 28.990 282.575 29.160 ;
        RECT 282.760 28.990 283.055 29.160 ;
        RECT 281.845 28.940 282.095 28.990 ;
        RECT 282.305 28.940 282.575 28.990 ;
        RECT 282.765 28.940 283.055 28.990 ;
        RECT 283.225 28.940 283.645 29.605 ;
        RECT 284.030 29.460 284.360 30.180 ;
        RECT 284.540 29.635 289.885 30.180 ;
        RECT 283.955 29.160 284.305 29.270 ;
        RECT 283.955 28.990 284.310 29.160 ;
        RECT 283.955 28.940 284.305 28.990 ;
        RECT 281.480 28.770 281.650 28.940 ;
        RECT 281.480 28.600 283.850 28.770 ;
        RECT 284.100 28.650 284.305 28.940 ;
        RECT 286.125 28.805 286.465 29.635 ;
        RECT 290.980 29.455 291.270 30.180 ;
        RECT 291.440 29.410 294.030 30.180 ;
        RECT 280.865 27.840 281.200 28.350 ;
        RECT 281.450 27.630 281.780 28.430 ;
        RECT 282.025 28.220 283.450 28.390 ;
        RECT 282.025 27.800 282.310 28.220 ;
        RECT 282.565 27.630 282.895 28.050 ;
        RECT 283.120 27.970 283.450 28.220 ;
        RECT 283.680 28.140 283.850 28.600 ;
        RECT 284.110 27.970 284.280 28.470 ;
        RECT 287.945 28.065 288.295 29.315 ;
        RECT 291.440 28.890 292.650 29.410 ;
        RECT 294.720 29.360 294.930 30.180 ;
        RECT 295.100 29.380 295.430 30.010 ;
        RECT 283.120 27.800 284.280 27.970 ;
        RECT 284.540 27.630 289.885 28.065 ;
        RECT 290.980 27.630 291.270 28.795 ;
        RECT 292.820 28.720 294.030 29.240 ;
        RECT 295.100 28.780 295.350 29.380 ;
        RECT 295.600 29.360 295.830 30.180 ;
        RECT 296.040 29.410 299.550 30.180 ;
        RECT 299.725 29.470 299.980 30.000 ;
        RECT 300.150 29.720 300.455 30.180 ;
        RECT 300.700 29.800 301.770 29.970 ;
        RECT 295.520 28.940 295.850 29.190 ;
        RECT 296.040 28.890 297.690 29.410 ;
        RECT 291.440 27.630 294.030 28.720 ;
        RECT 294.720 27.630 294.930 28.770 ;
        RECT 295.100 27.800 295.430 28.780 ;
        RECT 295.600 27.630 295.830 28.770 ;
        RECT 297.860 28.720 299.550 29.240 ;
        RECT 296.040 27.630 299.550 28.720 ;
        RECT 299.725 28.820 299.935 29.470 ;
        RECT 300.700 29.445 301.020 29.800 ;
        RECT 300.695 29.270 301.020 29.445 ;
        RECT 300.105 28.970 301.020 29.270 ;
        RECT 301.190 29.230 301.430 29.630 ;
        RECT 301.600 29.570 301.770 29.800 ;
        RECT 301.940 29.740 302.130 30.180 ;
        RECT 302.300 29.730 303.250 30.010 ;
        RECT 303.470 29.820 303.820 29.990 ;
        RECT 301.600 29.400 302.130 29.570 ;
        RECT 300.105 28.940 300.845 28.970 ;
        RECT 299.725 27.940 299.980 28.820 ;
        RECT 300.150 27.630 300.455 28.770 ;
        RECT 300.675 28.350 300.845 28.940 ;
        RECT 301.190 28.860 301.730 29.230 ;
        RECT 301.910 29.120 302.130 29.400 ;
        RECT 302.300 28.950 302.470 29.730 ;
        RECT 302.065 28.780 302.470 28.950 ;
        RECT 302.640 28.940 302.990 29.560 ;
        RECT 302.065 28.690 302.235 28.780 ;
        RECT 303.160 28.770 303.370 29.560 ;
        RECT 301.015 28.520 302.235 28.690 ;
        RECT 302.695 28.610 303.370 28.770 ;
        RECT 300.675 28.180 301.475 28.350 ;
        RECT 300.795 27.630 301.125 28.010 ;
        RECT 301.305 27.890 301.475 28.180 ;
        RECT 302.065 28.140 302.235 28.520 ;
        RECT 302.405 28.600 303.370 28.610 ;
        RECT 303.560 29.430 303.820 29.820 ;
        RECT 304.030 29.720 304.360 30.180 ;
        RECT 305.235 29.790 306.090 29.960 ;
        RECT 306.295 29.790 306.790 29.960 ;
        RECT 306.960 29.820 307.290 30.180 ;
        RECT 303.560 28.740 303.730 29.430 ;
        RECT 303.900 29.080 304.070 29.260 ;
        RECT 304.240 29.250 305.030 29.500 ;
        RECT 305.235 29.080 305.405 29.790 ;
        RECT 305.575 29.280 305.930 29.500 ;
        RECT 303.900 28.910 305.590 29.080 ;
        RECT 302.405 28.310 302.865 28.600 ;
        RECT 303.560 28.570 305.060 28.740 ;
        RECT 303.560 28.430 303.730 28.570 ;
        RECT 303.170 28.260 303.730 28.430 ;
        RECT 301.645 27.630 301.895 28.090 ;
        RECT 302.065 27.800 302.935 28.140 ;
        RECT 303.170 27.800 303.340 28.260 ;
        RECT 304.175 28.230 305.250 28.400 ;
        RECT 303.510 27.630 303.880 28.090 ;
        RECT 304.175 27.890 304.345 28.230 ;
        RECT 304.515 27.630 304.845 28.060 ;
        RECT 305.080 27.890 305.250 28.230 ;
        RECT 305.420 28.130 305.590 28.910 ;
        RECT 305.760 28.690 305.930 29.280 ;
        RECT 306.100 28.880 306.450 29.500 ;
        RECT 305.760 28.300 306.225 28.690 ;
        RECT 306.620 28.430 306.790 29.790 ;
        RECT 306.960 28.600 307.420 29.650 ;
        RECT 306.395 28.260 306.790 28.430 ;
        RECT 306.395 28.130 306.565 28.260 ;
        RECT 305.420 27.800 306.100 28.130 ;
        RECT 306.315 27.800 306.565 28.130 ;
        RECT 306.735 27.630 306.985 28.090 ;
        RECT 307.155 27.815 307.480 28.600 ;
        RECT 307.650 27.800 307.820 29.920 ;
        RECT 307.990 29.800 308.320 30.180 ;
        RECT 308.490 29.630 308.745 29.920 ;
        RECT 307.995 29.460 308.745 29.630 ;
        RECT 307.995 28.470 308.225 29.460 ;
        RECT 309.840 29.430 311.050 30.180 ;
        RECT 308.395 28.640 308.745 29.290 ;
        RECT 309.840 28.720 310.360 29.260 ;
        RECT 310.530 28.890 311.050 29.430 ;
        RECT 307.995 28.300 308.745 28.470 ;
        RECT 307.990 27.630 308.320 28.130 ;
        RECT 308.490 27.800 308.745 28.300 ;
        RECT 309.840 27.630 311.050 28.720 ;
        RECT 162.095 27.460 311.135 27.630 ;
        RECT 162.180 26.370 163.390 27.460 ;
        RECT 163.560 27.025 168.905 27.460 ;
        RECT 169.080 27.025 174.425 27.460 ;
        RECT 162.180 25.660 162.700 26.200 ;
        RECT 162.870 25.830 163.390 26.370 ;
        RECT 162.180 24.910 163.390 25.660 ;
        RECT 165.145 25.455 165.485 26.285 ;
        RECT 166.965 25.775 167.315 27.025 ;
        RECT 170.665 25.455 171.005 26.285 ;
        RECT 172.485 25.775 172.835 27.025 ;
        RECT 175.060 26.295 175.350 27.460 ;
        RECT 175.520 27.025 180.865 27.460 ;
        RECT 181.040 27.025 186.385 27.460 ;
        RECT 163.560 24.910 168.905 25.455 ;
        RECT 169.080 24.910 174.425 25.455 ;
        RECT 175.060 24.910 175.350 25.635 ;
        RECT 177.105 25.455 177.445 26.285 ;
        RECT 178.925 25.775 179.275 27.025 ;
        RECT 182.625 25.455 182.965 26.285 ;
        RECT 184.445 25.775 184.795 27.025 ;
        RECT 186.560 26.370 188.230 27.460 ;
        RECT 186.560 25.680 187.310 26.200 ;
        RECT 187.480 25.850 188.230 26.370 ;
        RECT 188.405 26.320 188.740 27.290 ;
        RECT 188.910 26.320 189.080 27.460 ;
        RECT 189.250 27.120 191.280 27.290 ;
        RECT 175.520 24.910 180.865 25.455 ;
        RECT 181.040 24.910 186.385 25.455 ;
        RECT 186.560 24.910 188.230 25.680 ;
        RECT 188.405 25.650 188.575 26.320 ;
        RECT 189.250 26.150 189.420 27.120 ;
        RECT 188.745 25.820 189.000 26.150 ;
        RECT 189.225 25.820 189.420 26.150 ;
        RECT 189.590 26.780 190.715 26.950 ;
        RECT 188.830 25.650 189.000 25.820 ;
        RECT 189.590 25.650 189.760 26.780 ;
        RECT 188.405 25.080 188.660 25.650 ;
        RECT 188.830 25.480 189.760 25.650 ;
        RECT 189.930 26.440 190.940 26.610 ;
        RECT 189.930 25.640 190.100 26.440 ;
        RECT 190.305 26.100 190.580 26.240 ;
        RECT 190.300 25.930 190.580 26.100 ;
        RECT 189.585 25.445 189.760 25.480 ;
        RECT 188.830 24.910 189.160 25.310 ;
        RECT 189.585 25.080 190.115 25.445 ;
        RECT 190.305 25.080 190.580 25.930 ;
        RECT 190.750 25.080 190.940 26.440 ;
        RECT 191.110 26.455 191.280 27.120 ;
        RECT 191.450 26.700 191.620 27.460 ;
        RECT 191.855 26.700 192.370 27.110 ;
        RECT 192.540 27.025 197.885 27.460 ;
        RECT 191.110 26.265 191.860 26.455 ;
        RECT 192.030 25.890 192.370 26.700 ;
        RECT 191.140 25.720 192.370 25.890 ;
        RECT 191.120 24.910 191.630 25.445 ;
        RECT 191.850 25.115 192.095 25.720 ;
        RECT 194.125 25.455 194.465 26.285 ;
        RECT 195.945 25.775 196.295 27.025 ;
        RECT 198.060 26.370 200.650 27.460 ;
        RECT 198.060 25.680 199.270 26.200 ;
        RECT 199.440 25.850 200.650 26.370 ;
        RECT 200.820 26.295 201.110 27.460 ;
        RECT 201.740 26.385 202.010 27.290 ;
        RECT 202.180 26.700 202.510 27.460 ;
        RECT 202.690 26.530 202.860 27.290 ;
        RECT 192.540 24.910 197.885 25.455 ;
        RECT 198.060 24.910 200.650 25.680 ;
        RECT 200.820 24.910 201.110 25.635 ;
        RECT 201.740 25.585 201.910 26.385 ;
        RECT 202.195 26.360 202.860 26.530 ;
        RECT 203.120 26.370 204.330 27.460 ;
        RECT 202.195 26.215 202.365 26.360 ;
        RECT 202.080 25.885 202.365 26.215 ;
        RECT 202.195 25.630 202.365 25.885 ;
        RECT 202.600 25.810 202.930 26.180 ;
        RECT 203.120 25.660 203.640 26.200 ;
        RECT 203.810 25.830 204.330 26.370 ;
        RECT 204.500 26.490 204.810 27.290 ;
        RECT 204.980 26.660 205.290 27.460 ;
        RECT 205.460 26.830 205.720 27.290 ;
        RECT 205.890 27.000 206.145 27.460 ;
        RECT 206.320 26.830 206.580 27.290 ;
        RECT 205.460 26.660 206.580 26.830 ;
        RECT 204.500 26.320 205.530 26.490 ;
        RECT 201.740 25.080 202.000 25.585 ;
        RECT 202.195 25.460 202.860 25.630 ;
        RECT 202.180 24.910 202.510 25.290 ;
        RECT 202.690 25.080 202.860 25.460 ;
        RECT 203.120 24.910 204.330 25.660 ;
        RECT 204.500 25.410 204.670 26.320 ;
        RECT 204.840 25.580 205.190 26.150 ;
        RECT 205.360 26.070 205.530 26.320 ;
        RECT 206.320 26.410 206.580 26.660 ;
        RECT 206.750 26.590 207.035 27.460 ;
        RECT 207.260 27.025 212.605 27.460 ;
        RECT 212.780 27.025 218.125 27.460 ;
        RECT 218.300 27.025 223.645 27.460 ;
        RECT 206.320 26.240 207.075 26.410 ;
        RECT 205.360 25.900 206.500 26.070 ;
        RECT 206.670 25.730 207.075 26.240 ;
        RECT 205.425 25.560 207.075 25.730 ;
        RECT 204.500 25.080 204.800 25.410 ;
        RECT 204.970 24.910 205.245 25.390 ;
        RECT 205.425 25.170 205.720 25.560 ;
        RECT 205.890 24.910 206.145 25.390 ;
        RECT 206.320 25.170 206.580 25.560 ;
        RECT 208.845 25.455 209.185 26.285 ;
        RECT 210.665 25.775 211.015 27.025 ;
        RECT 214.365 25.455 214.705 26.285 ;
        RECT 216.185 25.775 216.535 27.025 ;
        RECT 219.885 25.455 220.225 26.285 ;
        RECT 221.705 25.775 222.055 27.025 ;
        RECT 223.820 26.370 226.410 27.460 ;
        RECT 223.820 25.680 225.030 26.200 ;
        RECT 225.200 25.850 226.410 26.370 ;
        RECT 226.580 26.295 226.870 27.460 ;
        RECT 227.040 27.025 232.385 27.460 ;
        RECT 232.560 27.025 237.905 27.460 ;
        RECT 238.080 27.025 243.425 27.460 ;
        RECT 243.600 27.025 248.945 27.460 ;
        RECT 206.750 24.910 207.030 25.390 ;
        RECT 207.260 24.910 212.605 25.455 ;
        RECT 212.780 24.910 218.125 25.455 ;
        RECT 218.300 24.910 223.645 25.455 ;
        RECT 223.820 24.910 226.410 25.680 ;
        RECT 226.580 24.910 226.870 25.635 ;
        RECT 228.625 25.455 228.965 26.285 ;
        RECT 230.445 25.775 230.795 27.025 ;
        RECT 234.145 25.455 234.485 26.285 ;
        RECT 235.965 25.775 236.315 27.025 ;
        RECT 239.665 25.455 240.005 26.285 ;
        RECT 241.485 25.775 241.835 27.025 ;
        RECT 245.185 25.455 245.525 26.285 ;
        RECT 247.005 25.775 247.355 27.025 ;
        RECT 249.120 26.370 251.710 27.460 ;
        RECT 249.120 25.680 250.330 26.200 ;
        RECT 250.500 25.850 251.710 26.370 ;
        RECT 252.340 26.295 252.630 27.460 ;
        RECT 252.800 27.025 258.145 27.460 ;
        RECT 258.320 27.025 263.665 27.460 ;
        RECT 263.840 27.025 269.185 27.460 ;
        RECT 227.040 24.910 232.385 25.455 ;
        RECT 232.560 24.910 237.905 25.455 ;
        RECT 238.080 24.910 243.425 25.455 ;
        RECT 243.600 24.910 248.945 25.455 ;
        RECT 249.120 24.910 251.710 25.680 ;
        RECT 252.340 24.910 252.630 25.635 ;
        RECT 254.385 25.455 254.725 26.285 ;
        RECT 256.205 25.775 256.555 27.025 ;
        RECT 259.905 25.455 260.245 26.285 ;
        RECT 261.725 25.775 262.075 27.025 ;
        RECT 265.425 25.455 265.765 26.285 ;
        RECT 267.245 25.775 267.595 27.025 ;
        RECT 269.360 26.370 271.030 27.460 ;
        RECT 271.255 26.590 271.540 27.460 ;
        RECT 271.710 26.830 271.970 27.290 ;
        RECT 272.145 27.000 272.400 27.460 ;
        RECT 272.570 26.830 272.830 27.290 ;
        RECT 271.710 26.660 272.830 26.830 ;
        RECT 273.000 26.660 273.310 27.460 ;
        RECT 271.710 26.410 271.970 26.660 ;
        RECT 273.480 26.490 273.790 27.290 ;
        RECT 269.360 25.680 270.110 26.200 ;
        RECT 270.280 25.850 271.030 26.370 ;
        RECT 271.215 26.240 271.970 26.410 ;
        RECT 272.760 26.320 273.790 26.490 ;
        RECT 273.960 26.370 277.470 27.460 ;
        RECT 271.215 25.730 271.620 26.240 ;
        RECT 272.760 26.070 272.930 26.320 ;
        RECT 271.790 25.900 272.930 26.070 ;
        RECT 252.800 24.910 258.145 25.455 ;
        RECT 258.320 24.910 263.665 25.455 ;
        RECT 263.840 24.910 269.185 25.455 ;
        RECT 269.360 24.910 271.030 25.680 ;
        RECT 271.215 25.560 272.865 25.730 ;
        RECT 273.100 25.580 273.450 26.150 ;
        RECT 271.260 24.910 271.540 25.390 ;
        RECT 271.710 25.170 271.970 25.560 ;
        RECT 272.145 24.910 272.400 25.390 ;
        RECT 272.570 25.170 272.865 25.560 ;
        RECT 273.620 25.410 273.790 26.320 ;
        RECT 273.045 24.910 273.320 25.390 ;
        RECT 273.490 25.080 273.790 25.410 ;
        RECT 273.960 25.680 275.610 26.200 ;
        RECT 275.780 25.850 277.470 26.370 ;
        RECT 278.100 26.295 278.390 27.460 ;
        RECT 278.560 27.025 283.905 27.460 ;
        RECT 284.080 27.025 289.425 27.460 ;
        RECT 289.600 27.025 294.945 27.460 ;
        RECT 295.120 27.025 300.465 27.460 ;
        RECT 273.960 24.910 277.470 25.680 ;
        RECT 278.100 24.910 278.390 25.635 ;
        RECT 280.145 25.455 280.485 26.285 ;
        RECT 281.965 25.775 282.315 27.025 ;
        RECT 285.665 25.455 286.005 26.285 ;
        RECT 287.485 25.775 287.835 27.025 ;
        RECT 291.185 25.455 291.525 26.285 ;
        RECT 293.005 25.775 293.355 27.025 ;
        RECT 296.705 25.455 297.045 26.285 ;
        RECT 298.525 25.775 298.875 27.025 ;
        RECT 300.640 26.370 303.230 27.460 ;
        RECT 300.640 25.680 301.850 26.200 ;
        RECT 302.020 25.850 303.230 26.370 ;
        RECT 303.860 26.295 304.150 27.460 ;
        RECT 304.320 27.025 309.665 27.460 ;
        RECT 278.560 24.910 283.905 25.455 ;
        RECT 284.080 24.910 289.425 25.455 ;
        RECT 289.600 24.910 294.945 25.455 ;
        RECT 295.120 24.910 300.465 25.455 ;
        RECT 300.640 24.910 303.230 25.680 ;
        RECT 303.860 24.910 304.150 25.635 ;
        RECT 305.905 25.455 306.245 26.285 ;
        RECT 307.725 25.775 308.075 27.025 ;
        RECT 309.840 26.370 311.050 27.460 ;
        RECT 309.840 25.830 310.360 26.370 ;
        RECT 310.530 25.660 311.050 26.200 ;
        RECT 304.320 24.910 309.665 25.455 ;
        RECT 309.840 24.910 311.050 25.660 ;
        RECT 162.095 24.740 311.135 24.910 ;
        RECT 162.180 23.990 163.390 24.740 ;
        RECT 163.560 24.195 168.905 24.740 ;
        RECT 169.080 24.195 174.425 24.740 ;
        RECT 174.600 24.195 179.945 24.740 ;
        RECT 180.120 24.195 185.465 24.740 ;
        RECT 162.180 23.450 162.700 23.990 ;
        RECT 162.870 23.280 163.390 23.820 ;
        RECT 165.145 23.365 165.485 24.195 ;
        RECT 162.180 22.190 163.390 23.280 ;
        RECT 166.965 22.625 167.315 23.875 ;
        RECT 170.665 23.365 171.005 24.195 ;
        RECT 172.485 22.625 172.835 23.875 ;
        RECT 176.185 23.365 176.525 24.195 ;
        RECT 178.005 22.625 178.355 23.875 ;
        RECT 181.705 23.365 182.045 24.195 ;
        RECT 185.640 23.970 187.310 24.740 ;
        RECT 187.940 24.015 188.230 24.740 ;
        RECT 188.400 24.195 193.745 24.740 ;
        RECT 193.920 24.195 199.265 24.740 ;
        RECT 199.440 24.195 204.785 24.740 ;
        RECT 204.960 24.195 210.305 24.740 ;
        RECT 183.525 22.625 183.875 23.875 ;
        RECT 185.640 23.450 186.390 23.970 ;
        RECT 186.560 23.280 187.310 23.800 ;
        RECT 189.985 23.365 190.325 24.195 ;
        RECT 163.560 22.190 168.905 22.625 ;
        RECT 169.080 22.190 174.425 22.625 ;
        RECT 174.600 22.190 179.945 22.625 ;
        RECT 180.120 22.190 185.465 22.625 ;
        RECT 185.640 22.190 187.310 23.280 ;
        RECT 187.940 22.190 188.230 23.355 ;
        RECT 191.805 22.625 192.155 23.875 ;
        RECT 195.505 23.365 195.845 24.195 ;
        RECT 197.325 22.625 197.675 23.875 ;
        RECT 201.025 23.365 201.365 24.195 ;
        RECT 202.845 22.625 203.195 23.875 ;
        RECT 206.545 23.365 206.885 24.195 ;
        RECT 210.480 23.970 213.070 24.740 ;
        RECT 213.700 24.015 213.990 24.740 ;
        RECT 214.160 24.195 219.505 24.740 ;
        RECT 219.680 24.195 225.025 24.740 ;
        RECT 225.200 24.195 230.545 24.740 ;
        RECT 230.720 24.195 236.065 24.740 ;
        RECT 208.365 22.625 208.715 23.875 ;
        RECT 210.480 23.450 211.690 23.970 ;
        RECT 211.860 23.280 213.070 23.800 ;
        RECT 215.745 23.365 216.085 24.195 ;
        RECT 188.400 22.190 193.745 22.625 ;
        RECT 193.920 22.190 199.265 22.625 ;
        RECT 199.440 22.190 204.785 22.625 ;
        RECT 204.960 22.190 210.305 22.625 ;
        RECT 210.480 22.190 213.070 23.280 ;
        RECT 213.700 22.190 213.990 23.355 ;
        RECT 217.565 22.625 217.915 23.875 ;
        RECT 221.265 23.365 221.605 24.195 ;
        RECT 223.085 22.625 223.435 23.875 ;
        RECT 226.785 23.365 227.125 24.195 ;
        RECT 228.605 22.625 228.955 23.875 ;
        RECT 232.305 23.365 232.645 24.195 ;
        RECT 236.240 23.970 238.830 24.740 ;
        RECT 239.460 24.015 239.750 24.740 ;
        RECT 239.920 24.195 245.265 24.740 ;
        RECT 245.440 24.195 250.785 24.740 ;
        RECT 250.960 24.195 256.305 24.740 ;
        RECT 256.480 24.195 261.825 24.740 ;
        RECT 234.125 22.625 234.475 23.875 ;
        RECT 236.240 23.450 237.450 23.970 ;
        RECT 237.620 23.280 238.830 23.800 ;
        RECT 241.505 23.365 241.845 24.195 ;
        RECT 214.160 22.190 219.505 22.625 ;
        RECT 219.680 22.190 225.025 22.625 ;
        RECT 225.200 22.190 230.545 22.625 ;
        RECT 230.720 22.190 236.065 22.625 ;
        RECT 236.240 22.190 238.830 23.280 ;
        RECT 239.460 22.190 239.750 23.355 ;
        RECT 243.325 22.625 243.675 23.875 ;
        RECT 247.025 23.365 247.365 24.195 ;
        RECT 248.845 22.625 249.195 23.875 ;
        RECT 252.545 23.365 252.885 24.195 ;
        RECT 254.365 22.625 254.715 23.875 ;
        RECT 258.065 23.365 258.405 24.195 ;
        RECT 262.000 23.970 264.590 24.740 ;
        RECT 265.220 24.015 265.510 24.740 ;
        RECT 265.680 24.195 271.025 24.740 ;
        RECT 271.200 24.195 276.545 24.740 ;
        RECT 276.720 24.195 282.065 24.740 ;
        RECT 282.240 24.195 287.585 24.740 ;
        RECT 259.885 22.625 260.235 23.875 ;
        RECT 262.000 23.450 263.210 23.970 ;
        RECT 263.380 23.280 264.590 23.800 ;
        RECT 267.265 23.365 267.605 24.195 ;
        RECT 239.920 22.190 245.265 22.625 ;
        RECT 245.440 22.190 250.785 22.625 ;
        RECT 250.960 22.190 256.305 22.625 ;
        RECT 256.480 22.190 261.825 22.625 ;
        RECT 262.000 22.190 264.590 23.280 ;
        RECT 265.220 22.190 265.510 23.355 ;
        RECT 269.085 22.625 269.435 23.875 ;
        RECT 272.785 23.365 273.125 24.195 ;
        RECT 274.605 22.625 274.955 23.875 ;
        RECT 278.305 23.365 278.645 24.195 ;
        RECT 280.125 22.625 280.475 23.875 ;
        RECT 283.825 23.365 284.165 24.195 ;
        RECT 287.760 23.970 290.350 24.740 ;
        RECT 290.980 24.015 291.270 24.740 ;
        RECT 291.440 24.195 296.785 24.740 ;
        RECT 296.960 24.195 302.305 24.740 ;
        RECT 302.480 24.195 307.825 24.740 ;
        RECT 285.645 22.625 285.995 23.875 ;
        RECT 287.760 23.450 288.970 23.970 ;
        RECT 289.140 23.280 290.350 23.800 ;
        RECT 293.025 23.365 293.365 24.195 ;
        RECT 265.680 22.190 271.025 22.625 ;
        RECT 271.200 22.190 276.545 22.625 ;
        RECT 276.720 22.190 282.065 22.625 ;
        RECT 282.240 22.190 287.585 22.625 ;
        RECT 287.760 22.190 290.350 23.280 ;
        RECT 290.980 22.190 291.270 23.355 ;
        RECT 294.845 22.625 295.195 23.875 ;
        RECT 298.545 23.365 298.885 24.195 ;
        RECT 300.365 22.625 300.715 23.875 ;
        RECT 304.065 23.365 304.405 24.195 ;
        RECT 308.000 23.970 309.670 24.740 ;
        RECT 309.840 23.990 311.050 24.740 ;
        RECT 305.885 22.625 306.235 23.875 ;
        RECT 308.000 23.450 308.750 23.970 ;
        RECT 308.920 23.280 309.670 23.800 ;
        RECT 291.440 22.190 296.785 22.625 ;
        RECT 296.960 22.190 302.305 22.625 ;
        RECT 302.480 22.190 307.825 22.625 ;
        RECT 308.000 22.190 309.670 23.280 ;
        RECT 309.840 23.280 310.360 23.820 ;
        RECT 310.530 23.450 311.050 23.990 ;
        RECT 309.840 22.190 311.050 23.280 ;
        RECT 162.095 22.020 311.135 22.190 ;
        RECT 162.180 20.930 163.390 22.020 ;
        RECT 163.560 21.585 168.905 22.020 ;
        RECT 169.080 21.585 174.425 22.020 ;
        RECT 162.180 20.220 162.700 20.760 ;
        RECT 162.870 20.390 163.390 20.930 ;
        RECT 162.180 19.470 163.390 20.220 ;
        RECT 165.145 20.015 165.485 20.845 ;
        RECT 166.965 20.335 167.315 21.585 ;
        RECT 170.665 20.015 171.005 20.845 ;
        RECT 172.485 20.335 172.835 21.585 ;
        RECT 175.060 20.855 175.350 22.020 ;
        RECT 175.520 21.585 180.865 22.020 ;
        RECT 181.040 21.585 186.385 22.020 ;
        RECT 186.560 21.585 191.905 22.020 ;
        RECT 192.080 21.585 197.425 22.020 ;
        RECT 163.560 19.470 168.905 20.015 ;
        RECT 169.080 19.470 174.425 20.015 ;
        RECT 175.060 19.470 175.350 20.195 ;
        RECT 177.105 20.015 177.445 20.845 ;
        RECT 178.925 20.335 179.275 21.585 ;
        RECT 182.625 20.015 182.965 20.845 ;
        RECT 184.445 20.335 184.795 21.585 ;
        RECT 188.145 20.015 188.485 20.845 ;
        RECT 189.965 20.335 190.315 21.585 ;
        RECT 193.665 20.015 194.005 20.845 ;
        RECT 195.485 20.335 195.835 21.585 ;
        RECT 197.600 20.930 200.190 22.020 ;
        RECT 197.600 20.240 198.810 20.760 ;
        RECT 198.980 20.410 200.190 20.930 ;
        RECT 200.820 20.855 201.110 22.020 ;
        RECT 201.280 21.585 206.625 22.020 ;
        RECT 206.800 21.585 212.145 22.020 ;
        RECT 212.320 21.585 217.665 22.020 ;
        RECT 217.840 21.585 223.185 22.020 ;
        RECT 175.520 19.470 180.865 20.015 ;
        RECT 181.040 19.470 186.385 20.015 ;
        RECT 186.560 19.470 191.905 20.015 ;
        RECT 192.080 19.470 197.425 20.015 ;
        RECT 197.600 19.470 200.190 20.240 ;
        RECT 200.820 19.470 201.110 20.195 ;
        RECT 202.865 20.015 203.205 20.845 ;
        RECT 204.685 20.335 205.035 21.585 ;
        RECT 208.385 20.015 208.725 20.845 ;
        RECT 210.205 20.335 210.555 21.585 ;
        RECT 213.905 20.015 214.245 20.845 ;
        RECT 215.725 20.335 216.075 21.585 ;
        RECT 219.425 20.015 219.765 20.845 ;
        RECT 221.245 20.335 221.595 21.585 ;
        RECT 223.360 20.930 225.950 22.020 ;
        RECT 223.360 20.240 224.570 20.760 ;
        RECT 224.740 20.410 225.950 20.930 ;
        RECT 226.580 20.855 226.870 22.020 ;
        RECT 227.040 21.585 232.385 22.020 ;
        RECT 232.560 21.585 237.905 22.020 ;
        RECT 238.080 21.585 243.425 22.020 ;
        RECT 243.600 21.585 248.945 22.020 ;
        RECT 201.280 19.470 206.625 20.015 ;
        RECT 206.800 19.470 212.145 20.015 ;
        RECT 212.320 19.470 217.665 20.015 ;
        RECT 217.840 19.470 223.185 20.015 ;
        RECT 223.360 19.470 225.950 20.240 ;
        RECT 226.580 19.470 226.870 20.195 ;
        RECT 228.625 20.015 228.965 20.845 ;
        RECT 230.445 20.335 230.795 21.585 ;
        RECT 234.145 20.015 234.485 20.845 ;
        RECT 235.965 20.335 236.315 21.585 ;
        RECT 239.665 20.015 240.005 20.845 ;
        RECT 241.485 20.335 241.835 21.585 ;
        RECT 245.185 20.015 245.525 20.845 ;
        RECT 247.005 20.335 247.355 21.585 ;
        RECT 249.120 20.930 251.710 22.020 ;
        RECT 249.120 20.240 250.330 20.760 ;
        RECT 250.500 20.410 251.710 20.930 ;
        RECT 252.340 20.855 252.630 22.020 ;
        RECT 252.800 21.585 258.145 22.020 ;
        RECT 258.320 21.585 263.665 22.020 ;
        RECT 263.840 21.585 269.185 22.020 ;
        RECT 269.360 21.585 274.705 22.020 ;
        RECT 227.040 19.470 232.385 20.015 ;
        RECT 232.560 19.470 237.905 20.015 ;
        RECT 238.080 19.470 243.425 20.015 ;
        RECT 243.600 19.470 248.945 20.015 ;
        RECT 249.120 19.470 251.710 20.240 ;
        RECT 252.340 19.470 252.630 20.195 ;
        RECT 254.385 20.015 254.725 20.845 ;
        RECT 256.205 20.335 256.555 21.585 ;
        RECT 259.905 20.015 260.245 20.845 ;
        RECT 261.725 20.335 262.075 21.585 ;
        RECT 265.425 20.015 265.765 20.845 ;
        RECT 267.245 20.335 267.595 21.585 ;
        RECT 270.945 20.015 271.285 20.845 ;
        RECT 272.765 20.335 273.115 21.585 ;
        RECT 274.880 20.930 277.470 22.020 ;
        RECT 274.880 20.240 276.090 20.760 ;
        RECT 276.260 20.410 277.470 20.930 ;
        RECT 278.100 20.855 278.390 22.020 ;
        RECT 278.560 21.585 283.905 22.020 ;
        RECT 284.080 21.585 289.425 22.020 ;
        RECT 289.600 21.585 294.945 22.020 ;
        RECT 295.120 21.585 300.465 22.020 ;
        RECT 252.800 19.470 258.145 20.015 ;
        RECT 258.320 19.470 263.665 20.015 ;
        RECT 263.840 19.470 269.185 20.015 ;
        RECT 269.360 19.470 274.705 20.015 ;
        RECT 274.880 19.470 277.470 20.240 ;
        RECT 278.100 19.470 278.390 20.195 ;
        RECT 280.145 20.015 280.485 20.845 ;
        RECT 281.965 20.335 282.315 21.585 ;
        RECT 285.665 20.015 286.005 20.845 ;
        RECT 287.485 20.335 287.835 21.585 ;
        RECT 291.185 20.015 291.525 20.845 ;
        RECT 293.005 20.335 293.355 21.585 ;
        RECT 296.705 20.015 297.045 20.845 ;
        RECT 298.525 20.335 298.875 21.585 ;
        RECT 300.640 20.930 303.230 22.020 ;
        RECT 300.640 20.240 301.850 20.760 ;
        RECT 302.020 20.410 303.230 20.930 ;
        RECT 303.860 20.855 304.150 22.020 ;
        RECT 304.320 21.585 309.665 22.020 ;
        RECT 278.560 19.470 283.905 20.015 ;
        RECT 284.080 19.470 289.425 20.015 ;
        RECT 289.600 19.470 294.945 20.015 ;
        RECT 295.120 19.470 300.465 20.015 ;
        RECT 300.640 19.470 303.230 20.240 ;
        RECT 303.860 19.470 304.150 20.195 ;
        RECT 305.905 20.015 306.245 20.845 ;
        RECT 307.725 20.335 308.075 21.585 ;
        RECT 309.840 20.930 311.050 22.020 ;
        RECT 309.840 20.390 310.360 20.930 ;
        RECT 310.530 20.220 311.050 20.760 ;
        RECT 304.320 19.470 309.665 20.015 ;
        RECT 309.840 19.470 311.050 20.220 ;
        RECT 162.095 19.300 311.135 19.470 ;
        RECT 162.180 18.550 163.390 19.300 ;
        RECT 163.560 18.755 168.905 19.300 ;
        RECT 169.080 18.755 174.425 19.300 ;
        RECT 174.600 18.755 179.945 19.300 ;
        RECT 180.120 18.755 185.465 19.300 ;
        RECT 162.180 18.010 162.700 18.550 ;
        RECT 162.870 17.840 163.390 18.380 ;
        RECT 165.145 17.925 165.485 18.755 ;
        RECT 162.180 16.750 163.390 17.840 ;
        RECT 166.965 17.185 167.315 18.435 ;
        RECT 170.665 17.925 171.005 18.755 ;
        RECT 172.485 17.185 172.835 18.435 ;
        RECT 176.185 17.925 176.525 18.755 ;
        RECT 178.005 17.185 178.355 18.435 ;
        RECT 181.705 17.925 182.045 18.755 ;
        RECT 185.640 18.530 187.310 19.300 ;
        RECT 187.940 18.575 188.230 19.300 ;
        RECT 188.400 18.755 193.745 19.300 ;
        RECT 193.920 18.755 199.265 19.300 ;
        RECT 199.440 18.755 204.785 19.300 ;
        RECT 204.960 18.755 210.305 19.300 ;
        RECT 183.525 17.185 183.875 18.435 ;
        RECT 185.640 18.010 186.390 18.530 ;
        RECT 186.560 17.840 187.310 18.360 ;
        RECT 189.985 17.925 190.325 18.755 ;
        RECT 163.560 16.750 168.905 17.185 ;
        RECT 169.080 16.750 174.425 17.185 ;
        RECT 174.600 16.750 179.945 17.185 ;
        RECT 180.120 16.750 185.465 17.185 ;
        RECT 185.640 16.750 187.310 17.840 ;
        RECT 187.940 16.750 188.230 17.915 ;
        RECT 191.805 17.185 192.155 18.435 ;
        RECT 195.505 17.925 195.845 18.755 ;
        RECT 197.325 17.185 197.675 18.435 ;
        RECT 201.025 17.925 201.365 18.755 ;
        RECT 202.845 17.185 203.195 18.435 ;
        RECT 206.545 17.925 206.885 18.755 ;
        RECT 210.480 18.530 213.070 19.300 ;
        RECT 213.700 18.575 213.990 19.300 ;
        RECT 214.160 18.755 219.505 19.300 ;
        RECT 219.680 18.755 225.025 19.300 ;
        RECT 225.200 18.755 230.545 19.300 ;
        RECT 230.720 18.755 236.065 19.300 ;
        RECT 208.365 17.185 208.715 18.435 ;
        RECT 210.480 18.010 211.690 18.530 ;
        RECT 211.860 17.840 213.070 18.360 ;
        RECT 215.745 17.925 216.085 18.755 ;
        RECT 188.400 16.750 193.745 17.185 ;
        RECT 193.920 16.750 199.265 17.185 ;
        RECT 199.440 16.750 204.785 17.185 ;
        RECT 204.960 16.750 210.305 17.185 ;
        RECT 210.480 16.750 213.070 17.840 ;
        RECT 213.700 16.750 213.990 17.915 ;
        RECT 217.565 17.185 217.915 18.435 ;
        RECT 221.265 17.925 221.605 18.755 ;
        RECT 223.085 17.185 223.435 18.435 ;
        RECT 226.785 17.925 227.125 18.755 ;
        RECT 228.605 17.185 228.955 18.435 ;
        RECT 232.305 17.925 232.645 18.755 ;
        RECT 236.240 18.530 238.830 19.300 ;
        RECT 239.460 18.575 239.750 19.300 ;
        RECT 239.920 18.755 245.265 19.300 ;
        RECT 245.440 18.755 250.785 19.300 ;
        RECT 250.960 18.755 256.305 19.300 ;
        RECT 256.480 18.755 261.825 19.300 ;
        RECT 234.125 17.185 234.475 18.435 ;
        RECT 236.240 18.010 237.450 18.530 ;
        RECT 237.620 17.840 238.830 18.360 ;
        RECT 241.505 17.925 241.845 18.755 ;
        RECT 214.160 16.750 219.505 17.185 ;
        RECT 219.680 16.750 225.025 17.185 ;
        RECT 225.200 16.750 230.545 17.185 ;
        RECT 230.720 16.750 236.065 17.185 ;
        RECT 236.240 16.750 238.830 17.840 ;
        RECT 239.460 16.750 239.750 17.915 ;
        RECT 243.325 17.185 243.675 18.435 ;
        RECT 247.025 17.925 247.365 18.755 ;
        RECT 248.845 17.185 249.195 18.435 ;
        RECT 252.545 17.925 252.885 18.755 ;
        RECT 254.365 17.185 254.715 18.435 ;
        RECT 258.065 17.925 258.405 18.755 ;
        RECT 262.000 18.530 264.590 19.300 ;
        RECT 265.220 18.575 265.510 19.300 ;
        RECT 265.680 18.755 271.025 19.300 ;
        RECT 271.200 18.755 276.545 19.300 ;
        RECT 276.720 18.755 282.065 19.300 ;
        RECT 282.240 18.755 287.585 19.300 ;
        RECT 259.885 17.185 260.235 18.435 ;
        RECT 262.000 18.010 263.210 18.530 ;
        RECT 263.380 17.840 264.590 18.360 ;
        RECT 267.265 17.925 267.605 18.755 ;
        RECT 239.920 16.750 245.265 17.185 ;
        RECT 245.440 16.750 250.785 17.185 ;
        RECT 250.960 16.750 256.305 17.185 ;
        RECT 256.480 16.750 261.825 17.185 ;
        RECT 262.000 16.750 264.590 17.840 ;
        RECT 265.220 16.750 265.510 17.915 ;
        RECT 269.085 17.185 269.435 18.435 ;
        RECT 272.785 17.925 273.125 18.755 ;
        RECT 274.605 17.185 274.955 18.435 ;
        RECT 278.305 17.925 278.645 18.755 ;
        RECT 280.125 17.185 280.475 18.435 ;
        RECT 283.825 17.925 284.165 18.755 ;
        RECT 287.760 18.530 290.350 19.300 ;
        RECT 290.980 18.575 291.270 19.300 ;
        RECT 291.440 18.755 296.785 19.300 ;
        RECT 296.960 18.755 302.305 19.300 ;
        RECT 302.480 18.755 307.825 19.300 ;
        RECT 285.645 17.185 285.995 18.435 ;
        RECT 287.760 18.010 288.970 18.530 ;
        RECT 289.140 17.840 290.350 18.360 ;
        RECT 293.025 17.925 293.365 18.755 ;
        RECT 265.680 16.750 271.025 17.185 ;
        RECT 271.200 16.750 276.545 17.185 ;
        RECT 276.720 16.750 282.065 17.185 ;
        RECT 282.240 16.750 287.585 17.185 ;
        RECT 287.760 16.750 290.350 17.840 ;
        RECT 290.980 16.750 291.270 17.915 ;
        RECT 294.845 17.185 295.195 18.435 ;
        RECT 298.545 17.925 298.885 18.755 ;
        RECT 300.365 17.185 300.715 18.435 ;
        RECT 304.065 17.925 304.405 18.755 ;
        RECT 308.000 18.530 309.670 19.300 ;
        RECT 309.840 18.550 311.050 19.300 ;
        RECT 305.885 17.185 306.235 18.435 ;
        RECT 308.000 18.010 308.750 18.530 ;
        RECT 308.920 17.840 309.670 18.360 ;
        RECT 291.440 16.750 296.785 17.185 ;
        RECT 296.960 16.750 302.305 17.185 ;
        RECT 302.480 16.750 307.825 17.185 ;
        RECT 308.000 16.750 309.670 17.840 ;
        RECT 309.840 17.840 310.360 18.380 ;
        RECT 310.530 18.010 311.050 18.550 ;
        RECT 309.840 16.750 311.050 17.840 ;
        RECT 162.095 16.580 311.135 16.750 ;
        RECT 162.180 15.490 163.390 16.580 ;
        RECT 163.560 16.145 168.905 16.580 ;
        RECT 169.080 16.145 174.425 16.580 ;
        RECT 162.180 14.780 162.700 15.320 ;
        RECT 162.870 14.950 163.390 15.490 ;
        RECT 162.180 14.030 163.390 14.780 ;
        RECT 165.145 14.575 165.485 15.405 ;
        RECT 166.965 14.895 167.315 16.145 ;
        RECT 170.665 14.575 171.005 15.405 ;
        RECT 172.485 14.895 172.835 16.145 ;
        RECT 175.060 15.415 175.350 16.580 ;
        RECT 175.520 16.145 180.865 16.580 ;
        RECT 181.040 16.145 186.385 16.580 ;
        RECT 163.560 14.030 168.905 14.575 ;
        RECT 169.080 14.030 174.425 14.575 ;
        RECT 175.060 14.030 175.350 14.755 ;
        RECT 177.105 14.575 177.445 15.405 ;
        RECT 178.925 14.895 179.275 16.145 ;
        RECT 182.625 14.575 182.965 15.405 ;
        RECT 184.445 14.895 184.795 16.145 ;
        RECT 186.560 15.490 187.770 16.580 ;
        RECT 186.560 14.780 187.080 15.320 ;
        RECT 187.250 14.950 187.770 15.490 ;
        RECT 187.940 15.415 188.230 16.580 ;
        RECT 188.400 16.145 193.745 16.580 ;
        RECT 193.920 16.145 199.265 16.580 ;
        RECT 175.520 14.030 180.865 14.575 ;
        RECT 181.040 14.030 186.385 14.575 ;
        RECT 186.560 14.030 187.770 14.780 ;
        RECT 187.940 14.030 188.230 14.755 ;
        RECT 189.985 14.575 190.325 15.405 ;
        RECT 191.805 14.895 192.155 16.145 ;
        RECT 195.505 14.575 195.845 15.405 ;
        RECT 197.325 14.895 197.675 16.145 ;
        RECT 199.440 15.490 200.650 16.580 ;
        RECT 199.440 14.780 199.960 15.320 ;
        RECT 200.130 14.950 200.650 15.490 ;
        RECT 200.820 15.415 201.110 16.580 ;
        RECT 201.280 16.145 206.625 16.580 ;
        RECT 206.800 16.145 212.145 16.580 ;
        RECT 188.400 14.030 193.745 14.575 ;
        RECT 193.920 14.030 199.265 14.575 ;
        RECT 199.440 14.030 200.650 14.780 ;
        RECT 200.820 14.030 201.110 14.755 ;
        RECT 202.865 14.575 203.205 15.405 ;
        RECT 204.685 14.895 205.035 16.145 ;
        RECT 208.385 14.575 208.725 15.405 ;
        RECT 210.205 14.895 210.555 16.145 ;
        RECT 212.320 15.490 213.530 16.580 ;
        RECT 212.320 14.780 212.840 15.320 ;
        RECT 213.010 14.950 213.530 15.490 ;
        RECT 213.700 15.415 213.990 16.580 ;
        RECT 214.160 16.145 219.505 16.580 ;
        RECT 219.680 16.145 225.025 16.580 ;
        RECT 201.280 14.030 206.625 14.575 ;
        RECT 206.800 14.030 212.145 14.575 ;
        RECT 212.320 14.030 213.530 14.780 ;
        RECT 213.700 14.030 213.990 14.755 ;
        RECT 215.745 14.575 216.085 15.405 ;
        RECT 217.565 14.895 217.915 16.145 ;
        RECT 221.265 14.575 221.605 15.405 ;
        RECT 223.085 14.895 223.435 16.145 ;
        RECT 225.200 15.490 226.410 16.580 ;
        RECT 225.200 14.780 225.720 15.320 ;
        RECT 225.890 14.950 226.410 15.490 ;
        RECT 226.580 15.415 226.870 16.580 ;
        RECT 227.040 16.145 232.385 16.580 ;
        RECT 232.560 16.145 237.905 16.580 ;
        RECT 214.160 14.030 219.505 14.575 ;
        RECT 219.680 14.030 225.025 14.575 ;
        RECT 225.200 14.030 226.410 14.780 ;
        RECT 226.580 14.030 226.870 14.755 ;
        RECT 228.625 14.575 228.965 15.405 ;
        RECT 230.445 14.895 230.795 16.145 ;
        RECT 234.145 14.575 234.485 15.405 ;
        RECT 235.965 14.895 236.315 16.145 ;
        RECT 238.080 15.490 239.290 16.580 ;
        RECT 238.080 14.780 238.600 15.320 ;
        RECT 238.770 14.950 239.290 15.490 ;
        RECT 239.460 15.415 239.750 16.580 ;
        RECT 239.920 16.145 245.265 16.580 ;
        RECT 245.440 16.145 250.785 16.580 ;
        RECT 227.040 14.030 232.385 14.575 ;
        RECT 232.560 14.030 237.905 14.575 ;
        RECT 238.080 14.030 239.290 14.780 ;
        RECT 239.460 14.030 239.750 14.755 ;
        RECT 241.505 14.575 241.845 15.405 ;
        RECT 243.325 14.895 243.675 16.145 ;
        RECT 247.025 14.575 247.365 15.405 ;
        RECT 248.845 14.895 249.195 16.145 ;
        RECT 250.960 15.490 252.170 16.580 ;
        RECT 250.960 14.780 251.480 15.320 ;
        RECT 251.650 14.950 252.170 15.490 ;
        RECT 252.340 15.415 252.630 16.580 ;
        RECT 252.800 16.145 258.145 16.580 ;
        RECT 258.320 16.145 263.665 16.580 ;
        RECT 239.920 14.030 245.265 14.575 ;
        RECT 245.440 14.030 250.785 14.575 ;
        RECT 250.960 14.030 252.170 14.780 ;
        RECT 252.340 14.030 252.630 14.755 ;
        RECT 254.385 14.575 254.725 15.405 ;
        RECT 256.205 14.895 256.555 16.145 ;
        RECT 259.905 14.575 260.245 15.405 ;
        RECT 261.725 14.895 262.075 16.145 ;
        RECT 263.840 15.490 265.050 16.580 ;
        RECT 263.840 14.780 264.360 15.320 ;
        RECT 264.530 14.950 265.050 15.490 ;
        RECT 265.220 15.415 265.510 16.580 ;
        RECT 265.680 16.145 271.025 16.580 ;
        RECT 271.200 16.145 276.545 16.580 ;
        RECT 252.800 14.030 258.145 14.575 ;
        RECT 258.320 14.030 263.665 14.575 ;
        RECT 263.840 14.030 265.050 14.780 ;
        RECT 265.220 14.030 265.510 14.755 ;
        RECT 267.265 14.575 267.605 15.405 ;
        RECT 269.085 14.895 269.435 16.145 ;
        RECT 272.785 14.575 273.125 15.405 ;
        RECT 274.605 14.895 274.955 16.145 ;
        RECT 276.720 15.490 277.930 16.580 ;
        RECT 276.720 14.780 277.240 15.320 ;
        RECT 277.410 14.950 277.930 15.490 ;
        RECT 278.100 15.415 278.390 16.580 ;
        RECT 278.560 16.145 283.905 16.580 ;
        RECT 284.080 16.145 289.425 16.580 ;
        RECT 265.680 14.030 271.025 14.575 ;
        RECT 271.200 14.030 276.545 14.575 ;
        RECT 276.720 14.030 277.930 14.780 ;
        RECT 278.100 14.030 278.390 14.755 ;
        RECT 280.145 14.575 280.485 15.405 ;
        RECT 281.965 14.895 282.315 16.145 ;
        RECT 285.665 14.575 286.005 15.405 ;
        RECT 287.485 14.895 287.835 16.145 ;
        RECT 289.600 15.490 290.810 16.580 ;
        RECT 289.600 14.780 290.120 15.320 ;
        RECT 290.290 14.950 290.810 15.490 ;
        RECT 290.980 15.415 291.270 16.580 ;
        RECT 291.440 16.145 296.785 16.580 ;
        RECT 296.960 16.145 302.305 16.580 ;
        RECT 278.560 14.030 283.905 14.575 ;
        RECT 284.080 14.030 289.425 14.575 ;
        RECT 289.600 14.030 290.810 14.780 ;
        RECT 290.980 14.030 291.270 14.755 ;
        RECT 293.025 14.575 293.365 15.405 ;
        RECT 294.845 14.895 295.195 16.145 ;
        RECT 298.545 14.575 298.885 15.405 ;
        RECT 300.365 14.895 300.715 16.145 ;
        RECT 302.480 15.490 303.690 16.580 ;
        RECT 302.480 14.780 303.000 15.320 ;
        RECT 303.170 14.950 303.690 15.490 ;
        RECT 303.860 15.415 304.150 16.580 ;
        RECT 304.320 16.145 309.665 16.580 ;
        RECT 291.440 14.030 296.785 14.575 ;
        RECT 296.960 14.030 302.305 14.575 ;
        RECT 302.480 14.030 303.690 14.780 ;
        RECT 303.860 14.030 304.150 14.755 ;
        RECT 305.905 14.575 306.245 15.405 ;
        RECT 307.725 14.895 308.075 16.145 ;
        RECT 309.840 15.490 311.050 16.580 ;
        RECT 309.840 14.950 310.360 15.490 ;
        RECT 310.530 14.780 311.050 15.320 ;
        RECT 304.320 14.030 309.665 14.575 ;
        RECT 309.840 14.030 311.050 14.780 ;
        RECT 162.095 13.860 311.135 14.030 ;
        RECT 4.300 4.300 155.700 4.700 ;
      LAYER met1 ;
        RECT 45.390 225.410 246.965 225.710 ;
        RECT 45.390 224.810 45.690 225.410 ;
        RECT 59.190 224.810 236.370 225.110 ;
        RECT 246.665 225.010 246.965 225.410 ;
        RECT 62.000 224.210 226.710 224.510 ;
        RECT 236.070 224.410 236.370 224.810 ;
        RECT 226.410 223.810 226.710 224.210 ;
        RECT 4.100 216.515 102.825 222.630 ;
        RECT 106.340 220.315 153.245 220.715 ;
        RECT 106.340 217.515 108.920 220.315 ;
        RECT 109.605 219.705 110.565 219.935 ;
        RECT 110.895 219.705 111.855 220.055 ;
        RECT 109.325 219.255 109.555 219.500 ;
        RECT 110.615 219.255 110.845 219.500 ;
        RECT 111.905 219.255 112.135 219.500 ;
        RECT 109.290 217.755 109.590 219.255 ;
        RECT 110.580 217.755 110.880 219.255 ;
        RECT 111.870 217.755 112.170 219.255 ;
        RECT 4.100 212.490 63.455 216.515 ;
        RECT 64.175 215.825 80.135 216.055 ;
        RECT 81.805 215.825 97.765 216.055 ;
        RECT 63.895 214.620 64.125 215.620 ;
        RECT 80.185 214.620 81.755 215.620 ;
        RECT 97.815 214.620 98.045 215.620 ;
        RECT 64.175 214.185 80.135 214.415 ;
        RECT 81.805 214.185 97.765 214.415 ;
        RECT 77.595 213.035 78.595 213.270 ;
        RECT 83.345 213.035 84.345 213.270 ;
        RECT 64.175 212.805 80.135 213.035 ;
        RECT 81.805 212.805 97.765 213.035 ;
        RECT 4.100 211.660 56.570 212.490 ;
        RECT 4.100 191.850 9.525 211.660 ;
        RECT 10.245 210.970 18.205 211.200 ;
        RECT 18.535 210.970 26.495 211.200 ;
        RECT 28.165 210.970 36.125 211.200 ;
        RECT 36.455 210.970 44.415 211.200 ;
        RECT 9.965 210.465 10.195 210.765 ;
        RECT 9.925 209.065 10.225 210.465 ;
        RECT 9.965 202.765 10.195 209.065 ;
        RECT 18.255 207.465 18.485 210.765 ;
        RECT 18.215 206.065 18.515 207.465 ;
        RECT 18.255 202.765 18.485 206.065 ;
        RECT 26.545 204.465 26.775 210.765 ;
        RECT 27.885 204.465 28.115 210.765 ;
        RECT 36.175 207.465 36.405 210.765 ;
        RECT 44.465 210.465 44.695 210.765 ;
        RECT 44.425 209.065 44.725 210.465 ;
        RECT 45.135 210.150 56.570 211.660 ;
        RECT 36.165 206.065 36.465 207.465 ;
        RECT 26.505 203.065 26.805 204.465 ;
        RECT 27.845 203.065 28.145 204.465 ;
        RECT 26.505 202.560 28.145 203.065 ;
        RECT 36.175 202.765 36.405 206.065 ;
        RECT 44.465 202.765 44.695 209.065 ;
        RECT 45.135 207.460 50.745 210.150 ;
        RECT 54.835 209.565 56.570 210.150 ;
        RECT 51.315 207.460 51.905 209.565 ;
        RECT 52.485 207.460 54.245 209.565 ;
        RECT 54.825 207.460 56.570 209.565 ;
        RECT 10.245 202.330 18.205 202.560 ;
        RECT 18.535 202.330 36.125 202.560 ;
        RECT 36.455 202.330 44.415 202.560 ;
        RECT 10.245 201.180 44.415 202.330 ;
        RECT 10.245 200.950 18.205 201.180 ;
        RECT 18.535 200.950 36.125 201.180 ;
        RECT 36.455 200.950 44.415 201.180 ;
        RECT 9.965 194.445 10.195 200.745 ;
        RECT 18.255 197.445 18.485 200.745 ;
        RECT 26.505 200.445 28.145 200.950 ;
        RECT 26.505 199.045 26.805 200.445 ;
        RECT 27.845 199.045 28.145 200.445 ;
        RECT 18.215 196.045 18.515 197.445 ;
        RECT 9.925 193.045 10.225 194.445 ;
        RECT 9.965 192.745 10.195 193.045 ;
        RECT 18.255 192.745 18.485 196.045 ;
        RECT 26.545 192.745 26.775 199.045 ;
        RECT 27.885 192.745 28.115 199.045 ;
        RECT 36.175 197.445 36.405 200.745 ;
        RECT 36.165 196.045 36.465 197.445 ;
        RECT 36.175 192.745 36.405 196.045 ;
        RECT 44.465 194.445 44.695 200.745 ;
        RECT 44.425 193.045 44.725 194.445 ;
        RECT 44.465 192.745 44.695 193.045 ;
        RECT 10.245 192.310 18.205 192.540 ;
        RECT 18.535 192.310 26.495 192.540 ;
        RECT 28.165 192.310 36.125 192.540 ;
        RECT 36.455 192.310 44.415 192.540 ;
        RECT 45.135 191.850 49.450 207.460 ;
        RECT 4.100 190.670 49.450 191.850 ;
        RECT 4.100 180.880 9.525 190.670 ;
        RECT 9.965 189.980 12.205 190.210 ;
        RECT 12.535 189.980 14.495 190.210 ;
        RECT 9.965 184.050 10.195 189.980 ;
        RECT 12.535 189.775 13.090 189.980 ;
        RECT 12.255 189.350 13.090 189.775 ;
        RECT 9.930 182.650 10.230 184.050 ;
        RECT 9.965 181.570 10.195 182.650 ;
        RECT 12.255 181.775 12.485 189.350 ;
        RECT 14.545 188.900 14.775 189.775 ;
        RECT 14.510 187.500 14.810 188.900 ;
        RECT 14.545 181.775 14.775 187.500 ;
        RECT 9.965 181.340 12.205 181.570 ;
        RECT 12.535 181.340 14.495 181.570 ;
        RECT 15.215 180.880 16.545 190.670 ;
        RECT 45.135 190.570 49.450 190.670 ;
        RECT 56.110 190.570 56.570 207.460 ;
        RECT 17.265 189.980 19.225 190.210 ;
        RECT 19.555 189.980 21.515 190.210 ;
        RECT 21.845 189.980 23.805 190.210 ;
        RECT 24.135 189.980 26.095 190.210 ;
        RECT 26.425 189.980 28.385 190.210 ;
        RECT 28.715 189.980 30.675 190.210 ;
        RECT 31.005 189.980 32.965 190.210 ;
        RECT 33.295 189.980 35.255 190.210 ;
        RECT 35.585 189.980 37.545 190.210 ;
        RECT 37.875 189.980 39.835 190.210 ;
        RECT 40.165 189.980 42.125 190.210 ;
        RECT 42.455 189.980 44.415 190.210 ;
        RECT 16.985 189.645 17.215 189.775 ;
        RECT 16.950 188.245 17.250 189.645 ;
        RECT 16.985 181.775 17.215 188.245 ;
        RECT 19.275 186.555 19.505 189.775 ;
        RECT 21.565 189.645 21.795 189.775 ;
        RECT 21.530 188.245 21.830 189.645 ;
        RECT 19.240 184.995 19.540 186.555 ;
        RECT 19.275 181.775 19.505 184.995 ;
        RECT 21.565 181.775 21.795 188.245 ;
        RECT 23.855 186.555 24.085 189.775 ;
        RECT 26.145 189.645 26.375 189.775 ;
        RECT 26.110 188.245 26.410 189.645 ;
        RECT 23.820 184.995 24.120 186.555 ;
        RECT 23.855 181.775 24.085 184.995 ;
        RECT 26.145 181.775 26.375 188.245 ;
        RECT 28.435 186.555 28.665 189.775 ;
        RECT 30.725 189.645 30.955 189.775 ;
        RECT 30.690 188.245 30.990 189.645 ;
        RECT 28.400 184.995 28.700 186.555 ;
        RECT 28.435 181.775 28.665 184.995 ;
        RECT 30.725 181.775 30.955 188.245 ;
        RECT 33.015 186.555 33.245 189.775 ;
        RECT 35.305 189.645 35.535 189.775 ;
        RECT 35.270 188.245 35.570 189.645 ;
        RECT 32.980 184.995 33.280 186.555 ;
        RECT 33.015 181.775 33.245 184.995 ;
        RECT 35.305 181.775 35.535 188.245 ;
        RECT 37.595 186.555 37.825 189.775 ;
        RECT 39.885 189.645 40.115 189.775 ;
        RECT 39.850 188.245 40.150 189.645 ;
        RECT 37.560 184.995 37.860 186.555 ;
        RECT 37.595 181.775 37.825 184.995 ;
        RECT 39.885 181.775 40.115 188.245 ;
        RECT 42.175 186.555 42.405 189.775 ;
        RECT 44.465 189.645 44.695 189.775 ;
        RECT 44.430 188.245 44.730 189.645 ;
        RECT 42.140 184.995 42.440 186.555 ;
        RECT 42.175 181.775 42.405 184.995 ;
        RECT 44.465 181.775 44.695 188.245 ;
        RECT 45.135 187.880 50.745 190.570 ;
        RECT 51.315 188.465 53.075 190.570 ;
        RECT 53.655 188.465 54.245 190.570 ;
        RECT 54.825 188.465 56.570 190.570 ;
        RECT 54.835 187.880 56.570 188.465 ;
        RECT 45.135 187.650 56.570 187.880 ;
        RECT 17.465 181.570 19.025 181.605 ;
        RECT 19.755 181.570 21.315 181.605 ;
        RECT 22.045 181.570 23.605 181.605 ;
        RECT 24.335 181.570 25.895 181.605 ;
        RECT 26.625 181.570 28.185 181.605 ;
        RECT 28.915 181.570 30.475 181.605 ;
        RECT 31.205 181.570 32.765 181.605 ;
        RECT 33.495 181.570 35.055 181.605 ;
        RECT 35.785 181.570 37.345 181.605 ;
        RECT 38.075 181.570 39.635 181.605 ;
        RECT 40.365 181.570 41.925 181.605 ;
        RECT 42.655 181.570 44.215 181.605 ;
        RECT 17.265 181.340 44.415 181.570 ;
        RECT 17.465 181.305 19.025 181.340 ;
        RECT 19.755 181.305 21.315 181.340 ;
        RECT 22.045 181.305 23.605 181.340 ;
        RECT 24.335 181.305 25.895 181.340 ;
        RECT 26.625 181.305 28.185 181.340 ;
        RECT 28.915 181.305 30.475 181.340 ;
        RECT 31.205 181.305 32.765 181.340 ;
        RECT 33.495 181.305 35.055 181.340 ;
        RECT 35.785 181.305 37.345 181.340 ;
        RECT 38.075 181.305 39.635 181.340 ;
        RECT 40.365 181.305 41.925 181.340 ;
        RECT 42.655 181.305 44.215 181.340 ;
        RECT 45.135 180.880 46.085 187.650 ;
        RECT 4.100 180.050 46.085 180.880 ;
        RECT 4.100 127.485 4.900 180.050 ;
        RECT 5.910 178.420 53.180 179.250 ;
        RECT 5.910 168.720 9.530 178.420 ;
        RECT 17.400 177.960 18.800 178.130 ;
        RECT 19.690 177.960 21.090 178.130 ;
        RECT 26.560 177.960 27.960 178.130 ;
        RECT 28.850 177.960 30.250 178.130 ;
        RECT 35.720 177.960 37.120 178.130 ;
        RECT 38.010 177.960 39.410 178.130 ;
        RECT 44.880 177.960 46.280 178.130 ;
        RECT 47.170 177.960 48.570 178.130 ;
        RECT 49.460 177.960 50.860 178.130 ;
        RECT 10.250 177.730 12.210 177.960 ;
        RECT 12.540 177.730 14.500 177.960 ;
        RECT 14.830 177.730 16.790 177.960 ;
        RECT 17.120 177.730 19.080 177.960 ;
        RECT 19.410 177.730 21.370 177.960 ;
        RECT 21.700 177.730 23.660 177.960 ;
        RECT 23.990 177.730 25.950 177.960 ;
        RECT 26.280 177.730 28.240 177.960 ;
        RECT 28.570 177.730 30.530 177.960 ;
        RECT 30.860 177.730 32.820 177.960 ;
        RECT 33.150 177.730 35.110 177.960 ;
        RECT 35.440 177.730 37.400 177.960 ;
        RECT 37.730 177.730 39.690 177.960 ;
        RECT 40.020 177.730 41.980 177.960 ;
        RECT 42.310 177.730 44.270 177.960 ;
        RECT 44.600 177.730 46.560 177.960 ;
        RECT 46.890 177.730 48.850 177.960 ;
        RECT 49.180 177.730 51.140 177.960 ;
        RECT 9.970 174.270 10.200 177.570 ;
        RECT 12.260 174.270 12.490 177.570 ;
        RECT 14.550 176.670 14.780 177.570 ;
        RECT 14.465 175.270 14.865 176.670 ;
        RECT 9.885 172.870 10.285 174.270 ;
        RECT 12.175 172.870 12.575 174.270 ;
        RECT 9.970 169.570 10.200 172.870 ;
        RECT 12.260 169.570 12.490 172.870 ;
        RECT 14.550 169.570 14.780 175.270 ;
        RECT 16.840 174.270 17.070 177.570 ;
        RECT 16.755 172.870 17.155 174.270 ;
        RECT 16.840 169.570 17.070 172.870 ;
        RECT 19.130 171.870 19.360 177.570 ;
        RECT 21.420 174.270 21.650 177.570 ;
        RECT 23.710 176.670 23.940 177.570 ;
        RECT 23.625 175.270 24.025 176.670 ;
        RECT 21.335 172.870 21.735 174.270 ;
        RECT 19.045 170.470 19.445 171.870 ;
        RECT 19.130 169.570 19.360 170.470 ;
        RECT 21.420 169.570 21.650 172.870 ;
        RECT 23.710 169.570 23.940 175.270 ;
        RECT 26.000 174.270 26.230 177.570 ;
        RECT 25.915 172.870 26.315 174.270 ;
        RECT 26.000 169.570 26.230 172.870 ;
        RECT 28.290 171.870 28.520 177.570 ;
        RECT 30.580 174.270 30.810 177.570 ;
        RECT 32.870 176.670 33.100 177.570 ;
        RECT 32.785 175.270 33.185 176.670 ;
        RECT 30.495 172.870 30.895 174.270 ;
        RECT 28.205 170.470 28.605 171.870 ;
        RECT 28.290 169.570 28.520 170.470 ;
        RECT 30.580 169.570 30.810 172.870 ;
        RECT 32.870 169.570 33.100 175.270 ;
        RECT 35.160 174.270 35.390 177.570 ;
        RECT 35.075 172.870 35.475 174.270 ;
        RECT 35.160 169.570 35.390 172.870 ;
        RECT 37.450 171.870 37.680 177.570 ;
        RECT 39.740 174.270 39.970 177.570 ;
        RECT 42.030 176.670 42.260 177.570 ;
        RECT 41.945 175.270 42.345 176.670 ;
        RECT 39.655 172.870 40.055 174.270 ;
        RECT 37.365 170.470 37.765 171.870 ;
        RECT 37.450 169.570 37.680 170.470 ;
        RECT 39.740 169.570 39.970 172.870 ;
        RECT 42.030 169.570 42.260 175.270 ;
        RECT 44.320 174.270 44.550 177.570 ;
        RECT 44.235 172.870 44.635 174.270 ;
        RECT 44.320 169.570 44.550 172.870 ;
        RECT 46.610 171.870 46.840 177.570 ;
        RECT 48.900 174.270 49.130 177.570 ;
        RECT 51.190 174.270 51.420 177.570 ;
        RECT 48.815 172.870 49.215 174.270 ;
        RECT 51.105 172.870 51.505 174.270 ;
        RECT 46.525 170.470 46.925 171.870 ;
        RECT 46.610 169.570 46.840 170.470 ;
        RECT 48.900 169.570 49.130 172.870 ;
        RECT 51.190 169.570 51.420 172.870 ;
        RECT 10.250 169.180 12.210 169.410 ;
        RECT 12.540 169.180 14.500 169.410 ;
        RECT 14.830 169.180 16.790 169.410 ;
        RECT 17.120 169.180 19.080 169.410 ;
        RECT 19.410 169.180 21.370 169.410 ;
        RECT 21.700 169.180 23.660 169.410 ;
        RECT 23.990 169.180 25.950 169.410 ;
        RECT 26.280 169.180 28.240 169.410 ;
        RECT 28.570 169.180 30.530 169.410 ;
        RECT 30.860 169.180 32.820 169.410 ;
        RECT 33.150 169.180 35.110 169.410 ;
        RECT 35.440 169.180 37.400 169.410 ;
        RECT 37.730 169.180 39.690 169.410 ;
        RECT 40.020 169.180 41.980 169.410 ;
        RECT 42.310 169.180 44.270 169.410 ;
        RECT 44.600 169.180 46.560 169.410 ;
        RECT 46.890 169.180 48.850 169.410 ;
        RECT 49.180 169.180 51.140 169.410 ;
        RECT 10.530 169.010 11.930 169.180 ;
        RECT 12.820 169.010 14.220 169.180 ;
        RECT 15.110 169.010 16.510 169.180 ;
        RECT 21.980 169.010 23.380 169.180 ;
        RECT 24.270 169.010 25.670 169.180 ;
        RECT 31.140 169.010 32.540 169.180 ;
        RECT 33.430 169.010 34.830 169.180 ;
        RECT 40.300 169.010 41.700 169.180 ;
        RECT 42.590 169.010 43.990 169.180 ;
        RECT 51.860 168.720 53.180 178.420 ;
        RECT 5.910 167.830 53.180 168.720 ;
        RECT 5.910 148.290 9.530 167.830 ;
        RECT 10.310 167.140 12.270 167.370 ;
        RECT 12.600 167.140 14.560 167.370 ;
        RECT 16.350 167.140 18.310 167.370 ;
        RECT 18.640 167.140 20.600 167.370 ;
        RECT 22.390 167.140 24.350 167.370 ;
        RECT 24.680 167.140 26.640 167.370 ;
        RECT 28.430 167.140 30.390 167.370 ;
        RECT 30.720 167.140 32.680 167.370 ;
        RECT 34.470 167.140 36.430 167.370 ;
        RECT 36.760 167.140 38.720 167.370 ;
        RECT 40.510 167.140 42.470 167.370 ;
        RECT 42.800 167.140 44.760 167.370 ;
        RECT 46.550 167.140 48.510 167.370 ;
        RECT 48.840 167.140 50.800 167.370 ;
        RECT 10.030 161.265 10.260 166.980 ;
        RECT 12.320 161.265 12.550 166.980 ;
        RECT 14.610 161.265 14.840 166.980 ;
        RECT 16.070 161.265 16.300 166.980 ;
        RECT 18.360 166.565 18.590 166.980 ;
        RECT 18.325 165.865 18.625 166.565 ;
        RECT 9.995 159.865 10.295 161.265 ;
        RECT 12.285 159.865 12.585 161.265 ;
        RECT 14.575 159.865 14.875 161.265 ;
        RECT 16.035 159.865 16.335 161.265 ;
        RECT 10.030 158.820 10.260 159.865 ;
        RECT 12.320 158.820 12.550 159.865 ;
        RECT 14.610 158.820 14.840 159.865 ;
        RECT 16.070 158.980 16.300 159.865 ;
        RECT 18.360 158.980 18.590 165.865 ;
        RECT 20.650 161.265 20.880 166.980 ;
        RECT 22.110 161.265 22.340 166.980 ;
        RECT 24.400 166.565 24.630 166.980 ;
        RECT 24.365 165.865 24.665 166.565 ;
        RECT 20.615 159.865 20.915 161.265 ;
        RECT 22.075 159.865 22.375 161.265 ;
        RECT 20.650 158.980 20.880 159.865 ;
        RECT 22.110 158.980 22.340 159.865 ;
        RECT 24.400 158.980 24.630 165.865 ;
        RECT 26.690 161.265 26.920 166.980 ;
        RECT 28.150 161.265 28.380 166.980 ;
        RECT 30.440 162.965 30.670 166.980 ;
        RECT 30.405 162.265 30.705 162.965 ;
        RECT 26.655 159.865 26.955 161.265 ;
        RECT 28.115 159.865 28.415 161.265 ;
        RECT 26.690 158.980 26.920 159.865 ;
        RECT 28.150 158.980 28.380 159.865 ;
        RECT 30.440 158.980 30.670 162.265 ;
        RECT 32.730 161.265 32.960 166.980 ;
        RECT 34.190 161.265 34.420 166.980 ;
        RECT 36.480 166.565 36.710 166.980 ;
        RECT 36.445 165.865 36.745 166.565 ;
        RECT 32.695 159.865 32.995 161.265 ;
        RECT 34.155 159.865 34.455 161.265 ;
        RECT 32.730 158.980 32.960 159.865 ;
        RECT 34.190 158.980 34.420 159.865 ;
        RECT 36.480 158.980 36.710 165.865 ;
        RECT 38.770 161.265 39.000 166.980 ;
        RECT 40.230 161.265 40.460 166.980 ;
        RECT 42.520 166.565 42.750 166.980 ;
        RECT 42.485 165.865 42.785 166.565 ;
        RECT 38.735 159.865 39.035 161.265 ;
        RECT 40.195 159.865 40.495 161.265 ;
        RECT 38.770 158.980 39.000 159.865 ;
        RECT 40.230 158.980 40.460 159.865 ;
        RECT 42.520 158.980 42.750 165.865 ;
        RECT 44.810 161.265 45.040 166.980 ;
        RECT 46.270 161.265 46.500 166.980 ;
        RECT 48.560 161.265 48.790 166.980 ;
        RECT 50.850 161.265 51.080 166.980 ;
        RECT 44.775 159.865 45.075 161.265 ;
        RECT 46.235 159.865 46.535 161.265 ;
        RECT 48.525 159.865 48.825 161.265 ;
        RECT 50.815 159.865 51.115 161.265 ;
        RECT 44.810 158.980 45.040 159.865 ;
        RECT 46.270 158.820 46.500 159.865 ;
        RECT 48.560 158.820 48.790 159.865 ;
        RECT 50.850 158.820 51.080 159.865 ;
        RECT 10.030 158.590 14.840 158.820 ;
        RECT 10.030 157.210 14.840 157.440 ;
        RECT 16.350 157.210 44.760 158.820 ;
        RECT 46.270 158.590 51.080 158.820 ;
        RECT 46.270 157.210 51.080 157.440 ;
        RECT 10.030 156.165 10.260 157.210 ;
        RECT 12.320 156.165 12.550 157.210 ;
        RECT 14.610 156.165 14.840 157.210 ;
        RECT 16.070 156.165 16.300 157.050 ;
        RECT 9.995 154.765 10.295 156.165 ;
        RECT 12.285 154.765 12.585 156.165 ;
        RECT 14.575 154.765 14.875 156.165 ;
        RECT 16.035 154.765 16.335 156.165 ;
        RECT 10.030 149.050 10.260 154.765 ;
        RECT 12.320 149.050 12.550 154.765 ;
        RECT 14.610 149.050 14.840 154.765 ;
        RECT 16.070 149.050 16.300 154.765 ;
        RECT 18.360 150.165 18.590 157.050 ;
        RECT 20.650 156.165 20.880 157.050 ;
        RECT 22.110 156.165 22.340 157.050 ;
        RECT 20.615 154.765 20.915 156.165 ;
        RECT 22.075 154.765 22.375 156.165 ;
        RECT 18.325 149.465 18.625 150.165 ;
        RECT 18.360 149.050 18.590 149.465 ;
        RECT 20.650 149.050 20.880 154.765 ;
        RECT 22.110 149.050 22.340 154.765 ;
        RECT 24.400 151.965 24.630 157.050 ;
        RECT 26.690 156.165 26.920 157.050 ;
        RECT 28.150 156.165 28.380 157.050 ;
        RECT 26.655 154.765 26.955 156.165 ;
        RECT 28.115 154.765 28.415 156.165 ;
        RECT 24.365 151.265 24.665 151.965 ;
        RECT 24.400 149.050 24.630 151.265 ;
        RECT 26.690 149.050 26.920 154.765 ;
        RECT 28.150 149.050 28.380 154.765 ;
        RECT 30.440 149.050 30.670 157.210 ;
        RECT 32.730 156.165 32.960 157.050 ;
        RECT 32.695 154.765 32.995 156.165 ;
        RECT 32.730 149.050 32.960 154.765 ;
        RECT 34.190 149.050 34.420 157.210 ;
        RECT 36.480 149.050 36.710 157.210 ;
        RECT 38.770 149.050 39.000 157.210 ;
        RECT 40.230 156.165 40.460 157.050 ;
        RECT 40.195 154.765 40.495 156.165 ;
        RECT 40.230 149.050 40.460 154.765 ;
        RECT 42.520 150.165 42.750 157.050 ;
        RECT 44.810 156.165 45.040 157.050 ;
        RECT 46.270 156.165 46.500 157.210 ;
        RECT 48.560 156.165 48.790 157.210 ;
        RECT 50.850 156.165 51.080 157.210 ;
        RECT 44.775 154.765 45.075 156.165 ;
        RECT 46.235 154.765 46.535 156.165 ;
        RECT 48.525 154.765 48.825 156.165 ;
        RECT 50.815 154.765 51.115 156.165 ;
        RECT 42.485 149.465 42.785 150.165 ;
        RECT 42.520 149.050 42.750 149.465 ;
        RECT 44.810 149.050 45.040 154.765 ;
        RECT 46.270 149.050 46.500 154.765 ;
        RECT 48.560 149.050 48.790 154.765 ;
        RECT 50.850 149.050 51.080 154.765 ;
        RECT 10.310 148.660 12.270 148.890 ;
        RECT 12.600 148.660 14.560 148.890 ;
        RECT 16.350 148.660 18.310 148.890 ;
        RECT 18.640 148.660 20.600 148.890 ;
        RECT 22.390 148.660 24.350 148.890 ;
        RECT 24.680 148.660 26.640 148.890 ;
        RECT 28.430 148.660 30.390 148.890 ;
        RECT 30.720 148.660 32.680 148.890 ;
        RECT 34.470 148.660 36.430 148.890 ;
        RECT 36.760 148.660 38.720 148.890 ;
        RECT 40.510 148.660 42.470 148.890 ;
        RECT 42.800 148.660 44.760 148.890 ;
        RECT 46.550 148.660 48.510 148.890 ;
        RECT 48.840 148.660 50.800 148.890 ;
        RECT 51.580 148.290 53.180 167.830 ;
        RECT 5.910 143.745 53.180 148.290 ;
        RECT 62.865 171.445 63.455 212.490 ;
        RECT 63.895 211.600 64.595 212.600 ;
        RECT 77.595 212.570 78.595 212.805 ;
        RECT 77.595 211.395 78.595 211.630 ;
        RECT 80.185 211.600 81.755 212.600 ;
        RECT 83.345 212.570 84.345 212.805 ;
        RECT 83.345 211.395 84.345 211.630 ;
        RECT 97.345 211.600 98.045 212.600 ;
        RECT 64.175 211.165 80.135 211.395 ;
        RECT 81.805 211.165 97.765 211.395 ;
        RECT 77.595 210.930 78.595 211.165 ;
        RECT 83.345 210.930 84.345 211.165 ;
        RECT 77.595 210.015 78.595 210.250 ;
        RECT 83.345 210.015 84.345 210.250 ;
        RECT 64.175 209.785 80.135 210.015 ;
        RECT 81.805 209.785 97.765 210.015 ;
        RECT 63.895 208.580 64.595 209.580 ;
        RECT 77.595 209.550 78.595 209.785 ;
        RECT 77.595 208.375 78.595 208.610 ;
        RECT 80.185 208.580 81.755 209.580 ;
        RECT 83.345 209.550 84.345 209.785 ;
        RECT 83.345 208.375 84.345 208.610 ;
        RECT 97.345 208.580 98.045 209.580 ;
        RECT 64.175 208.145 80.135 208.375 ;
        RECT 81.805 208.145 97.765 208.375 ;
        RECT 77.595 207.910 78.595 208.145 ;
        RECT 83.345 207.910 84.345 208.145 ;
        RECT 77.595 206.995 78.595 207.230 ;
        RECT 83.345 206.995 84.345 207.230 ;
        RECT 64.175 206.765 80.135 206.995 ;
        RECT 81.805 206.765 97.765 206.995 ;
        RECT 63.895 205.560 64.595 206.560 ;
        RECT 77.595 206.530 78.595 206.765 ;
        RECT 77.595 205.355 78.595 205.590 ;
        RECT 80.185 205.560 81.755 206.560 ;
        RECT 83.345 206.530 84.345 206.765 ;
        RECT 83.345 205.355 84.345 205.590 ;
        RECT 97.345 205.560 98.045 206.560 ;
        RECT 64.175 205.125 80.135 205.355 ;
        RECT 81.805 205.125 97.765 205.355 ;
        RECT 77.595 204.890 78.595 205.125 ;
        RECT 83.345 204.890 84.345 205.125 ;
        RECT 77.595 203.975 78.595 204.210 ;
        RECT 83.345 203.975 84.345 204.210 ;
        RECT 64.175 203.745 80.135 203.975 ;
        RECT 81.805 203.745 97.765 203.975 ;
        RECT 63.895 202.540 75.695 203.540 ;
        RECT 77.595 203.510 78.595 203.745 ;
        RECT 77.595 202.335 78.595 202.570 ;
        RECT 80.185 202.540 81.755 203.540 ;
        RECT 83.345 203.510 84.345 203.745 ;
        RECT 83.345 202.335 84.345 202.570 ;
        RECT 86.245 202.540 98.045 203.540 ;
        RECT 64.175 202.105 80.135 202.335 ;
        RECT 81.805 202.105 97.765 202.335 ;
        RECT 77.595 201.870 78.595 202.105 ;
        RECT 83.345 201.870 84.345 202.105 ;
        RECT 77.595 200.955 78.595 201.190 ;
        RECT 83.345 200.955 84.345 201.190 ;
        RECT 64.175 200.725 80.135 200.955 ;
        RECT 81.805 200.725 97.765 200.955 ;
        RECT 63.895 199.520 70.195 200.520 ;
        RECT 77.595 200.490 78.595 200.725 ;
        RECT 77.595 199.315 78.595 199.550 ;
        RECT 80.185 199.520 81.755 200.520 ;
        RECT 83.345 200.490 84.345 200.725 ;
        RECT 83.345 199.315 84.345 199.550 ;
        RECT 91.745 199.520 98.045 200.520 ;
        RECT 64.175 199.085 80.135 199.315 ;
        RECT 81.805 199.085 97.765 199.315 ;
        RECT 77.595 198.850 78.595 199.085 ;
        RECT 83.345 198.850 84.345 199.085 ;
        RECT 77.595 197.935 78.595 198.170 ;
        RECT 83.345 197.935 84.345 198.170 ;
        RECT 64.175 197.705 80.135 197.935 ;
        RECT 81.805 197.705 97.765 197.935 ;
        RECT 63.895 196.500 67.445 197.500 ;
        RECT 77.595 197.470 78.595 197.705 ;
        RECT 77.595 196.295 78.595 196.530 ;
        RECT 80.185 196.500 81.755 197.500 ;
        RECT 83.345 197.470 84.345 197.705 ;
        RECT 83.345 196.295 84.345 196.530 ;
        RECT 94.495 196.500 98.045 197.500 ;
        RECT 64.175 196.065 80.135 196.295 ;
        RECT 81.805 196.065 97.765 196.295 ;
        RECT 77.595 195.830 78.595 196.065 ;
        RECT 83.345 195.830 84.345 196.065 ;
        RECT 77.595 194.915 78.595 195.150 ;
        RECT 83.345 194.915 84.345 195.150 ;
        RECT 64.175 194.685 80.135 194.915 ;
        RECT 81.805 194.685 97.765 194.915 ;
        RECT 63.895 193.480 72.945 194.480 ;
        RECT 77.595 194.450 78.595 194.685 ;
        RECT 77.595 193.275 78.595 193.510 ;
        RECT 80.185 193.480 81.755 194.480 ;
        RECT 83.345 194.450 84.345 194.685 ;
        RECT 83.345 193.275 84.345 193.510 ;
        RECT 88.995 193.480 98.045 194.480 ;
        RECT 64.175 193.045 80.135 193.275 ;
        RECT 81.805 193.045 97.765 193.275 ;
        RECT 77.595 192.810 78.595 193.045 ;
        RECT 83.345 192.810 84.345 193.045 ;
        RECT 77.595 191.895 78.595 192.130 ;
        RECT 83.345 191.895 84.345 192.130 ;
        RECT 64.175 191.665 80.135 191.895 ;
        RECT 81.805 191.665 97.765 191.895 ;
        RECT 63.895 190.460 67.445 191.460 ;
        RECT 77.595 191.430 78.595 191.665 ;
        RECT 77.595 190.255 78.595 190.490 ;
        RECT 80.185 190.460 81.755 191.460 ;
        RECT 83.345 191.430 84.345 191.665 ;
        RECT 83.345 190.255 84.345 190.490 ;
        RECT 94.495 190.460 98.045 191.460 ;
        RECT 64.175 190.025 80.135 190.255 ;
        RECT 81.805 190.025 97.765 190.255 ;
        RECT 77.595 189.790 78.595 190.025 ;
        RECT 83.345 189.790 84.345 190.025 ;
        RECT 77.595 188.875 78.595 189.110 ;
        RECT 83.345 188.875 84.345 189.110 ;
        RECT 64.175 188.645 80.135 188.875 ;
        RECT 81.805 188.645 97.765 188.875 ;
        RECT 63.895 187.440 70.195 188.440 ;
        RECT 77.595 188.410 78.595 188.645 ;
        RECT 77.595 187.235 78.595 187.470 ;
        RECT 80.185 187.440 81.755 188.440 ;
        RECT 83.345 188.410 84.345 188.645 ;
        RECT 83.345 187.235 84.345 187.470 ;
        RECT 91.745 187.440 98.045 188.440 ;
        RECT 64.175 187.005 80.135 187.235 ;
        RECT 81.805 187.005 97.765 187.235 ;
        RECT 77.595 186.770 78.595 187.005 ;
        RECT 83.345 186.770 84.345 187.005 ;
        RECT 77.595 185.855 78.595 186.090 ;
        RECT 83.345 185.855 84.345 186.090 ;
        RECT 64.175 185.625 80.135 185.855 ;
        RECT 81.805 185.625 97.765 185.855 ;
        RECT 63.895 184.420 75.695 185.420 ;
        RECT 77.595 185.390 78.595 185.625 ;
        RECT 77.595 184.215 78.595 184.450 ;
        RECT 80.185 184.420 81.755 185.420 ;
        RECT 83.345 185.390 84.345 185.625 ;
        RECT 83.345 184.215 84.345 184.450 ;
        RECT 86.245 184.420 98.045 185.420 ;
        RECT 64.175 183.985 80.135 184.215 ;
        RECT 81.805 183.985 97.765 184.215 ;
        RECT 77.595 183.750 78.595 183.985 ;
        RECT 83.345 183.750 84.345 183.985 ;
        RECT 77.595 182.835 78.595 183.070 ;
        RECT 83.345 182.835 84.345 183.070 ;
        RECT 64.175 182.605 80.135 182.835 ;
        RECT 81.805 182.605 97.765 182.835 ;
        RECT 98.485 182.710 102.825 216.515 ;
        RECT 108.520 216.690 108.920 217.515 ;
        RECT 109.325 217.500 109.555 217.755 ;
        RECT 110.615 217.500 110.845 217.755 ;
        RECT 111.905 217.500 112.135 217.755 ;
        RECT 109.605 216.945 110.565 217.295 ;
        RECT 110.895 217.065 111.855 217.295 ;
        RECT 112.545 216.690 112.950 220.315 ;
        RECT 113.635 219.705 114.595 219.935 ;
        RECT 114.925 219.705 115.885 220.055 ;
        RECT 113.355 219.255 113.585 219.500 ;
        RECT 114.645 219.255 114.875 219.500 ;
        RECT 115.935 219.255 116.165 219.500 ;
        RECT 113.320 217.755 113.620 219.255 ;
        RECT 114.610 217.755 114.910 219.255 ;
        RECT 115.900 217.755 116.200 219.255 ;
        RECT 113.355 217.500 113.585 217.755 ;
        RECT 114.645 217.500 114.875 217.755 ;
        RECT 115.935 217.500 116.165 217.755 ;
        RECT 113.635 216.945 114.595 217.295 ;
        RECT 114.925 217.065 115.885 217.295 ;
        RECT 116.575 216.690 116.980 220.315 ;
        RECT 117.665 219.705 118.625 219.935 ;
        RECT 118.955 219.705 119.915 220.055 ;
        RECT 117.385 219.255 117.615 219.500 ;
        RECT 118.675 219.255 118.905 219.500 ;
        RECT 119.965 219.255 120.195 219.500 ;
        RECT 117.350 217.755 117.650 219.255 ;
        RECT 118.640 217.755 118.940 219.255 ;
        RECT 119.930 217.755 120.230 219.255 ;
        RECT 117.385 217.500 117.615 217.755 ;
        RECT 118.675 217.500 118.905 217.755 ;
        RECT 119.965 217.500 120.195 217.755 ;
        RECT 117.665 216.945 118.625 217.295 ;
        RECT 118.955 217.065 119.915 217.295 ;
        RECT 120.605 216.690 121.010 220.315 ;
        RECT 121.695 219.705 122.655 219.935 ;
        RECT 122.985 219.705 123.945 220.055 ;
        RECT 121.415 219.255 121.645 219.500 ;
        RECT 122.705 219.255 122.935 219.500 ;
        RECT 123.995 219.255 124.225 219.500 ;
        RECT 121.380 217.755 121.680 219.255 ;
        RECT 122.670 217.755 122.970 219.255 ;
        RECT 123.960 217.755 124.260 219.255 ;
        RECT 121.415 217.500 121.645 217.755 ;
        RECT 122.705 217.500 122.935 217.755 ;
        RECT 123.995 217.500 124.225 217.755 ;
        RECT 121.695 216.945 122.655 217.295 ;
        RECT 122.985 217.065 123.945 217.295 ;
        RECT 124.635 216.690 125.040 220.315 ;
        RECT 125.725 219.705 126.685 219.935 ;
        RECT 127.015 219.705 127.975 220.055 ;
        RECT 125.445 219.255 125.675 219.500 ;
        RECT 126.735 219.255 126.965 219.500 ;
        RECT 128.025 219.255 128.255 219.500 ;
        RECT 125.410 217.755 125.710 219.255 ;
        RECT 126.700 217.755 127.000 219.255 ;
        RECT 127.990 217.755 128.290 219.255 ;
        RECT 125.445 217.500 125.675 217.755 ;
        RECT 126.735 217.500 126.965 217.755 ;
        RECT 128.025 217.500 128.255 217.755 ;
        RECT 125.725 216.945 126.685 217.295 ;
        RECT 127.015 217.065 127.975 217.295 ;
        RECT 128.665 216.690 129.070 220.315 ;
        RECT 129.755 219.705 130.715 219.935 ;
        RECT 131.045 219.705 132.005 220.055 ;
        RECT 129.475 219.255 129.705 219.500 ;
        RECT 130.765 219.255 130.995 219.500 ;
        RECT 132.055 219.255 132.285 219.500 ;
        RECT 129.440 217.755 129.740 219.255 ;
        RECT 130.730 217.755 131.030 219.255 ;
        RECT 132.020 217.755 132.320 219.255 ;
        RECT 129.475 217.500 129.705 217.755 ;
        RECT 130.765 217.500 130.995 217.755 ;
        RECT 132.055 217.500 132.285 217.755 ;
        RECT 129.755 216.945 130.715 217.295 ;
        RECT 131.045 217.065 132.005 217.295 ;
        RECT 132.695 216.690 133.100 220.315 ;
        RECT 133.785 219.705 134.745 219.935 ;
        RECT 135.075 219.705 136.035 220.055 ;
        RECT 133.505 219.255 133.735 219.500 ;
        RECT 134.795 219.255 135.025 219.500 ;
        RECT 136.085 219.255 136.315 219.500 ;
        RECT 133.470 217.755 133.770 219.255 ;
        RECT 134.760 217.755 135.060 219.255 ;
        RECT 136.050 217.755 136.350 219.255 ;
        RECT 133.505 217.500 133.735 217.755 ;
        RECT 134.795 217.500 135.025 217.755 ;
        RECT 136.085 217.500 136.315 217.755 ;
        RECT 133.785 216.945 134.745 217.295 ;
        RECT 135.075 217.065 136.035 217.295 ;
        RECT 136.725 216.690 137.130 220.315 ;
        RECT 137.815 219.705 138.775 219.935 ;
        RECT 139.105 219.705 140.065 220.055 ;
        RECT 137.535 219.255 137.765 219.500 ;
        RECT 138.825 219.255 139.055 219.500 ;
        RECT 140.115 219.255 140.345 219.500 ;
        RECT 137.500 217.755 137.800 219.255 ;
        RECT 138.790 217.755 139.090 219.255 ;
        RECT 140.080 217.755 140.380 219.255 ;
        RECT 137.535 217.500 137.765 217.755 ;
        RECT 138.825 217.500 139.055 217.755 ;
        RECT 140.115 217.500 140.345 217.755 ;
        RECT 137.815 216.945 138.775 217.295 ;
        RECT 139.105 217.065 140.065 217.295 ;
        RECT 140.755 216.690 141.160 220.315 ;
        RECT 141.845 219.705 142.805 219.935 ;
        RECT 143.135 219.705 144.095 220.055 ;
        RECT 141.565 219.255 141.795 219.500 ;
        RECT 142.855 219.255 143.085 219.500 ;
        RECT 144.145 219.255 144.375 219.500 ;
        RECT 141.530 217.755 141.830 219.255 ;
        RECT 142.820 217.755 143.120 219.255 ;
        RECT 144.110 217.755 144.410 219.255 ;
        RECT 141.565 217.500 141.795 217.755 ;
        RECT 142.855 217.500 143.085 217.755 ;
        RECT 144.145 217.500 144.375 217.755 ;
        RECT 141.845 216.945 142.805 217.295 ;
        RECT 143.135 217.065 144.095 217.295 ;
        RECT 144.785 216.690 145.190 220.315 ;
        RECT 145.875 219.705 146.835 219.935 ;
        RECT 147.165 219.705 148.125 220.055 ;
        RECT 145.595 219.255 145.825 219.500 ;
        RECT 146.885 219.255 147.115 219.500 ;
        RECT 148.175 219.255 148.405 219.500 ;
        RECT 145.560 217.755 145.860 219.255 ;
        RECT 146.850 217.755 147.150 219.255 ;
        RECT 148.140 217.755 148.440 219.255 ;
        RECT 145.595 217.500 145.825 217.755 ;
        RECT 146.885 217.500 147.115 217.755 ;
        RECT 148.175 217.500 148.405 217.755 ;
        RECT 145.875 216.945 146.835 217.295 ;
        RECT 147.165 217.065 148.125 217.295 ;
        RECT 148.815 216.690 149.220 220.315 ;
        RECT 149.905 219.705 150.865 219.935 ;
        RECT 151.195 219.705 152.155 220.055 ;
        RECT 149.625 219.255 149.855 219.500 ;
        RECT 150.915 219.255 151.145 219.500 ;
        RECT 152.205 219.255 152.435 219.500 ;
        RECT 149.590 217.755 149.890 219.255 ;
        RECT 150.880 217.755 151.180 219.255 ;
        RECT 152.170 217.755 152.470 219.255 ;
        RECT 149.625 217.500 149.855 217.755 ;
        RECT 150.915 217.500 151.145 217.755 ;
        RECT 152.205 217.500 152.435 217.755 ;
        RECT 149.905 216.945 150.865 217.295 ;
        RECT 151.195 217.065 152.155 217.295 ;
        RECT 152.845 216.690 153.245 220.315 ;
        RECT 108.520 216.290 153.245 216.690 ;
        RECT 106.415 213.340 153.245 213.740 ;
        RECT 106.415 210.540 108.915 213.340 ;
        RECT 109.605 212.735 110.565 212.965 ;
        RECT 110.895 212.735 111.855 212.965 ;
        RECT 108.515 203.720 108.915 210.540 ;
        RECT 109.325 205.495 109.555 212.530 ;
        RECT 110.615 211.190 110.845 212.530 ;
        RECT 110.580 209.690 110.880 211.190 ;
        RECT 109.290 204.795 109.590 205.495 ;
        RECT 109.325 204.530 109.555 204.795 ;
        RECT 110.615 204.530 110.845 209.690 ;
        RECT 111.905 206.705 112.135 212.530 ;
        RECT 111.870 206.005 112.170 206.705 ;
        RECT 111.905 204.530 112.135 206.005 ;
        RECT 109.605 203.995 110.565 204.325 ;
        RECT 110.895 203.995 111.855 204.325 ;
        RECT 112.545 203.720 112.945 213.340 ;
        RECT 113.635 212.735 114.595 212.965 ;
        RECT 114.925 212.735 115.885 212.965 ;
        RECT 113.355 205.495 113.585 212.530 ;
        RECT 114.645 211.190 114.875 212.530 ;
        RECT 114.610 209.690 114.910 211.190 ;
        RECT 113.320 204.795 113.620 205.495 ;
        RECT 113.355 204.530 113.585 204.795 ;
        RECT 114.645 204.530 114.875 209.690 ;
        RECT 115.935 206.705 116.165 212.530 ;
        RECT 115.900 206.005 116.200 206.705 ;
        RECT 115.935 204.530 116.165 206.005 ;
        RECT 113.635 203.995 114.595 204.325 ;
        RECT 114.925 203.995 115.885 204.325 ;
        RECT 116.575 203.720 116.975 213.340 ;
        RECT 117.665 212.735 118.625 212.965 ;
        RECT 118.955 212.735 119.915 212.965 ;
        RECT 117.385 205.495 117.615 212.530 ;
        RECT 118.675 211.190 118.905 212.530 ;
        RECT 118.640 209.690 118.940 211.190 ;
        RECT 117.350 204.795 117.650 205.495 ;
        RECT 117.385 204.530 117.615 204.795 ;
        RECT 118.675 204.530 118.905 209.690 ;
        RECT 119.965 206.705 120.195 212.530 ;
        RECT 119.930 206.005 120.230 206.705 ;
        RECT 119.965 204.530 120.195 206.005 ;
        RECT 117.665 203.995 118.625 204.325 ;
        RECT 118.955 203.995 119.915 204.325 ;
        RECT 120.605 203.720 121.005 213.340 ;
        RECT 121.695 212.735 122.655 212.965 ;
        RECT 122.985 212.735 123.945 212.965 ;
        RECT 121.415 205.495 121.645 212.530 ;
        RECT 122.705 211.190 122.935 212.530 ;
        RECT 122.670 209.690 122.970 211.190 ;
        RECT 121.380 204.795 121.680 205.495 ;
        RECT 121.415 204.530 121.645 204.795 ;
        RECT 122.705 204.530 122.935 209.690 ;
        RECT 123.995 206.705 124.225 212.530 ;
        RECT 123.960 206.005 124.260 206.705 ;
        RECT 123.995 204.530 124.225 206.005 ;
        RECT 121.695 203.995 122.655 204.325 ;
        RECT 122.985 203.995 123.945 204.325 ;
        RECT 124.635 203.720 125.035 213.340 ;
        RECT 125.725 212.735 126.685 212.965 ;
        RECT 127.015 212.735 127.975 212.965 ;
        RECT 125.445 205.495 125.675 212.530 ;
        RECT 126.735 211.190 126.965 212.530 ;
        RECT 126.700 209.690 127.000 211.190 ;
        RECT 125.410 204.795 125.710 205.495 ;
        RECT 125.445 204.530 125.675 204.795 ;
        RECT 126.735 204.530 126.965 209.690 ;
        RECT 128.025 206.705 128.255 212.530 ;
        RECT 127.990 206.005 128.290 206.705 ;
        RECT 128.025 204.530 128.255 206.005 ;
        RECT 125.725 203.995 126.685 204.325 ;
        RECT 127.015 203.995 127.975 204.325 ;
        RECT 128.665 203.720 129.065 213.340 ;
        RECT 129.755 212.735 130.715 212.965 ;
        RECT 131.045 212.735 132.005 212.965 ;
        RECT 129.475 205.495 129.705 212.530 ;
        RECT 130.765 211.190 130.995 212.530 ;
        RECT 130.730 209.690 131.030 211.190 ;
        RECT 129.440 204.795 129.740 205.495 ;
        RECT 129.475 204.530 129.705 204.795 ;
        RECT 130.765 204.530 130.995 209.690 ;
        RECT 132.055 206.705 132.285 212.530 ;
        RECT 132.020 206.005 132.320 206.705 ;
        RECT 132.055 204.530 132.285 206.005 ;
        RECT 129.755 203.995 130.715 204.325 ;
        RECT 131.045 203.995 132.005 204.325 ;
        RECT 132.695 203.720 133.095 213.340 ;
        RECT 133.785 212.735 134.745 212.965 ;
        RECT 135.075 212.735 136.035 212.965 ;
        RECT 133.505 205.495 133.735 212.530 ;
        RECT 134.795 211.190 135.025 212.530 ;
        RECT 134.760 209.690 135.060 211.190 ;
        RECT 133.470 204.795 133.770 205.495 ;
        RECT 133.505 204.530 133.735 204.795 ;
        RECT 134.795 204.530 135.025 209.690 ;
        RECT 136.085 206.705 136.315 212.530 ;
        RECT 136.050 206.005 136.350 206.705 ;
        RECT 136.085 204.530 136.315 206.005 ;
        RECT 133.785 203.995 134.745 204.325 ;
        RECT 135.075 203.995 136.035 204.325 ;
        RECT 136.725 203.720 137.125 213.340 ;
        RECT 137.815 212.735 138.775 212.965 ;
        RECT 139.105 212.735 140.065 212.965 ;
        RECT 137.535 205.495 137.765 212.530 ;
        RECT 138.825 211.190 139.055 212.530 ;
        RECT 138.790 209.690 139.090 211.190 ;
        RECT 137.500 204.795 137.800 205.495 ;
        RECT 137.535 204.530 137.765 204.795 ;
        RECT 138.825 204.530 139.055 209.690 ;
        RECT 140.115 206.705 140.345 212.530 ;
        RECT 140.080 206.005 140.380 206.705 ;
        RECT 140.115 204.530 140.345 206.005 ;
        RECT 137.815 203.995 138.775 204.325 ;
        RECT 139.105 203.995 140.065 204.325 ;
        RECT 140.755 203.720 141.155 213.340 ;
        RECT 141.845 212.735 142.805 212.965 ;
        RECT 143.135 212.735 144.095 212.965 ;
        RECT 141.565 205.495 141.795 212.530 ;
        RECT 142.855 211.190 143.085 212.530 ;
        RECT 142.820 209.690 143.120 211.190 ;
        RECT 141.530 204.795 141.830 205.495 ;
        RECT 141.565 204.530 141.795 204.795 ;
        RECT 142.855 204.530 143.085 209.690 ;
        RECT 144.145 206.705 144.375 212.530 ;
        RECT 144.110 206.005 144.410 206.705 ;
        RECT 144.145 204.530 144.375 206.005 ;
        RECT 141.845 203.995 142.805 204.325 ;
        RECT 143.135 203.995 144.095 204.325 ;
        RECT 144.785 203.720 145.185 213.340 ;
        RECT 145.875 212.735 146.835 212.965 ;
        RECT 147.165 212.735 148.125 212.965 ;
        RECT 145.595 205.495 145.825 212.530 ;
        RECT 146.885 211.190 147.115 212.530 ;
        RECT 146.850 209.690 147.150 211.190 ;
        RECT 145.560 204.795 145.860 205.495 ;
        RECT 145.595 204.530 145.825 204.795 ;
        RECT 146.885 204.530 147.115 209.690 ;
        RECT 148.175 206.705 148.405 212.530 ;
        RECT 148.140 206.005 148.440 206.705 ;
        RECT 148.175 204.530 148.405 206.005 ;
        RECT 145.875 203.995 146.835 204.325 ;
        RECT 147.165 203.995 148.125 204.325 ;
        RECT 148.815 203.720 149.215 213.340 ;
        RECT 149.905 212.735 150.865 212.965 ;
        RECT 151.195 212.735 152.155 212.965 ;
        RECT 149.625 205.495 149.855 212.530 ;
        RECT 150.915 211.190 151.145 212.530 ;
        RECT 150.880 209.690 151.180 211.190 ;
        RECT 149.590 204.795 149.890 205.495 ;
        RECT 149.625 204.530 149.855 204.795 ;
        RECT 150.915 204.530 151.145 209.690 ;
        RECT 152.205 206.705 152.435 212.530 ;
        RECT 152.170 206.005 152.470 206.705 ;
        RECT 152.205 204.530 152.435 206.005 ;
        RECT 149.905 203.995 150.865 204.325 ;
        RECT 151.195 203.995 152.155 204.325 ;
        RECT 152.845 203.720 153.245 213.340 ;
        RECT 108.515 203.320 153.245 203.720 ;
        RECT 165.150 201.250 239.210 201.730 ;
        RECT 108.515 200.625 153.245 201.025 ;
        RECT 168.440 200.850 168.760 201.110 ;
        RECT 178.100 201.050 178.420 201.110 ;
        RECT 179.495 201.050 179.785 201.095 ;
        RECT 178.100 200.910 179.785 201.050 ;
        RECT 178.100 200.850 178.420 200.910 ;
        RECT 179.495 200.865 179.785 200.910 ;
        RECT 187.760 201.050 188.080 201.110 ;
        RECT 188.695 201.050 188.985 201.095 ;
        RECT 187.760 200.910 188.985 201.050 ;
        RECT 187.760 200.850 188.080 200.910 ;
        RECT 188.695 200.865 188.985 200.910 ;
        RECT 197.420 201.050 197.740 201.110 ;
        RECT 198.355 201.050 198.645 201.095 ;
        RECT 197.420 200.910 198.645 201.050 ;
        RECT 197.420 200.850 197.740 200.910 ;
        RECT 198.355 200.865 198.645 200.910 ;
        RECT 207.080 201.050 207.400 201.110 ;
        RECT 208.015 201.050 208.305 201.095 ;
        RECT 207.080 200.910 208.305 201.050 ;
        RECT 207.080 200.850 207.400 200.910 ;
        RECT 208.015 200.865 208.305 200.910 ;
        RECT 216.740 201.050 217.060 201.110 ;
        RECT 218.135 201.050 218.425 201.095 ;
        RECT 216.740 200.910 218.425 201.050 ;
        RECT 216.740 200.850 217.060 200.910 ;
        RECT 218.135 200.865 218.425 200.910 ;
        RECT 226.400 201.050 226.720 201.110 ;
        RECT 227.795 201.050 228.085 201.095 ;
        RECT 226.400 200.910 228.085 201.050 ;
        RECT 226.400 200.850 226.720 200.910 ;
        RECT 227.795 200.865 228.085 200.910 ;
        RECT 236.060 201.050 236.380 201.110 ;
        RECT 236.995 201.050 237.285 201.095 ;
        RECT 236.060 200.910 237.285 201.050 ;
        RECT 236.060 200.850 236.380 200.910 ;
        RECT 236.995 200.865 237.285 200.910 ;
        RECT 108.515 195.095 108.915 200.625 ;
        RECT 109.735 200.250 110.435 200.320 ;
        RECT 111.025 200.250 111.725 200.320 ;
        RECT 109.605 200.020 110.565 200.250 ;
        RECT 110.895 200.020 111.855 200.250 ;
        RECT 109.325 199.635 109.555 199.860 ;
        RECT 109.290 198.935 109.590 199.635 ;
        RECT 110.615 198.955 110.845 199.860 ;
        RECT 111.905 199.635 112.135 199.860 ;
        RECT 109.325 195.860 109.555 198.935 ;
        RECT 110.580 196.855 110.880 198.955 ;
        RECT 111.870 198.935 112.170 199.635 ;
        RECT 110.615 195.860 110.845 196.855 ;
        RECT 111.905 195.860 112.135 198.935 ;
        RECT 109.605 195.470 110.565 195.700 ;
        RECT 110.895 195.470 111.855 195.700 ;
        RECT 112.545 195.095 112.945 200.625 ;
        RECT 113.765 200.250 114.465 200.320 ;
        RECT 115.055 200.250 115.755 200.320 ;
        RECT 113.635 200.020 114.595 200.250 ;
        RECT 114.925 200.020 115.885 200.250 ;
        RECT 113.355 199.635 113.585 199.860 ;
        RECT 113.320 198.935 113.620 199.635 ;
        RECT 114.645 198.955 114.875 199.860 ;
        RECT 115.935 199.635 116.165 199.860 ;
        RECT 113.355 195.860 113.585 198.935 ;
        RECT 114.610 196.855 114.910 198.955 ;
        RECT 115.900 198.935 116.200 199.635 ;
        RECT 114.645 195.860 114.875 196.855 ;
        RECT 115.935 195.860 116.165 198.935 ;
        RECT 113.635 195.470 114.595 195.700 ;
        RECT 114.925 195.470 115.885 195.700 ;
        RECT 116.575 195.095 116.975 200.625 ;
        RECT 117.795 200.250 118.495 200.320 ;
        RECT 119.085 200.250 119.785 200.320 ;
        RECT 117.665 200.020 118.625 200.250 ;
        RECT 118.955 200.020 119.915 200.250 ;
        RECT 117.385 199.635 117.615 199.860 ;
        RECT 117.350 198.935 117.650 199.635 ;
        RECT 118.675 198.955 118.905 199.860 ;
        RECT 119.965 199.635 120.195 199.860 ;
        RECT 117.385 195.860 117.615 198.935 ;
        RECT 118.640 196.855 118.940 198.955 ;
        RECT 119.930 198.935 120.230 199.635 ;
        RECT 118.675 195.860 118.905 196.855 ;
        RECT 119.965 195.860 120.195 198.935 ;
        RECT 117.665 195.470 118.625 195.700 ;
        RECT 118.955 195.470 119.915 195.700 ;
        RECT 120.605 195.095 121.005 200.625 ;
        RECT 121.825 200.250 122.525 200.320 ;
        RECT 123.115 200.250 123.815 200.320 ;
        RECT 121.695 200.020 122.655 200.250 ;
        RECT 122.985 200.020 123.945 200.250 ;
        RECT 121.415 199.635 121.645 199.860 ;
        RECT 121.380 198.935 121.680 199.635 ;
        RECT 122.705 198.955 122.935 199.860 ;
        RECT 123.995 199.635 124.225 199.860 ;
        RECT 121.415 195.860 121.645 198.935 ;
        RECT 122.670 196.855 122.970 198.955 ;
        RECT 123.960 198.935 124.260 199.635 ;
        RECT 122.705 195.860 122.935 196.855 ;
        RECT 123.995 195.860 124.225 198.935 ;
        RECT 121.695 195.470 122.655 195.700 ;
        RECT 122.985 195.470 123.945 195.700 ;
        RECT 124.635 195.095 125.035 200.625 ;
        RECT 125.855 200.250 126.555 200.320 ;
        RECT 127.145 200.250 127.845 200.320 ;
        RECT 125.725 200.020 126.685 200.250 ;
        RECT 127.015 200.020 127.975 200.250 ;
        RECT 125.445 199.635 125.675 199.860 ;
        RECT 125.410 198.935 125.710 199.635 ;
        RECT 126.735 198.955 126.965 199.860 ;
        RECT 128.025 199.635 128.255 199.860 ;
        RECT 125.445 195.860 125.675 198.935 ;
        RECT 126.700 196.855 127.000 198.955 ;
        RECT 127.990 198.935 128.290 199.635 ;
        RECT 126.735 195.860 126.965 196.855 ;
        RECT 128.025 195.860 128.255 198.935 ;
        RECT 125.725 195.470 126.685 195.700 ;
        RECT 127.015 195.470 127.975 195.700 ;
        RECT 128.665 195.095 129.065 200.625 ;
        RECT 129.885 200.250 130.585 200.320 ;
        RECT 131.175 200.250 131.875 200.320 ;
        RECT 129.755 200.020 130.715 200.250 ;
        RECT 131.045 200.020 132.005 200.250 ;
        RECT 129.475 199.635 129.705 199.860 ;
        RECT 129.440 198.935 129.740 199.635 ;
        RECT 130.765 198.955 130.995 199.860 ;
        RECT 132.055 199.635 132.285 199.860 ;
        RECT 129.475 195.860 129.705 198.935 ;
        RECT 130.730 196.855 131.030 198.955 ;
        RECT 132.020 198.935 132.320 199.635 ;
        RECT 130.765 195.860 130.995 196.855 ;
        RECT 132.055 195.860 132.285 198.935 ;
        RECT 129.755 195.470 130.715 195.700 ;
        RECT 131.045 195.470 132.005 195.700 ;
        RECT 132.695 195.095 133.095 200.625 ;
        RECT 133.915 200.250 134.615 200.320 ;
        RECT 135.205 200.250 135.905 200.320 ;
        RECT 133.785 200.020 134.745 200.250 ;
        RECT 135.075 200.020 136.035 200.250 ;
        RECT 133.505 199.635 133.735 199.860 ;
        RECT 133.470 198.935 133.770 199.635 ;
        RECT 134.795 198.955 135.025 199.860 ;
        RECT 136.085 199.635 136.315 199.860 ;
        RECT 133.505 195.860 133.735 198.935 ;
        RECT 134.760 196.855 135.060 198.955 ;
        RECT 136.050 198.935 136.350 199.635 ;
        RECT 134.795 195.860 135.025 196.855 ;
        RECT 136.085 195.860 136.315 198.935 ;
        RECT 133.785 195.470 134.745 195.700 ;
        RECT 135.075 195.470 136.035 195.700 ;
        RECT 136.725 195.095 137.125 200.625 ;
        RECT 137.945 200.250 138.645 200.320 ;
        RECT 139.235 200.250 139.935 200.320 ;
        RECT 137.815 200.020 138.775 200.250 ;
        RECT 139.105 200.020 140.065 200.250 ;
        RECT 137.535 199.635 137.765 199.860 ;
        RECT 137.500 198.935 137.800 199.635 ;
        RECT 138.825 198.955 139.055 199.860 ;
        RECT 140.115 199.635 140.345 199.860 ;
        RECT 137.535 195.860 137.765 198.935 ;
        RECT 138.790 196.855 139.090 198.955 ;
        RECT 140.080 198.935 140.380 199.635 ;
        RECT 138.825 195.860 139.055 196.855 ;
        RECT 140.115 195.860 140.345 198.935 ;
        RECT 137.815 195.470 138.775 195.700 ;
        RECT 139.105 195.470 140.065 195.700 ;
        RECT 140.755 195.095 141.155 200.625 ;
        RECT 141.975 200.250 142.675 200.320 ;
        RECT 143.265 200.250 143.965 200.320 ;
        RECT 141.845 200.020 142.805 200.250 ;
        RECT 143.135 200.020 144.095 200.250 ;
        RECT 141.565 199.635 141.795 199.860 ;
        RECT 141.530 198.935 141.830 199.635 ;
        RECT 142.855 198.955 143.085 199.860 ;
        RECT 144.145 199.635 144.375 199.860 ;
        RECT 141.565 195.860 141.795 198.935 ;
        RECT 142.820 196.855 143.120 198.955 ;
        RECT 144.110 198.935 144.410 199.635 ;
        RECT 142.855 195.860 143.085 196.855 ;
        RECT 144.145 195.860 144.375 198.935 ;
        RECT 141.845 195.470 142.805 195.700 ;
        RECT 143.135 195.470 144.095 195.700 ;
        RECT 144.785 195.095 145.185 200.625 ;
        RECT 146.005 200.250 146.705 200.320 ;
        RECT 147.295 200.250 147.995 200.320 ;
        RECT 145.875 200.020 146.835 200.250 ;
        RECT 147.165 200.020 148.125 200.250 ;
        RECT 145.595 199.635 145.825 199.860 ;
        RECT 145.560 198.935 145.860 199.635 ;
        RECT 146.885 198.955 147.115 199.860 ;
        RECT 148.175 199.635 148.405 199.860 ;
        RECT 145.595 195.860 145.825 198.935 ;
        RECT 146.850 196.855 147.150 198.955 ;
        RECT 148.140 198.935 148.440 199.635 ;
        RECT 146.885 195.860 147.115 196.855 ;
        RECT 148.175 195.860 148.405 198.935 ;
        RECT 145.875 195.470 146.835 195.700 ;
        RECT 147.165 195.470 148.125 195.700 ;
        RECT 148.815 195.095 149.215 200.625 ;
        RECT 150.035 200.250 150.735 200.320 ;
        RECT 151.325 200.250 152.025 200.320 ;
        RECT 149.905 200.020 150.865 200.250 ;
        RECT 151.195 200.020 152.155 200.250 ;
        RECT 149.625 199.635 149.855 199.860 ;
        RECT 149.590 198.935 149.890 199.635 ;
        RECT 150.915 198.955 151.145 199.860 ;
        RECT 152.205 199.635 152.435 199.860 ;
        RECT 149.625 195.860 149.855 198.935 ;
        RECT 150.880 196.855 151.180 198.955 ;
        RECT 152.170 198.935 152.470 199.635 ;
        RECT 150.915 195.860 151.145 196.855 ;
        RECT 152.205 195.860 152.435 198.935 ;
        RECT 149.905 195.470 150.865 195.700 ;
        RECT 151.195 195.470 152.155 195.700 ;
        RECT 152.845 195.095 153.245 200.625 ;
        RECT 166.600 200.030 166.920 200.090 ;
        RECT 170.755 200.030 171.045 200.075 ;
        RECT 166.600 199.890 171.045 200.030 ;
        RECT 166.600 199.830 166.920 199.890 ;
        RECT 170.755 199.845 171.045 199.890 ;
        RECT 178.560 199.830 178.880 200.090 ;
        RECT 189.600 199.830 189.920 200.090 ;
        RECT 199.260 199.830 199.580 200.090 ;
        RECT 208.920 199.830 209.240 200.090 ;
        RECT 226.860 199.830 227.180 200.090 ;
        RECT 236.060 199.830 236.380 200.090 ;
        RECT 169.820 199.490 170.140 199.750 ;
        RECT 217.200 199.690 217.520 199.750 ;
        RECT 217.675 199.690 217.965 199.735 ;
        RECT 217.200 199.550 217.965 199.690 ;
        RECT 217.200 199.490 217.520 199.550 ;
        RECT 217.675 199.505 217.965 199.550 ;
        RECT 171.675 199.350 171.965 199.395 ;
        RECT 172.120 199.350 172.440 199.410 ;
        RECT 182.240 199.350 182.560 199.410 ;
        RECT 171.675 199.210 182.560 199.350 ;
        RECT 171.675 199.165 171.965 199.210 ;
        RECT 172.120 199.150 172.440 199.210 ;
        RECT 182.240 199.150 182.560 199.210 ;
        RECT 165.150 198.530 239.990 199.010 ;
        RECT 165.150 195.810 239.210 196.290 ;
        RECT 189.155 195.610 189.445 195.655 ;
        RECT 189.600 195.610 189.920 195.670 ;
        RECT 189.155 195.470 189.920 195.610 ;
        RECT 189.155 195.425 189.445 195.470 ;
        RECT 189.600 195.410 189.920 195.470 ;
        RECT 190.150 195.470 191.670 195.610 ;
        RECT 190.150 195.270 190.290 195.470 ;
        RECT 108.515 194.695 153.245 195.095 ;
        RECT 108.515 185.165 108.915 194.695 ;
        RECT 109.605 194.320 110.305 194.390 ;
        RECT 111.155 194.320 111.855 194.390 ;
        RECT 109.605 194.090 110.565 194.320 ;
        RECT 110.895 194.090 111.855 194.320 ;
        RECT 109.325 192.835 109.555 193.930 ;
        RECT 109.290 191.335 109.590 192.835 ;
        RECT 109.325 185.930 109.555 191.335 ;
        RECT 110.615 189.090 110.845 193.930 ;
        RECT 111.905 192.835 112.135 193.930 ;
        RECT 111.870 191.335 112.170 192.835 ;
        RECT 110.580 187.590 110.880 189.090 ;
        RECT 110.615 185.930 110.845 187.590 ;
        RECT 111.905 185.930 112.135 191.335 ;
        RECT 109.605 185.540 110.565 185.770 ;
        RECT 110.895 185.540 111.855 185.770 ;
        RECT 112.545 185.165 112.945 194.695 ;
        RECT 113.635 194.320 114.335 194.390 ;
        RECT 115.185 194.320 115.885 194.390 ;
        RECT 113.635 194.090 114.595 194.320 ;
        RECT 114.925 194.090 115.885 194.320 ;
        RECT 113.355 192.835 113.585 193.930 ;
        RECT 113.320 191.335 113.620 192.835 ;
        RECT 113.355 185.930 113.585 191.335 ;
        RECT 114.645 189.090 114.875 193.930 ;
        RECT 115.935 192.835 116.165 193.930 ;
        RECT 115.900 191.335 116.200 192.835 ;
        RECT 114.610 187.590 114.910 189.090 ;
        RECT 114.645 185.930 114.875 187.590 ;
        RECT 115.935 185.930 116.165 191.335 ;
        RECT 113.635 185.540 114.595 185.770 ;
        RECT 114.925 185.540 115.885 185.770 ;
        RECT 116.575 185.165 116.975 194.695 ;
        RECT 117.665 194.320 118.365 194.390 ;
        RECT 119.215 194.320 119.915 194.390 ;
        RECT 117.665 194.090 118.625 194.320 ;
        RECT 118.955 194.090 119.915 194.320 ;
        RECT 117.385 192.835 117.615 193.930 ;
        RECT 117.350 191.335 117.650 192.835 ;
        RECT 117.385 185.930 117.615 191.335 ;
        RECT 118.675 189.090 118.905 193.930 ;
        RECT 119.965 192.835 120.195 193.930 ;
        RECT 119.930 191.335 120.230 192.835 ;
        RECT 118.640 187.590 118.940 189.090 ;
        RECT 118.675 185.930 118.905 187.590 ;
        RECT 119.965 185.930 120.195 191.335 ;
        RECT 117.665 185.540 118.625 185.770 ;
        RECT 118.955 185.540 119.915 185.770 ;
        RECT 120.605 185.165 121.005 194.695 ;
        RECT 121.695 194.320 122.395 194.390 ;
        RECT 123.245 194.320 123.945 194.390 ;
        RECT 121.695 194.090 122.655 194.320 ;
        RECT 122.985 194.090 123.945 194.320 ;
        RECT 121.415 192.835 121.645 193.930 ;
        RECT 121.380 191.335 121.680 192.835 ;
        RECT 121.415 185.930 121.645 191.335 ;
        RECT 122.705 189.090 122.935 193.930 ;
        RECT 123.995 192.835 124.225 193.930 ;
        RECT 123.960 191.335 124.260 192.835 ;
        RECT 122.670 187.590 122.970 189.090 ;
        RECT 122.705 185.930 122.935 187.590 ;
        RECT 123.995 185.930 124.225 191.335 ;
        RECT 121.695 185.540 122.655 185.770 ;
        RECT 122.985 185.540 123.945 185.770 ;
        RECT 124.635 185.165 125.035 194.695 ;
        RECT 125.725 194.320 126.425 194.390 ;
        RECT 127.275 194.320 127.975 194.390 ;
        RECT 125.725 194.090 126.685 194.320 ;
        RECT 127.015 194.090 127.975 194.320 ;
        RECT 125.445 192.835 125.675 193.930 ;
        RECT 125.410 191.335 125.710 192.835 ;
        RECT 125.445 185.930 125.675 191.335 ;
        RECT 126.735 189.090 126.965 193.930 ;
        RECT 128.025 192.835 128.255 193.930 ;
        RECT 127.990 191.335 128.290 192.835 ;
        RECT 126.700 187.590 127.000 189.090 ;
        RECT 126.735 185.930 126.965 187.590 ;
        RECT 128.025 185.930 128.255 191.335 ;
        RECT 125.725 185.540 126.685 185.770 ;
        RECT 127.015 185.540 127.975 185.770 ;
        RECT 128.665 185.165 129.065 194.695 ;
        RECT 129.755 194.320 130.455 194.390 ;
        RECT 131.305 194.320 132.005 194.390 ;
        RECT 129.755 194.090 130.715 194.320 ;
        RECT 131.045 194.090 132.005 194.320 ;
        RECT 129.475 192.835 129.705 193.930 ;
        RECT 129.440 191.335 129.740 192.835 ;
        RECT 129.475 185.930 129.705 191.335 ;
        RECT 130.765 189.090 130.995 193.930 ;
        RECT 132.055 192.835 132.285 193.930 ;
        RECT 132.020 191.335 132.320 192.835 ;
        RECT 130.730 187.590 131.030 189.090 ;
        RECT 130.765 185.930 130.995 187.590 ;
        RECT 132.055 185.930 132.285 191.335 ;
        RECT 129.755 185.540 130.715 185.770 ;
        RECT 131.045 185.540 132.005 185.770 ;
        RECT 132.695 185.165 133.095 194.695 ;
        RECT 133.785 194.320 134.485 194.390 ;
        RECT 135.335 194.320 136.035 194.390 ;
        RECT 133.785 194.090 134.745 194.320 ;
        RECT 135.075 194.090 136.035 194.320 ;
        RECT 133.505 192.835 133.735 193.930 ;
        RECT 133.470 191.335 133.770 192.835 ;
        RECT 133.505 185.930 133.735 191.335 ;
        RECT 134.795 189.090 135.025 193.930 ;
        RECT 136.085 192.835 136.315 193.930 ;
        RECT 136.050 191.335 136.350 192.835 ;
        RECT 134.760 187.590 135.060 189.090 ;
        RECT 134.795 185.930 135.025 187.590 ;
        RECT 136.085 185.930 136.315 191.335 ;
        RECT 133.785 185.540 134.745 185.770 ;
        RECT 135.075 185.540 136.035 185.770 ;
        RECT 136.725 185.165 137.125 194.695 ;
        RECT 137.815 194.320 138.515 194.390 ;
        RECT 139.365 194.320 140.065 194.390 ;
        RECT 137.815 194.090 138.775 194.320 ;
        RECT 139.105 194.090 140.065 194.320 ;
        RECT 137.535 192.835 137.765 193.930 ;
        RECT 137.500 191.335 137.800 192.835 ;
        RECT 137.535 185.930 137.765 191.335 ;
        RECT 138.825 189.090 139.055 193.930 ;
        RECT 140.115 192.835 140.345 193.930 ;
        RECT 140.080 191.335 140.380 192.835 ;
        RECT 138.790 187.590 139.090 189.090 ;
        RECT 138.825 185.930 139.055 187.590 ;
        RECT 140.115 185.930 140.345 191.335 ;
        RECT 137.815 185.540 138.775 185.770 ;
        RECT 139.105 185.540 140.065 185.770 ;
        RECT 140.755 185.165 141.155 194.695 ;
        RECT 141.845 194.320 142.545 194.390 ;
        RECT 143.395 194.320 144.095 194.390 ;
        RECT 141.845 194.090 142.805 194.320 ;
        RECT 143.135 194.090 144.095 194.320 ;
        RECT 141.565 192.835 141.795 193.930 ;
        RECT 141.530 191.335 141.830 192.835 ;
        RECT 141.565 185.930 141.795 191.335 ;
        RECT 142.855 189.090 143.085 193.930 ;
        RECT 144.145 192.835 144.375 193.930 ;
        RECT 144.110 191.335 144.410 192.835 ;
        RECT 142.820 187.590 143.120 189.090 ;
        RECT 142.855 185.930 143.085 187.590 ;
        RECT 144.145 185.930 144.375 191.335 ;
        RECT 141.845 185.540 142.805 185.770 ;
        RECT 143.135 185.540 144.095 185.770 ;
        RECT 144.785 185.165 145.185 194.695 ;
        RECT 145.875 194.320 146.575 194.390 ;
        RECT 147.425 194.320 148.125 194.390 ;
        RECT 145.875 194.090 146.835 194.320 ;
        RECT 147.165 194.090 148.125 194.320 ;
        RECT 145.595 192.835 145.825 193.930 ;
        RECT 145.560 191.335 145.860 192.835 ;
        RECT 145.595 185.930 145.825 191.335 ;
        RECT 146.885 189.090 147.115 193.930 ;
        RECT 148.175 192.835 148.405 193.930 ;
        RECT 148.140 191.335 148.440 192.835 ;
        RECT 146.850 187.590 147.150 189.090 ;
        RECT 146.885 185.930 147.115 187.590 ;
        RECT 148.175 185.930 148.405 191.335 ;
        RECT 145.875 185.540 146.835 185.770 ;
        RECT 147.165 185.540 148.125 185.770 ;
        RECT 148.815 185.165 149.215 194.695 ;
        RECT 149.905 194.320 150.605 194.390 ;
        RECT 151.455 194.320 152.155 194.390 ;
        RECT 149.905 194.090 150.865 194.320 ;
        RECT 151.195 194.090 152.155 194.320 ;
        RECT 149.625 192.835 149.855 193.930 ;
        RECT 149.590 191.335 149.890 192.835 ;
        RECT 149.625 185.930 149.855 191.335 ;
        RECT 150.915 189.090 151.145 193.930 ;
        RECT 152.205 192.835 152.435 193.930 ;
        RECT 152.170 191.335 152.470 192.835 ;
        RECT 150.880 187.590 151.180 189.090 ;
        RECT 150.915 185.930 151.145 187.590 ;
        RECT 152.205 185.930 152.435 191.335 ;
        RECT 152.845 187.965 153.245 194.695 ;
        RECT 189.690 195.130 190.290 195.270 ;
        RECT 180.400 194.590 180.720 194.650 ;
        RECT 189.690 194.590 189.830 195.130 ;
        RECT 190.520 195.070 190.840 195.330 ;
        RECT 190.980 195.070 191.300 195.330 ;
        RECT 190.610 194.635 190.750 195.070 ;
        RECT 191.530 194.635 191.670 195.470 ;
        RECT 192.360 194.930 192.680 194.990 ;
        RECT 192.360 194.790 195.810 194.930 ;
        RECT 192.360 194.730 192.680 194.790 ;
        RECT 180.400 194.450 189.830 194.590 ;
        RECT 190.375 194.450 190.750 194.635 ;
        RECT 191.455 194.590 191.745 194.635 ;
        RECT 195.120 194.590 195.440 194.650 ;
        RECT 195.670 194.635 195.810 194.790 ;
        RECT 191.455 194.450 195.440 194.590 ;
        RECT 180.400 194.390 180.720 194.450 ;
        RECT 190.375 194.405 190.665 194.450 ;
        RECT 191.455 194.405 191.745 194.450 ;
        RECT 195.120 194.390 195.440 194.450 ;
        RECT 195.595 194.405 195.885 194.635 ;
        RECT 179.940 194.250 180.260 194.310 ;
        RECT 207.540 194.250 207.860 194.310 ;
        RECT 179.940 194.110 207.860 194.250 ;
        RECT 179.940 194.050 180.260 194.110 ;
        RECT 207.540 194.050 207.860 194.110 ;
        RECT 176.720 193.910 177.040 193.970 ;
        RECT 194.660 193.910 194.980 193.970 ;
        RECT 176.720 193.770 194.980 193.910 ;
        RECT 176.720 193.710 177.040 193.770 ;
        RECT 194.660 193.710 194.980 193.770 ;
        RECT 196.040 193.710 196.360 193.970 ;
        RECT 165.150 193.090 239.990 193.570 ;
        RECT 178.115 192.890 178.405 192.935 ;
        RECT 178.560 192.890 178.880 192.950 ;
        RECT 178.115 192.750 178.880 192.890 ;
        RECT 178.115 192.705 178.405 192.750 ;
        RECT 178.560 192.690 178.880 192.750 ;
        RECT 186.855 192.890 187.145 192.935 ;
        RECT 190.520 192.890 190.840 192.950 ;
        RECT 186.855 192.750 190.840 192.890 ;
        RECT 186.855 192.705 187.145 192.750 ;
        RECT 190.520 192.690 190.840 192.750 ;
        RECT 199.260 192.690 199.580 192.950 ;
        RECT 190.060 192.550 190.380 192.610 ;
        RECT 180.950 192.410 190.380 192.550 ;
        RECT 175.340 192.010 175.660 192.270 ;
        RECT 175.800 192.210 176.120 192.270 ;
        RECT 177.195 192.210 177.485 192.255 ;
        RECT 175.800 192.070 177.485 192.210 ;
        RECT 175.800 192.010 176.120 192.070 ;
        RECT 177.195 192.025 177.485 192.070 ;
        RECT 178.560 192.210 178.880 192.270 ;
        RECT 180.950 192.255 181.090 192.410 ;
        RECT 179.035 192.210 179.325 192.255 ;
        RECT 180.875 192.210 181.165 192.255 ;
        RECT 178.560 192.070 179.325 192.210 ;
        RECT 178.560 192.010 178.880 192.070 ;
        RECT 179.035 192.025 179.325 192.070 ;
        RECT 179.570 192.070 181.165 192.210 ;
        RECT 171.200 191.870 171.520 191.930 ;
        RECT 179.570 191.870 179.710 192.070 ;
        RECT 180.875 192.025 181.165 192.070 ;
        RECT 182.240 192.210 182.560 192.270 ;
        RECT 184.540 192.255 184.860 192.270 ;
        RECT 183.635 192.210 183.925 192.255 ;
        RECT 182.240 192.070 183.925 192.210 ;
        RECT 182.240 192.010 182.560 192.070 ;
        RECT 183.635 192.025 183.925 192.070 ;
        RECT 184.375 192.025 184.860 192.255 ;
        RECT 184.540 192.010 184.860 192.025 ;
        RECT 185.000 192.010 185.320 192.270 ;
        RECT 188.310 192.255 188.450 192.410 ;
        RECT 190.060 192.350 190.380 192.410 ;
        RECT 191.440 192.550 191.760 192.610 ;
        RECT 200.640 192.550 200.960 192.610 ;
        RECT 191.440 192.410 193.055 192.550 ;
        RECT 191.440 192.350 191.760 192.410 ;
        RECT 185.475 192.025 185.765 192.255 ;
        RECT 185.960 192.025 186.250 192.255 ;
        RECT 188.235 192.025 188.525 192.255 ;
        RECT 190.980 192.210 191.300 192.270 ;
        RECT 192.360 192.210 192.680 192.270 ;
        RECT 192.915 192.255 193.055 192.410 ;
        RECT 193.830 192.410 200.960 192.550 ;
        RECT 193.830 192.255 193.970 192.410 ;
        RECT 200.640 192.350 200.960 192.410 ;
        RECT 194.660 192.255 194.980 192.270 ;
        RECT 190.150 192.070 192.680 192.210 ;
        RECT 171.200 191.730 179.710 191.870 ;
        RECT 171.200 191.670 171.520 191.730 ;
        RECT 179.940 191.670 180.260 191.930 ;
        RECT 180.400 191.670 180.720 191.930 ;
        RECT 183.175 191.870 183.465 191.915 ;
        RECT 185.550 191.870 185.690 192.025 ;
        RECT 183.175 191.730 185.690 191.870 ;
        RECT 183.175 191.685 183.465 191.730 ;
        RECT 168.900 191.530 169.220 191.590 ;
        RECT 181.780 191.530 182.100 191.590 ;
        RECT 186.035 191.530 186.175 192.025 ;
        RECT 190.150 191.870 190.290 192.070 ;
        RECT 190.980 192.010 191.300 192.070 ;
        RECT 192.360 192.010 192.680 192.070 ;
        RECT 192.840 192.025 193.130 192.255 ;
        RECT 193.755 192.025 194.045 192.255 ;
        RECT 194.215 192.025 194.505 192.255 ;
        RECT 194.660 192.025 194.990 192.255 ;
        RECT 200.195 192.210 200.485 192.255 ;
        RECT 195.670 192.070 200.485 192.210 ;
        RECT 168.900 191.390 181.550 191.530 ;
        RECT 168.900 191.330 169.220 191.390 ;
        RECT 173.040 191.190 173.360 191.250 ;
        RECT 174.435 191.190 174.725 191.235 ;
        RECT 173.040 191.050 174.725 191.190 ;
        RECT 173.040 190.990 173.360 191.050 ;
        RECT 174.435 191.005 174.725 191.050 ;
        RECT 176.260 190.990 176.580 191.250 ;
        RECT 181.410 191.235 181.550 191.390 ;
        RECT 181.780 191.390 186.175 191.530 ;
        RECT 188.310 191.730 190.290 191.870 ;
        RECT 190.535 191.870 190.825 191.915 ;
        RECT 194.290 191.870 194.430 192.025 ;
        RECT 194.660 192.010 194.980 192.025 ;
        RECT 190.535 191.730 194.430 191.870 ;
        RECT 181.780 191.330 182.100 191.390 ;
        RECT 181.335 191.005 181.625 191.235 ;
        RECT 182.240 191.190 182.560 191.250 ;
        RECT 188.310 191.190 188.450 191.730 ;
        RECT 190.535 191.685 190.825 191.730 ;
        RECT 195.670 191.575 195.810 192.070 ;
        RECT 200.195 192.025 200.485 192.070 ;
        RECT 196.040 191.870 196.360 191.930 ;
        RECT 201.575 191.870 201.865 191.915 ;
        RECT 196.040 191.730 210.070 191.870 ;
        RECT 196.040 191.670 196.360 191.730 ;
        RECT 201.575 191.685 201.865 191.730 ;
        RECT 195.595 191.345 195.885 191.575 ;
        RECT 209.930 191.250 210.070 191.730 ;
        RECT 182.240 191.050 188.450 191.190 ;
        RECT 182.240 190.990 182.560 191.050 ;
        RECT 188.680 190.990 189.000 191.250 ;
        RECT 201.115 191.190 201.405 191.235 ;
        RECT 204.320 191.190 204.640 191.250 ;
        RECT 201.115 191.050 204.640 191.190 ;
        RECT 201.115 191.005 201.405 191.050 ;
        RECT 204.320 190.990 204.640 191.050 ;
        RECT 209.840 190.990 210.160 191.250 ;
        RECT 165.150 190.370 239.210 190.850 ;
        RECT 169.820 190.170 170.140 190.230 ;
        RECT 176.260 190.170 176.580 190.230 ;
        RECT 169.820 190.030 173.730 190.170 ;
        RECT 169.820 189.970 170.140 190.030 ;
        RECT 166.600 188.950 166.920 189.210 ;
        RECT 171.675 189.150 171.965 189.195 ;
        RECT 172.580 189.150 172.900 189.210 ;
        RECT 171.675 189.010 172.900 189.150 ;
        RECT 171.675 188.965 171.965 189.010 ;
        RECT 172.580 188.950 172.900 189.010 ;
        RECT 173.055 188.965 173.345 189.195 ;
        RECT 173.130 188.810 173.270 188.965 ;
        RECT 171.750 188.670 173.270 188.810 ;
        RECT 173.590 188.810 173.730 190.030 ;
        RECT 174.050 190.030 176.580 190.170 ;
        RECT 174.050 189.195 174.190 190.030 ;
        RECT 176.260 189.970 176.580 190.030 ;
        RECT 180.400 189.970 180.720 190.230 ;
        RECT 184.555 190.170 184.845 190.215 ;
        RECT 188.680 190.170 189.000 190.230 ;
        RECT 184.555 190.030 189.000 190.170 ;
        RECT 184.555 189.985 184.845 190.030 ;
        RECT 188.680 189.970 189.000 190.030 ;
        RECT 190.535 189.985 190.825 190.215 ;
        RECT 208.475 190.170 208.765 190.215 ;
        RECT 208.920 190.170 209.240 190.230 ;
        RECT 208.475 190.030 209.240 190.170 ;
        RECT 208.475 189.985 208.765 190.030 ;
        RECT 180.490 189.490 180.630 189.970 ;
        RECT 182.240 189.830 182.560 189.890 ;
        RECT 190.610 189.830 190.750 189.985 ;
        RECT 208.920 189.970 209.240 190.030 ;
        RECT 226.415 190.170 226.705 190.215 ;
        RECT 226.860 190.170 227.180 190.230 ;
        RECT 226.415 190.030 227.180 190.170 ;
        RECT 226.415 189.985 226.705 190.030 ;
        RECT 226.860 189.970 227.180 190.030 ;
        RECT 182.240 189.690 190.750 189.830 ;
        RECT 191.070 189.690 196.755 189.830 ;
        RECT 182.240 189.630 182.560 189.690 ;
        RECT 180.875 189.490 181.165 189.535 ;
        RECT 191.070 189.490 191.210 189.690 ;
        RECT 180.490 189.350 181.165 189.490 ;
        RECT 180.875 189.305 181.165 189.350 ;
        RECT 183.250 189.350 191.210 189.490 ;
        RECT 192.375 189.490 192.665 189.535 ;
        RECT 192.375 189.350 196.270 189.490 ;
        RECT 173.975 188.965 174.265 189.195 ;
        RECT 174.880 189.150 175.200 189.210 ;
        RECT 175.355 189.150 175.645 189.195 ;
        RECT 174.880 189.010 175.645 189.150 ;
        RECT 174.880 188.950 175.200 189.010 ;
        RECT 175.355 188.965 175.645 189.010 ;
        RECT 176.735 189.150 177.025 189.195 ;
        RECT 179.020 189.150 179.340 189.210 ;
        RECT 176.735 189.010 179.340 189.150 ;
        RECT 176.735 188.965 177.025 189.010 ;
        RECT 179.020 188.950 179.340 189.010 ;
        RECT 179.495 188.965 179.785 189.195 ;
        RECT 178.575 188.810 178.865 188.855 ;
        RECT 173.590 188.670 178.865 188.810 ;
        RECT 171.750 188.530 171.890 188.670 ;
        RECT 178.575 188.625 178.865 188.670 ;
        RECT 167.535 188.470 167.825 188.515 ;
        RECT 170.280 188.470 170.600 188.530 ;
        RECT 167.535 188.330 170.600 188.470 ;
        RECT 167.535 188.285 167.825 188.330 ;
        RECT 170.280 188.270 170.600 188.330 ;
        RECT 171.660 188.270 171.980 188.530 ;
        RECT 172.595 188.470 172.885 188.515 ;
        RECT 173.500 188.470 173.820 188.530 ;
        RECT 172.595 188.330 173.820 188.470 ;
        RECT 172.595 188.285 172.885 188.330 ;
        RECT 173.500 188.270 173.820 188.330 ;
        RECT 176.275 188.470 176.565 188.515 ;
        RECT 176.720 188.470 177.040 188.530 ;
        RECT 176.275 188.330 177.040 188.470 ;
        RECT 176.275 188.285 176.565 188.330 ;
        RECT 176.720 188.270 177.040 188.330 ;
        RECT 177.640 188.270 177.960 188.530 ;
        RECT 178.100 188.470 178.420 188.530 ;
        RECT 179.570 188.470 179.710 188.965 ;
        RECT 180.400 188.950 180.720 189.210 ;
        RECT 181.320 189.150 181.640 189.210 ;
        RECT 182.715 189.150 183.005 189.195 ;
        RECT 181.320 189.010 183.005 189.150 ;
        RECT 181.320 188.950 181.640 189.010 ;
        RECT 182.715 188.965 183.005 189.010 ;
        RECT 183.250 188.810 183.390 189.350 ;
        RECT 192.375 189.305 192.665 189.350 ;
        RECT 183.635 189.150 183.925 189.195 ;
        RECT 185.000 189.150 185.320 189.210 ;
        RECT 183.635 189.010 185.320 189.150 ;
        RECT 183.635 188.965 183.925 189.010 ;
        RECT 185.000 188.950 185.320 189.010 ;
        RECT 185.460 188.950 185.780 189.210 ;
        RECT 187.300 188.950 187.620 189.210 ;
        RECT 189.600 188.950 189.920 189.210 ;
        RECT 190.060 188.950 190.380 189.210 ;
        RECT 191.440 188.950 191.760 189.210 ;
        RECT 191.900 189.150 192.220 189.210 ;
        RECT 192.795 189.150 193.085 189.195 ;
        RECT 191.900 189.010 193.085 189.150 ;
        RECT 191.900 188.950 192.220 189.010 ;
        RECT 192.795 188.965 193.085 189.010 ;
        RECT 193.280 189.150 193.600 189.210 ;
        RECT 196.130 189.195 196.270 189.350 ;
        RECT 196.615 189.195 196.755 189.690 ;
        RECT 197.435 189.645 197.725 189.875 ;
        RECT 225.940 189.830 226.260 189.890 ;
        RECT 235.140 189.830 235.460 189.890 ;
        RECT 225.940 189.690 235.460 189.830 ;
        RECT 197.510 189.490 197.650 189.645 ;
        RECT 225.940 189.630 226.260 189.690 ;
        RECT 235.140 189.630 235.460 189.690 ;
        RECT 209.840 189.490 210.160 189.550 ;
        RECT 226.860 189.490 227.180 189.550 ;
        RECT 232.840 189.490 233.160 189.550 ;
        RECT 197.510 189.350 209.610 189.490 ;
        RECT 194.215 189.150 194.505 189.195 ;
        RECT 193.280 189.010 194.505 189.150 ;
        RECT 193.280 188.950 193.600 189.010 ;
        RECT 194.215 188.965 194.505 189.010 ;
        RECT 194.680 188.965 194.970 189.195 ;
        RECT 196.055 188.965 196.345 189.195 ;
        RECT 196.540 188.965 196.830 189.195 ;
        RECT 197.420 189.150 197.740 189.210 ;
        RECT 209.470 189.195 209.610 189.350 ;
        RECT 209.840 189.350 210.990 189.490 ;
        RECT 209.840 189.290 210.160 189.350 ;
        RECT 198.815 189.150 199.105 189.195 ;
        RECT 197.420 189.010 199.105 189.150 ;
        RECT 180.490 188.670 183.390 188.810 ;
        RECT 185.920 188.810 186.240 188.870 ;
        RECT 191.530 188.810 191.670 188.950 ;
        RECT 194.755 188.810 194.895 188.965 ;
        RECT 197.420 188.950 197.740 189.010 ;
        RECT 198.815 188.965 199.105 189.010 ;
        RECT 209.395 188.965 209.685 189.195 ;
        RECT 210.300 188.950 210.620 189.210 ;
        RECT 210.850 189.195 210.990 189.350 ;
        RECT 226.860 189.350 231.230 189.490 ;
        RECT 226.860 189.290 227.180 189.350 ;
        RECT 210.775 189.150 211.065 189.195 ;
        RECT 210.775 189.010 222.030 189.150 ;
        RECT 210.775 188.965 211.065 189.010 ;
        RECT 195.120 188.810 195.440 188.870 ;
        RECT 185.920 188.670 188.910 188.810 ;
        RECT 191.530 188.670 195.440 188.810 ;
        RECT 180.490 188.530 180.630 188.670 ;
        RECT 185.920 188.610 186.240 188.670 ;
        RECT 178.100 188.330 179.710 188.470 ;
        RECT 178.100 188.270 178.420 188.330 ;
        RECT 180.400 188.270 180.720 188.530 ;
        RECT 181.780 188.270 182.100 188.530 ;
        RECT 186.380 188.270 186.700 188.530 ;
        RECT 188.220 188.270 188.540 188.530 ;
        RECT 188.770 188.515 188.910 188.670 ;
        RECT 195.120 188.610 195.440 188.670 ;
        RECT 195.580 188.610 195.900 188.870 ;
        RECT 221.890 188.530 222.030 189.010 ;
        RECT 227.320 188.950 227.640 189.210 ;
        RECT 228.255 188.965 228.545 189.195 ;
        RECT 228.700 189.150 229.020 189.210 ;
        RECT 230.540 189.150 230.860 189.210 ;
        RECT 231.090 189.195 231.230 189.350 ;
        RECT 231.550 189.350 233.160 189.490 ;
        RECT 231.550 189.195 231.690 189.350 ;
        RECT 232.840 189.290 233.160 189.350 ;
        RECT 228.700 189.010 230.860 189.150 ;
        RECT 226.400 188.810 226.720 188.870 ;
        RECT 227.780 188.810 228.100 188.870 ;
        RECT 226.400 188.670 228.100 188.810 ;
        RECT 228.330 188.810 228.470 188.965 ;
        RECT 228.700 188.950 229.020 189.010 ;
        RECT 230.540 188.950 230.860 189.010 ;
        RECT 231.015 188.965 231.305 189.195 ;
        RECT 231.475 188.965 231.765 189.195 ;
        RECT 231.920 189.150 232.240 189.210 ;
        RECT 233.775 189.150 234.065 189.195 ;
        RECT 231.920 189.010 234.065 189.150 ;
        RECT 231.920 188.950 232.240 189.010 ;
        RECT 233.775 188.965 234.065 189.010 ;
        RECT 229.160 188.810 229.480 188.870 ;
        RECT 228.330 188.670 229.480 188.810 ;
        RECT 226.400 188.610 226.720 188.670 ;
        RECT 227.780 188.610 228.100 188.670 ;
        RECT 229.160 188.610 229.480 188.670 ;
        RECT 188.695 188.285 188.985 188.515 ;
        RECT 190.980 188.470 191.300 188.530 ;
        RECT 193.280 188.470 193.600 188.530 ;
        RECT 190.980 188.330 193.600 188.470 ;
        RECT 190.980 188.270 191.300 188.330 ;
        RECT 193.280 188.270 193.600 188.330 ;
        RECT 193.740 188.270 194.060 188.530 ;
        RECT 197.895 188.470 198.185 188.515 ;
        RECT 199.720 188.470 200.040 188.530 ;
        RECT 197.895 188.330 200.040 188.470 ;
        RECT 197.895 188.285 198.185 188.330 ;
        RECT 199.720 188.270 200.040 188.330 ;
        RECT 221.800 188.470 222.120 188.530 ;
        RECT 228.700 188.470 229.020 188.530 ;
        RECT 221.800 188.330 229.020 188.470 ;
        RECT 221.800 188.270 222.120 188.330 ;
        RECT 228.700 188.270 229.020 188.330 ;
        RECT 230.080 188.270 230.400 188.530 ;
        RECT 231.460 188.470 231.780 188.530 ;
        RECT 232.395 188.470 232.685 188.515 ;
        RECT 231.460 188.330 232.685 188.470 ;
        RECT 231.460 188.270 231.780 188.330 ;
        RECT 232.395 188.285 232.685 188.330 ;
        RECT 232.855 188.470 233.145 188.515 ;
        RECT 233.300 188.470 233.620 188.530 ;
        RECT 232.855 188.330 233.620 188.470 ;
        RECT 232.855 188.285 233.145 188.330 ;
        RECT 233.300 188.270 233.620 188.330 ;
        RECT 149.905 185.540 150.865 185.770 ;
        RECT 151.195 185.540 152.155 185.770 ;
        RECT 152.845 185.165 155.165 187.965 ;
        RECT 165.150 187.650 239.990 188.130 ;
        RECT 170.740 187.250 171.060 187.510 ;
        RECT 172.135 187.450 172.425 187.495 ;
        RECT 179.020 187.450 179.340 187.510 ;
        RECT 180.860 187.450 181.180 187.510 ;
        RECT 172.135 187.310 175.570 187.450 ;
        RECT 172.135 187.265 172.425 187.310 ;
        RECT 174.880 187.110 175.200 187.170 ;
        RECT 171.290 186.970 175.200 187.110 ;
        RECT 168.455 186.585 168.745 186.815 ;
        RECT 168.530 186.430 168.670 186.585 ;
        RECT 169.820 186.570 170.140 186.830 ;
        RECT 170.280 186.770 170.600 186.830 ;
        RECT 171.290 186.815 171.430 186.970 ;
        RECT 174.880 186.910 175.200 186.970 ;
        RECT 171.215 186.770 171.505 186.815 ;
        RECT 170.280 186.630 171.505 186.770 ;
        RECT 170.280 186.570 170.600 186.630 ;
        RECT 171.215 186.585 171.505 186.630 ;
        RECT 171.660 186.770 171.980 186.830 ;
        RECT 173.055 186.770 173.345 186.815 ;
        RECT 171.660 186.630 173.345 186.770 ;
        RECT 171.660 186.570 171.980 186.630 ;
        RECT 173.055 186.585 173.345 186.630 ;
        RECT 173.960 186.570 174.280 186.830 ;
        RECT 170.740 186.430 171.060 186.490 ;
        RECT 168.530 186.290 171.060 186.430 ;
        RECT 174.970 186.430 175.110 186.910 ;
        RECT 175.430 186.830 175.570 187.310 ;
        RECT 175.890 187.310 179.340 187.450 ;
        RECT 175.340 186.570 175.660 186.830 ;
        RECT 175.890 186.430 176.030 187.310 ;
        RECT 179.020 187.250 179.340 187.310 ;
        RECT 180.490 187.310 181.180 187.450 ;
        RECT 176.275 187.110 176.565 187.155 ;
        RECT 180.490 187.110 180.630 187.310 ;
        RECT 180.860 187.250 181.180 187.310 ;
        RECT 182.240 187.250 182.560 187.510 ;
        RECT 183.620 187.250 183.940 187.510 ;
        RECT 184.630 187.310 190.290 187.450 ;
        RECT 184.630 187.170 184.770 187.310 ;
        RECT 184.540 187.110 184.860 187.170 ;
        RECT 187.300 187.110 187.620 187.170 ;
        RECT 176.275 186.970 180.630 187.110 ;
        RECT 180.950 186.970 184.860 187.110 ;
        RECT 176.275 186.925 176.565 186.970 ;
        RECT 180.950 186.830 181.090 186.970 ;
        RECT 184.540 186.910 184.860 186.970 ;
        RECT 185.550 186.970 187.620 187.110 ;
        RECT 176.720 186.570 177.040 186.830 ;
        RECT 177.655 186.585 177.945 186.815 ;
        RECT 176.260 186.430 176.580 186.490 ;
        RECT 174.970 186.290 176.580 186.430 ;
        RECT 170.740 186.230 171.060 186.290 ;
        RECT 176.260 186.230 176.580 186.290 ;
        RECT 167.520 186.090 167.840 186.150 ;
        RECT 177.730 186.090 177.870 186.585 ;
        RECT 179.020 186.570 179.340 186.830 ;
        RECT 179.940 186.570 180.260 186.830 ;
        RECT 180.860 186.570 181.180 186.830 ;
        RECT 181.335 186.770 181.625 186.815 ;
        RECT 182.240 186.770 182.560 186.830 ;
        RECT 185.550 186.815 185.690 186.970 ;
        RECT 187.300 186.910 187.620 186.970 ;
        RECT 187.760 187.110 188.080 187.170 ;
        RECT 189.140 187.110 189.460 187.170 ;
        RECT 187.760 186.970 189.460 187.110 ;
        RECT 190.150 187.110 190.290 187.310 ;
        RECT 190.520 187.250 190.840 187.510 ;
        RECT 191.900 187.450 192.220 187.510 ;
        RECT 195.595 187.450 195.885 187.495 ;
        RECT 196.500 187.450 196.820 187.510 ;
        RECT 191.900 187.310 194.430 187.450 ;
        RECT 191.900 187.250 192.220 187.310 ;
        RECT 191.440 187.110 191.760 187.170 ;
        RECT 194.290 187.155 194.430 187.310 ;
        RECT 195.595 187.310 196.820 187.450 ;
        RECT 195.595 187.265 195.885 187.310 ;
        RECT 196.500 187.250 196.820 187.310 ;
        RECT 200.275 187.310 202.710 187.450 ;
        RECT 190.150 186.970 193.055 187.110 ;
        RECT 187.760 186.910 188.080 186.970 ;
        RECT 189.140 186.910 189.460 186.970 ;
        RECT 191.440 186.910 191.760 186.970 ;
        RECT 181.335 186.630 182.560 186.770 ;
        RECT 181.335 186.585 181.625 186.630 ;
        RECT 182.240 186.570 182.560 186.630 ;
        RECT 182.715 186.585 183.005 186.815 ;
        RECT 185.015 186.585 185.305 186.815 ;
        RECT 185.475 186.585 185.765 186.815 ;
        RECT 186.855 186.770 187.145 186.815 ;
        RECT 188.235 186.770 188.525 186.815 ;
        RECT 190.060 186.770 190.380 186.830 ;
        RECT 186.855 186.630 187.990 186.770 ;
        RECT 186.855 186.585 187.145 186.630 ;
        RECT 167.520 185.950 177.870 186.090 ;
        RECT 180.400 186.090 180.720 186.150 ;
        RECT 182.790 186.090 182.930 186.585 ;
        RECT 185.090 186.090 185.230 186.585 ;
        RECT 186.380 186.230 186.700 186.490 ;
        RECT 187.850 186.430 187.990 186.630 ;
        RECT 188.235 186.630 190.380 186.770 ;
        RECT 188.235 186.585 188.525 186.630 ;
        RECT 190.060 186.570 190.380 186.630 ;
        RECT 190.980 186.770 191.300 186.830 ;
        RECT 192.915 186.815 193.055 186.970 ;
        RECT 194.215 186.925 194.505 187.155 ;
        RECT 195.120 187.110 195.440 187.170 ;
        RECT 200.275 187.110 200.415 187.310 ;
        RECT 201.575 187.110 201.865 187.155 ;
        RECT 195.120 186.970 200.415 187.110 ;
        RECT 195.120 186.910 195.440 186.970 ;
        RECT 192.375 186.770 192.665 186.815 ;
        RECT 190.980 186.630 192.665 186.770 ;
        RECT 190.980 186.570 191.300 186.630 ;
        RECT 192.375 186.585 192.665 186.630 ;
        RECT 192.840 186.585 193.130 186.815 ;
        RECT 193.740 186.570 194.060 186.830 ;
        RECT 196.590 186.815 196.730 186.970 ;
        RECT 194.700 186.770 194.990 186.815 ;
        RECT 194.290 186.630 194.990 186.770 ;
        RECT 189.600 186.430 189.920 186.490 ;
        RECT 187.850 186.290 189.920 186.430 ;
        RECT 189.600 186.230 189.920 186.290 ;
        RECT 190.520 186.430 190.840 186.490 ;
        RECT 194.290 186.430 194.430 186.630 ;
        RECT 194.700 186.585 194.990 186.630 ;
        RECT 196.055 186.585 196.345 186.815 ;
        RECT 196.520 186.585 196.810 186.815 ;
        RECT 196.130 186.430 196.270 186.585 ;
        RECT 197.420 186.570 197.740 186.830 ;
        RECT 197.880 186.570 198.200 186.830 ;
        RECT 198.340 186.815 198.660 186.830 ;
        RECT 200.275 186.815 200.415 186.970 ;
        RECT 200.730 186.970 201.865 187.110 ;
        RECT 198.340 186.585 198.670 186.815 ;
        RECT 199.735 186.585 200.025 186.815 ;
        RECT 200.200 186.585 200.490 186.815 ;
        RECT 198.340 186.570 198.660 186.585 ;
        RECT 199.810 186.430 199.950 186.585 ;
        RECT 190.520 186.290 194.430 186.430 ;
        RECT 195.210 186.290 199.950 186.430 ;
        RECT 190.520 186.230 190.840 186.290 ;
        RECT 180.400 185.950 182.930 186.090 ;
        RECT 183.710 185.950 185.230 186.090 ;
        RECT 186.470 186.090 186.610 186.230 ;
        RECT 187.775 186.090 188.065 186.135 ;
        RECT 193.280 186.090 193.600 186.150 ;
        RECT 195.210 186.090 195.350 186.290 ;
        RECT 198.800 186.090 199.120 186.150 ;
        RECT 186.470 185.950 187.070 186.090 ;
        RECT 167.520 185.890 167.840 185.950 ;
        RECT 180.400 185.890 180.720 185.950 ;
        RECT 169.375 185.750 169.665 185.795 ;
        RECT 169.820 185.750 170.140 185.810 ;
        RECT 169.375 185.610 170.140 185.750 ;
        RECT 169.375 185.565 169.665 185.610 ;
        RECT 169.820 185.550 170.140 185.610 ;
        RECT 170.740 185.750 171.060 185.810 ;
        RECT 176.720 185.750 177.040 185.810 ;
        RECT 182.700 185.750 183.020 185.810 ;
        RECT 170.740 185.610 183.020 185.750 ;
        RECT 170.740 185.550 171.060 185.610 ;
        RECT 176.720 185.550 177.040 185.610 ;
        RECT 182.700 185.550 183.020 185.610 ;
        RECT 183.160 185.750 183.480 185.810 ;
        RECT 183.710 185.750 183.850 185.950 ;
        RECT 183.160 185.610 183.850 185.750 ;
        RECT 184.095 185.750 184.385 185.795 ;
        RECT 184.540 185.750 184.860 185.810 ;
        RECT 184.095 185.610 184.860 185.750 ;
        RECT 183.160 185.550 183.480 185.610 ;
        RECT 184.095 185.565 184.385 185.610 ;
        RECT 184.540 185.550 184.860 185.610 ;
        RECT 186.380 185.550 186.700 185.810 ;
        RECT 186.930 185.750 187.070 185.950 ;
        RECT 187.775 185.950 192.130 186.090 ;
        RECT 187.775 185.905 188.065 185.950 ;
        RECT 188.695 185.750 188.985 185.795 ;
        RECT 186.930 185.610 188.985 185.750 ;
        RECT 191.990 185.750 192.130 185.950 ;
        RECT 193.280 185.950 195.350 186.090 ;
        RECT 197.970 185.950 199.120 186.090 ;
        RECT 193.280 185.890 193.600 185.950 ;
        RECT 197.970 185.750 198.110 185.950 ;
        RECT 198.800 185.890 199.120 185.950 ;
        RECT 199.260 185.890 199.580 186.150 ;
        RECT 200.180 186.090 200.500 186.150 ;
        RECT 200.730 186.090 200.870 186.970 ;
        RECT 201.575 186.925 201.865 186.970 ;
        RECT 202.020 186.815 202.340 186.830 ;
        RECT 201.115 186.585 201.405 186.815 ;
        RECT 202.020 186.585 202.350 186.815 ;
        RECT 200.180 185.950 200.870 186.090 ;
        RECT 200.180 185.890 200.500 185.950 ;
        RECT 191.990 185.610 198.110 185.750 ;
        RECT 198.340 185.750 198.660 185.810 ;
        RECT 201.190 185.750 201.330 186.585 ;
        RECT 202.020 186.570 202.340 186.585 ;
        RECT 202.570 186.090 202.710 187.310 ;
        RECT 202.955 187.265 203.245 187.495 ;
        RECT 211.695 187.450 211.985 187.495 ;
        RECT 216.740 187.450 217.060 187.510 ;
        RECT 211.695 187.310 217.060 187.450 ;
        RECT 211.695 187.265 211.985 187.310 ;
        RECT 203.030 187.110 203.170 187.265 ;
        RECT 216.740 187.250 217.060 187.310 ;
        RECT 217.200 187.250 217.520 187.510 ;
        RECT 219.040 187.450 219.360 187.510 ;
        RECT 221.355 187.450 221.645 187.495 ;
        RECT 219.040 187.310 221.645 187.450 ;
        RECT 219.040 187.250 219.360 187.310 ;
        RECT 221.355 187.265 221.645 187.310 ;
        RECT 225.020 187.450 225.340 187.510 ;
        RECT 234.695 187.450 234.985 187.495 ;
        RECT 236.060 187.450 236.380 187.510 ;
        RECT 225.020 187.310 231.230 187.450 ;
        RECT 225.020 187.250 225.340 187.310 ;
        RECT 224.120 187.110 224.410 187.155 ;
        RECT 229.640 187.110 229.930 187.155 ;
        RECT 230.560 187.110 230.850 187.155 ;
        RECT 203.030 186.970 218.350 187.110 ;
        RECT 208.935 186.770 209.225 186.815 ;
        RECT 209.840 186.770 210.160 186.830 ;
        RECT 210.775 186.770 211.065 186.815 ;
        RECT 208.935 186.630 209.335 186.770 ;
        RECT 209.840 186.630 211.065 186.770 ;
        RECT 208.935 186.585 209.225 186.630 ;
        RECT 208.000 186.430 208.320 186.490 ;
        RECT 209.010 186.430 209.150 186.585 ;
        RECT 209.840 186.570 210.160 186.630 ;
        RECT 210.775 186.585 211.065 186.630 ;
        RECT 212.140 186.570 212.460 186.830 ;
        RECT 213.520 186.570 213.840 186.830 ;
        RECT 214.900 186.570 215.220 186.830 ;
        RECT 218.210 186.815 218.350 186.970 ;
        RECT 224.120 186.970 230.850 187.110 ;
        RECT 231.090 187.110 231.230 187.310 ;
        RECT 234.695 187.310 236.380 187.450 ;
        RECT 234.695 187.265 234.985 187.310 ;
        RECT 236.060 187.250 236.380 187.310 ;
        RECT 236.535 187.265 236.825 187.495 ;
        RECT 236.610 187.110 236.750 187.265 ;
        RECT 231.090 186.970 236.750 187.110 ;
        RECT 224.120 186.925 224.410 186.970 ;
        RECT 229.640 186.925 229.930 186.970 ;
        RECT 230.560 186.925 230.850 186.970 ;
        RECT 218.135 186.585 218.425 186.815 ;
        RECT 219.960 186.570 220.280 186.830 ;
        RECT 221.800 186.570 222.120 186.830 ;
        RECT 222.260 186.570 222.580 186.830 ;
        RECT 225.040 186.770 225.330 186.815 ;
        RECT 226.880 186.770 227.170 186.815 ;
        RECT 225.040 186.630 227.170 186.770 ;
        RECT 225.040 186.585 225.330 186.630 ;
        RECT 226.880 186.585 227.170 186.630 ;
        RECT 227.320 186.570 227.640 186.830 ;
        RECT 227.780 186.815 228.100 186.830 ;
        RECT 227.780 186.585 228.315 186.815 ;
        RECT 227.780 186.570 228.100 186.585 ;
        RECT 228.700 186.570 229.020 186.830 ;
        RECT 229.225 186.770 229.515 186.815 ;
        RECT 231.065 186.770 231.355 186.815 ;
        RECT 229.225 186.630 231.355 186.770 ;
        RECT 229.225 186.585 229.515 186.630 ;
        RECT 231.065 186.585 231.355 186.630 ;
        RECT 231.920 186.570 232.240 186.830 ;
        RECT 232.380 186.570 232.700 186.830 ;
        RECT 233.775 186.585 234.065 186.815 ;
        RECT 213.060 186.430 213.380 186.490 ;
        RECT 208.000 186.290 213.380 186.430 ;
        RECT 208.000 186.230 208.320 186.290 ;
        RECT 213.060 186.230 213.380 186.290 ;
        RECT 219.515 186.430 219.805 186.475 ;
        RECT 221.890 186.430 222.030 186.570 ;
        RECT 219.515 186.290 222.030 186.430 ;
        RECT 219.515 186.245 219.805 186.290 ;
        RECT 222.720 186.230 223.040 186.490 ;
        RECT 223.180 186.430 223.500 186.490 ;
        RECT 223.655 186.430 223.945 186.475 ;
        RECT 232.010 186.430 232.150 186.570 ;
        RECT 233.850 186.430 233.990 186.585 ;
        RECT 236.060 186.570 236.380 186.830 ;
        RECT 237.440 186.570 237.760 186.830 ;
        RECT 223.180 186.290 223.945 186.430 ;
        RECT 223.180 186.230 223.500 186.290 ;
        RECT 223.655 186.245 223.945 186.290 ;
        RECT 225.110 186.290 226.630 186.430 ;
        RECT 232.010 186.290 233.990 186.430 ;
        RECT 209.840 186.090 210.160 186.150 ;
        RECT 202.570 185.950 210.160 186.090 ;
        RECT 209.840 185.890 210.160 185.950 ;
        RECT 214.455 186.090 214.745 186.135 ;
        RECT 217.200 186.090 217.520 186.150 ;
        RECT 214.455 185.950 217.520 186.090 ;
        RECT 214.455 185.905 214.745 185.950 ;
        RECT 217.200 185.890 217.520 185.950 ;
        RECT 219.055 186.090 219.345 186.135 ;
        RECT 225.110 186.090 225.250 186.290 ;
        RECT 219.055 185.950 225.250 186.090 ;
        RECT 219.055 185.905 219.345 185.950 ;
        RECT 225.955 185.905 226.245 186.135 ;
        RECT 198.340 185.610 201.330 185.750 ;
        RECT 213.075 185.750 213.365 185.795 ;
        RECT 214.900 185.750 215.220 185.810 ;
        RECT 213.075 185.610 215.220 185.750 ;
        RECT 188.695 185.565 188.985 185.610 ;
        RECT 198.340 185.550 198.660 185.610 ;
        RECT 213.075 185.565 213.365 185.610 ;
        RECT 214.900 185.550 215.220 185.610 ;
        RECT 215.820 185.550 216.140 185.810 ;
        RECT 219.500 185.750 219.820 185.810 ;
        RECT 220.895 185.750 221.185 185.795 ;
        RECT 219.500 185.610 221.185 185.750 ;
        RECT 219.500 185.550 219.820 185.610 ;
        RECT 220.895 185.565 221.185 185.610 ;
        RECT 223.640 185.750 223.960 185.810 ;
        RECT 226.030 185.750 226.170 185.905 ;
        RECT 223.640 185.610 226.170 185.750 ;
        RECT 226.490 185.750 226.630 186.290 ;
        RECT 226.915 186.090 227.205 186.135 ;
        RECT 230.145 186.090 230.435 186.135 ;
        RECT 226.915 185.950 230.435 186.090 ;
        RECT 226.915 185.905 227.205 185.950 ;
        RECT 230.145 185.905 230.435 185.950 ;
        RECT 234.220 186.090 234.540 186.150 ;
        RECT 235.155 186.090 235.445 186.135 ;
        RECT 234.220 185.950 235.445 186.090 ;
        RECT 234.220 185.890 234.540 185.950 ;
        RECT 235.155 185.905 235.445 185.950 ;
        RECT 231.935 185.750 232.225 185.795 ;
        RECT 226.490 185.610 232.225 185.750 ;
        RECT 223.640 185.550 223.960 185.610 ;
        RECT 231.935 185.565 232.225 185.610 ;
        RECT 232.380 185.750 232.700 185.810 ;
        RECT 232.855 185.750 233.145 185.795 ;
        RECT 232.380 185.610 233.145 185.750 ;
        RECT 232.380 185.550 232.700 185.610 ;
        RECT 232.855 185.565 233.145 185.610 ;
        RECT 108.515 184.765 155.165 185.165 ;
        RECT 165.150 184.930 239.210 185.410 ;
        RECT 167.520 184.530 167.840 184.790 ;
        RECT 170.280 184.530 170.600 184.790 ;
        RECT 172.120 184.730 172.440 184.790 ;
        RECT 178.100 184.730 178.420 184.790 ;
        RECT 172.120 184.590 173.730 184.730 ;
        RECT 172.120 184.530 172.440 184.590 ;
        RECT 168.915 184.205 169.205 184.435 ;
        RECT 170.370 184.390 170.510 184.530 ;
        RECT 170.370 184.250 173.270 184.390 ;
        RECT 168.990 184.050 169.130 184.205 ;
        RECT 168.990 183.910 171.890 184.050 ;
        RECT 166.600 183.510 166.920 183.770 ;
        RECT 167.980 183.510 168.300 183.770 ;
        RECT 169.375 183.525 169.665 183.755 ;
        RECT 169.450 183.370 169.590 183.525 ;
        RECT 170.740 183.510 171.060 183.770 ;
        RECT 171.750 183.755 171.890 183.910 ;
        RECT 173.130 183.755 173.270 184.250 ;
        RECT 173.590 184.050 173.730 184.590 ;
        RECT 174.510 184.590 178.420 184.730 ;
        RECT 173.960 184.190 174.280 184.450 ;
        RECT 174.510 184.435 174.650 184.590 ;
        RECT 178.100 184.530 178.420 184.590 ;
        RECT 178.560 184.530 178.880 184.790 ;
        RECT 183.620 184.730 183.940 184.790 ;
        RECT 188.695 184.730 188.985 184.775 ;
        RECT 183.620 184.590 188.985 184.730 ;
        RECT 183.620 184.530 183.940 184.590 ;
        RECT 188.695 184.545 188.985 184.590 ;
        RECT 191.440 184.530 191.760 184.790 ;
        RECT 194.675 184.730 194.965 184.775 ;
        RECT 195.580 184.730 195.900 184.790 ;
        RECT 194.675 184.590 195.900 184.730 ;
        RECT 194.675 184.545 194.965 184.590 ;
        RECT 195.580 184.530 195.900 184.590 ;
        RECT 197.880 184.530 198.200 184.790 ;
        RECT 207.540 184.530 207.860 184.790 ;
        RECT 214.900 184.730 215.220 184.790 ;
        RECT 219.515 184.730 219.805 184.775 ;
        RECT 222.720 184.730 223.040 184.790 ;
        RECT 208.090 184.590 213.750 184.730 ;
        RECT 174.435 184.205 174.725 184.435 ;
        RECT 180.860 184.390 181.180 184.450 ;
        RECT 177.265 184.250 181.180 184.390 ;
        RECT 173.590 183.910 176.950 184.050 ;
        RECT 175.340 183.755 175.660 183.770 ;
        RECT 171.675 183.525 171.965 183.755 ;
        RECT 173.055 183.525 173.345 183.755 ;
        RECT 175.330 183.525 175.660 183.755 ;
        RECT 175.340 183.510 175.660 183.525 ;
        RECT 175.800 183.510 176.120 183.770 ;
        RECT 172.580 183.370 172.900 183.430 ;
        RECT 169.450 183.230 172.900 183.370 ;
        RECT 172.580 183.170 172.900 183.230 ;
        RECT 176.275 183.185 176.565 183.415 ;
        RECT 176.810 183.370 176.950 183.910 ;
        RECT 177.265 183.755 177.405 184.250 ;
        RECT 180.860 184.190 181.180 184.250 ;
        RECT 184.080 184.190 184.400 184.450 ;
        RECT 185.475 184.390 185.765 184.435 ;
        RECT 185.475 184.250 190.290 184.390 ;
        RECT 185.475 184.205 185.765 184.250 ;
        RECT 177.190 183.525 177.480 183.755 ;
        RECT 177.655 183.525 177.945 183.755 ;
        RECT 178.100 183.710 178.420 183.770 ;
        RECT 179.470 183.710 179.760 183.755 ;
        RECT 178.100 183.570 179.760 183.710 ;
        RECT 177.730 183.370 177.870 183.525 ;
        RECT 178.100 183.510 178.420 183.570 ;
        RECT 179.470 183.525 179.760 183.570 ;
        RECT 179.940 183.510 180.260 183.770 ;
        RECT 180.860 183.755 181.180 183.770 ;
        RECT 180.860 183.525 181.345 183.755 ;
        RECT 181.795 183.525 182.085 183.755 ;
        RECT 180.860 183.510 181.180 183.525 ;
        RECT 176.810 183.230 180.170 183.370 ;
        RECT 170.280 182.830 170.600 183.090 ;
        RECT 176.350 183.030 176.490 183.185 ;
        RECT 178.560 183.030 178.880 183.090 ;
        RECT 176.350 182.890 178.880 183.030 ;
        RECT 180.030 183.030 180.170 183.230 ;
        RECT 180.400 183.170 180.720 183.430 ;
        RECT 181.870 183.370 182.010 183.525 ;
        RECT 182.240 183.510 182.560 183.770 ;
        RECT 183.175 183.525 183.465 183.755 ;
        RECT 184.170 183.710 184.310 184.190 ;
        RECT 187.760 184.050 188.080 184.110 ;
        RECT 185.090 183.910 188.080 184.050 ;
        RECT 190.150 184.050 190.290 184.250 ;
        RECT 190.520 184.190 190.840 184.450 ;
        RECT 193.295 184.390 193.585 184.435 ;
        RECT 197.970 184.390 198.110 184.530 ;
        RECT 193.295 184.250 198.110 184.390 ;
        RECT 193.295 184.205 193.585 184.250 ;
        RECT 192.360 184.050 192.680 184.110 ;
        RECT 196.500 184.050 196.820 184.110 ;
        RECT 190.150 183.910 192.130 184.050 ;
        RECT 184.555 183.710 184.845 183.755 ;
        RECT 184.170 183.570 184.845 183.710 ;
        RECT 184.555 183.525 184.845 183.570 ;
        RECT 180.950 183.230 182.010 183.370 ;
        RECT 183.250 183.370 183.390 183.525 ;
        RECT 185.090 183.370 185.230 183.910 ;
        RECT 187.760 183.850 188.080 183.910 ;
        RECT 186.855 183.525 187.145 183.755 ;
        RECT 188.235 183.710 188.525 183.755 ;
        RECT 190.060 183.710 190.380 183.770 ;
        RECT 190.995 183.710 191.285 183.755 ;
        RECT 188.235 183.570 191.285 183.710 ;
        RECT 191.990 183.710 192.130 183.910 ;
        RECT 192.360 183.910 196.820 184.050 ;
        RECT 192.360 183.850 192.680 183.910 ;
        RECT 196.500 183.850 196.820 183.910 ;
        RECT 197.435 183.865 197.725 184.095 ;
        RECT 203.860 184.050 204.180 184.110 ;
        RECT 198.890 183.910 204.180 184.050 ;
        RECT 195.120 183.710 195.440 183.770 ;
        RECT 191.990 183.570 195.440 183.710 ;
        RECT 188.235 183.525 188.525 183.570 ;
        RECT 183.250 183.230 185.230 183.370 ;
        RECT 186.930 183.370 187.070 183.525 ;
        RECT 190.060 183.510 190.380 183.570 ;
        RECT 190.995 183.525 191.285 183.570 ;
        RECT 195.120 183.510 195.440 183.570 ;
        RECT 196.960 183.710 197.280 183.770 ;
        RECT 197.510 183.710 197.650 183.865 ;
        RECT 196.960 183.570 197.650 183.710 ;
        RECT 196.960 183.510 197.280 183.570 ;
        RECT 191.900 183.370 192.220 183.430 ;
        RECT 186.930 183.230 192.220 183.370 ;
        RECT 180.950 183.030 181.090 183.230 ;
        RECT 191.900 183.170 192.220 183.230 ;
        RECT 196.500 183.170 196.820 183.430 ;
        RECT 197.510 183.370 197.650 183.570 ;
        RECT 198.890 183.370 199.030 183.910 ;
        RECT 203.860 183.850 204.180 183.910 ;
        RECT 200.180 183.710 200.500 183.770 ;
        RECT 202.955 183.710 203.245 183.755 ;
        RECT 200.180 183.570 203.245 183.710 ;
        RECT 200.180 183.510 200.500 183.570 ;
        RECT 202.955 183.525 203.245 183.570 ;
        RECT 203.400 183.710 203.720 183.770 ;
        RECT 204.335 183.710 204.625 183.755 ;
        RECT 203.400 183.570 204.625 183.710 ;
        RECT 203.400 183.510 203.720 183.570 ;
        RECT 204.335 183.525 204.625 183.570 ;
        RECT 206.160 183.510 206.480 183.770 ;
        RECT 197.510 183.230 199.030 183.370 ;
        RECT 199.260 183.170 199.580 183.430 ;
        RECT 208.090 183.370 208.230 184.590 ;
        RECT 213.610 184.450 213.750 184.590 ;
        RECT 214.070 184.590 214.670 184.730 ;
        RECT 209.345 184.390 209.635 184.435 ;
        RECT 212.575 184.390 212.865 184.435 ;
        RECT 209.345 184.250 212.865 184.390 ;
        RECT 209.345 184.205 209.635 184.250 ;
        RECT 212.575 184.205 212.865 184.250 ;
        RECT 213.520 184.190 213.840 184.450 ;
        RECT 209.840 184.050 210.160 184.110 ;
        RECT 210.775 184.050 211.065 184.095 ;
        RECT 209.840 183.910 211.065 184.050 ;
        RECT 209.840 183.850 210.160 183.910 ;
        RECT 210.775 183.865 211.065 183.910 ;
        RECT 212.155 184.050 212.445 184.095 ;
        RECT 214.070 184.050 214.210 184.590 ;
        RECT 214.530 184.450 214.670 184.590 ;
        RECT 214.900 184.590 216.970 184.730 ;
        RECT 214.900 184.530 215.220 184.590 ;
        RECT 214.440 184.190 214.760 184.450 ;
        RECT 216.830 184.095 216.970 184.590 ;
        RECT 219.515 184.590 223.040 184.730 ;
        RECT 219.515 184.545 219.805 184.590 ;
        RECT 222.720 184.530 223.040 184.590 ;
        RECT 229.175 184.730 229.465 184.775 ;
        RECT 232.380 184.730 232.700 184.790 ;
        RECT 229.175 184.590 232.700 184.730 ;
        RECT 229.175 184.545 229.465 184.590 ;
        RECT 232.380 184.530 232.700 184.590 ;
        RECT 218.580 184.390 218.900 184.450 ;
        RECT 222.260 184.390 222.580 184.450 ;
        RECT 218.580 184.250 222.580 184.390 ;
        RECT 218.580 184.190 218.900 184.250 ;
        RECT 222.260 184.190 222.580 184.250 ;
        RECT 224.155 184.390 224.445 184.435 ;
        RECT 227.385 184.390 227.675 184.435 ;
        RECT 224.155 184.250 227.675 184.390 ;
        RECT 224.155 184.205 224.445 184.250 ;
        RECT 227.385 184.205 227.675 184.250 ;
        RECT 231.015 184.390 231.305 184.435 ;
        RECT 231.920 184.390 232.240 184.450 ;
        RECT 231.015 184.250 232.240 184.390 ;
        RECT 231.015 184.205 231.305 184.250 ;
        RECT 231.920 184.190 232.240 184.250 ;
        RECT 232.855 184.205 233.145 184.435 ;
        RECT 212.155 183.910 214.210 184.050 ;
        RECT 214.990 183.910 216.510 184.050 ;
        RECT 212.155 183.865 212.445 183.910 ;
        RECT 214.990 183.770 215.130 183.910 ;
        RECT 211.680 183.755 212.000 183.770 ;
        RECT 208.425 183.710 208.715 183.755 ;
        RECT 210.265 183.710 210.555 183.755 ;
        RECT 208.425 183.570 210.555 183.710 ;
        RECT 208.425 183.525 208.715 183.570 ;
        RECT 210.265 183.525 210.555 183.570 ;
        RECT 211.570 183.525 212.000 183.755 ;
        RECT 212.610 183.710 212.900 183.755 ;
        RECT 214.450 183.710 214.740 183.755 ;
        RECT 212.610 183.570 214.740 183.710 ;
        RECT 212.610 183.525 212.900 183.570 ;
        RECT 214.450 183.525 214.740 183.570 ;
        RECT 211.680 183.510 212.000 183.525 ;
        RECT 214.900 183.510 215.220 183.770 ;
        RECT 215.820 183.510 216.140 183.770 ;
        RECT 216.370 183.710 216.510 183.910 ;
        RECT 216.755 183.865 217.045 184.095 ;
        RECT 221.340 184.050 221.660 184.110 ;
        RECT 217.290 183.910 218.810 184.050 ;
        RECT 217.290 183.710 217.430 183.910 ;
        RECT 216.370 183.570 217.430 183.710 ;
        RECT 218.120 183.510 218.440 183.770 ;
        RECT 218.670 183.755 218.810 183.910 ;
        RECT 220.050 183.910 221.660 184.050 ;
        RECT 220.050 183.755 220.190 183.910 ;
        RECT 221.340 183.850 221.660 183.910 ;
        RECT 223.195 184.050 223.485 184.095 ;
        RECT 223.640 184.050 223.960 184.110 ;
        RECT 223.195 183.910 223.960 184.050 ;
        RECT 223.195 183.865 223.485 183.910 ;
        RECT 223.640 183.850 223.960 183.910 ;
        RECT 224.560 183.850 224.880 184.110 ;
        RECT 225.265 184.050 225.555 184.095 ;
        RECT 232.930 184.050 233.070 184.205 ;
        RECT 234.220 184.190 234.540 184.450 ;
        RECT 225.265 183.910 233.070 184.050 ;
        RECT 225.265 183.865 225.555 183.910 ;
        RECT 218.595 183.525 218.885 183.755 ;
        RECT 219.975 183.525 220.265 183.755 ;
        RECT 220.895 183.710 221.185 183.755 ;
        RECT 220.510 183.570 221.185 183.710 ;
        RECT 199.810 183.230 208.230 183.370 ;
        RECT 208.930 183.370 209.220 183.415 ;
        RECT 209.850 183.370 210.140 183.415 ;
        RECT 215.370 183.370 215.660 183.415 ;
        RECT 220.510 183.370 220.650 183.570 ;
        RECT 220.895 183.525 221.185 183.570 ;
        RECT 222.280 183.710 222.570 183.755 ;
        RECT 224.120 183.710 224.410 183.755 ;
        RECT 222.280 183.570 224.410 183.710 ;
        RECT 222.280 183.525 222.570 183.570 ;
        RECT 224.120 183.525 224.410 183.570 ;
        RECT 225.940 183.510 226.260 183.770 ;
        RECT 226.465 183.710 226.755 183.755 ;
        RECT 228.305 183.710 228.595 183.755 ;
        RECT 226.465 183.570 228.595 183.710 ;
        RECT 226.465 183.525 226.755 183.570 ;
        RECT 228.305 183.525 228.595 183.570 ;
        RECT 230.095 183.525 230.385 183.755 ;
        RECT 208.930 183.230 215.660 183.370 ;
        RECT 180.030 182.890 181.090 183.030 ;
        RECT 183.160 183.030 183.480 183.090 ;
        RECT 187.300 183.030 187.620 183.090 ;
        RECT 183.160 182.890 187.620 183.030 ;
        RECT 178.560 182.830 178.880 182.890 ;
        RECT 183.160 182.830 183.480 182.890 ;
        RECT 187.300 182.830 187.620 182.890 ;
        RECT 187.775 183.030 188.065 183.075 ;
        RECT 190.980 183.030 191.300 183.090 ;
        RECT 187.775 182.890 191.300 183.030 ;
        RECT 187.775 182.845 188.065 182.890 ;
        RECT 190.980 182.830 191.300 182.890 ;
        RECT 191.440 183.030 191.760 183.090 ;
        RECT 196.975 183.030 197.265 183.075 ;
        RECT 191.440 182.890 197.265 183.030 ;
        RECT 191.440 182.830 191.760 182.890 ;
        RECT 196.975 182.845 197.265 182.890 ;
        RECT 197.880 183.030 198.200 183.090 ;
        RECT 199.810 183.075 199.950 183.230 ;
        RECT 208.930 183.185 209.220 183.230 ;
        RECT 209.850 183.185 210.140 183.230 ;
        RECT 215.370 183.185 215.660 183.230 ;
        RECT 215.910 183.230 220.650 183.370 ;
        RECT 221.360 183.370 221.650 183.415 ;
        RECT 226.880 183.370 227.170 183.415 ;
        RECT 227.800 183.370 228.090 183.415 ;
        RECT 221.360 183.230 228.090 183.370 ;
        RECT 199.735 183.030 200.025 183.075 ;
        RECT 197.880 182.890 200.025 183.030 ;
        RECT 197.880 182.830 198.200 182.890 ;
        RECT 199.735 182.845 200.025 182.890 ;
        RECT 200.180 183.030 200.500 183.090 ;
        RECT 202.035 183.030 202.325 183.075 ;
        RECT 200.180 182.890 202.325 183.030 ;
        RECT 200.180 182.830 200.500 182.890 ;
        RECT 202.035 182.845 202.325 182.890 ;
        RECT 205.255 183.030 205.545 183.075 ;
        RECT 206.620 183.030 206.940 183.090 ;
        RECT 205.255 182.890 206.940 183.030 ;
        RECT 205.255 182.845 205.545 182.890 ;
        RECT 206.620 182.830 206.940 182.890 ;
        RECT 207.095 183.030 207.385 183.075 ;
        RECT 215.910 183.030 216.050 183.230 ;
        RECT 221.360 183.185 221.650 183.230 ;
        RECT 226.880 183.185 227.170 183.230 ;
        RECT 227.800 183.185 228.090 183.230 ;
        RECT 207.095 182.890 216.050 183.030 ;
        RECT 216.280 183.030 216.600 183.090 ;
        RECT 217.215 183.030 217.505 183.075 ;
        RECT 216.280 182.890 217.505 183.030 ;
        RECT 207.095 182.845 207.385 182.890 ;
        RECT 216.280 182.830 216.600 182.890 ;
        RECT 217.215 182.845 217.505 182.890 ;
        RECT 217.660 183.030 217.980 183.090 ;
        RECT 219.960 183.030 220.280 183.090 ;
        RECT 217.660 182.890 220.280 183.030 ;
        RECT 217.660 182.830 217.980 182.890 ;
        RECT 219.960 182.830 220.280 182.890 ;
        RECT 224.560 183.030 224.880 183.090 ;
        RECT 230.170 183.030 230.310 183.525 ;
        RECT 232.380 183.510 232.700 183.770 ;
        RECT 233.775 183.710 234.065 183.755 ;
        RECT 234.680 183.710 235.000 183.770 ;
        RECT 233.775 183.570 235.000 183.710 ;
        RECT 233.775 183.525 234.065 183.570 ;
        RECT 234.680 183.510 235.000 183.570 ;
        RECT 235.140 183.510 235.460 183.770 ;
        RECT 236.535 183.710 236.825 183.755 ;
        RECT 237.900 183.710 238.220 183.770 ;
        RECT 236.535 183.570 238.220 183.710 ;
        RECT 236.535 183.525 236.825 183.570 ;
        RECT 237.900 183.510 238.220 183.570 ;
        RECT 224.560 182.890 230.310 183.030 ;
        RECT 231.475 183.030 231.765 183.075 ;
        RECT 232.380 183.030 232.700 183.090 ;
        RECT 231.475 182.890 232.700 183.030 ;
        RECT 224.560 182.830 224.880 182.890 ;
        RECT 231.475 182.845 231.765 182.890 ;
        RECT 232.380 182.830 232.700 182.890 ;
        RECT 235.600 182.830 235.920 183.090 ;
        RECT 63.895 181.400 64.595 182.400 ;
        RECT 77.595 182.370 78.595 182.605 ;
        RECT 77.595 181.195 78.595 181.430 ;
        RECT 80.185 181.400 81.755 182.400 ;
        RECT 83.345 182.370 84.345 182.605 ;
        RECT 83.345 181.195 84.345 181.430 ;
        RECT 97.345 181.400 98.045 182.400 ;
        RECT 64.175 180.965 80.135 181.195 ;
        RECT 81.805 180.965 97.765 181.195 ;
        RECT 77.595 180.730 78.595 180.965 ;
        RECT 83.345 180.730 84.345 180.965 ;
        RECT 98.485 180.110 155.900 182.710 ;
        RECT 165.150 182.210 239.990 182.690 ;
        RECT 168.900 182.010 169.220 182.070 ;
        RECT 169.375 182.010 169.665 182.055 ;
        RECT 168.900 181.870 169.665 182.010 ;
        RECT 168.900 181.810 169.220 181.870 ;
        RECT 169.375 181.825 169.665 181.870 ;
        RECT 174.895 182.010 175.185 182.055 ;
        RECT 178.100 182.010 178.420 182.070 ;
        RECT 174.895 181.870 178.420 182.010 ;
        RECT 174.895 181.825 175.185 181.870 ;
        RECT 178.100 181.810 178.420 181.870 ;
        RECT 179.035 182.010 179.325 182.055 ;
        RECT 179.940 182.010 180.260 182.070 ;
        RECT 179.035 181.870 180.260 182.010 ;
        RECT 179.035 181.825 179.325 181.870 ;
        RECT 179.940 181.810 180.260 181.870 ;
        RECT 180.400 182.010 180.720 182.070 ;
        RECT 182.715 182.010 183.005 182.055 ;
        RECT 180.400 181.870 183.005 182.010 ;
        RECT 180.400 181.810 180.720 181.870 ;
        RECT 182.715 181.825 183.005 181.870 ;
        RECT 184.555 182.010 184.845 182.055 ;
        RECT 185.920 182.010 186.240 182.070 ;
        RECT 184.555 181.870 186.240 182.010 ;
        RECT 184.555 181.825 184.845 181.870 ;
        RECT 185.920 181.810 186.240 181.870 ;
        RECT 186.380 181.810 186.700 182.070 ;
        RECT 186.855 182.010 187.145 182.055 ;
        RECT 189.140 182.010 189.460 182.070 ;
        RECT 186.855 181.870 189.460 182.010 ;
        RECT 186.855 181.825 187.145 181.870 ;
        RECT 189.140 181.810 189.460 181.870 ;
        RECT 194.215 182.010 194.505 182.055 ;
        RECT 194.660 182.010 194.980 182.070 ;
        RECT 194.215 181.870 194.980 182.010 ;
        RECT 194.215 181.825 194.505 181.870 ;
        RECT 194.660 181.810 194.980 181.870 ;
        RECT 196.055 181.825 196.345 182.055 ;
        RECT 196.515 182.010 196.805 182.055 ;
        RECT 197.420 182.010 197.740 182.070 ;
        RECT 196.515 181.870 197.740 182.010 ;
        RECT 196.515 181.825 196.805 181.870 ;
        RECT 176.720 181.670 177.040 181.730 ;
        RECT 184.080 181.670 184.400 181.730 ;
        RECT 185.000 181.670 185.320 181.730 ;
        RECT 170.370 181.530 176.490 181.670 ;
        RECT 170.370 181.390 170.510 181.530 ;
        RECT 167.060 181.130 167.380 181.390 ;
        RECT 168.455 181.330 168.745 181.375 ;
        RECT 169.360 181.330 169.680 181.390 ;
        RECT 168.455 181.190 169.680 181.330 ;
        RECT 168.455 181.145 168.745 181.190 ;
        RECT 169.360 181.130 169.680 181.190 ;
        RECT 170.280 181.130 170.600 181.390 ;
        RECT 170.740 181.330 171.060 181.390 ;
        RECT 171.660 181.330 171.980 181.390 ;
        RECT 170.740 181.190 171.980 181.330 ;
        RECT 170.740 181.130 171.060 181.190 ;
        RECT 171.660 181.130 171.980 181.190 ;
        RECT 172.595 181.330 172.885 181.375 ;
        RECT 173.500 181.330 173.820 181.390 ;
        RECT 172.595 181.190 173.820 181.330 ;
        RECT 172.595 181.145 172.885 181.190 ;
        RECT 173.500 181.130 173.820 181.190 ;
        RECT 173.960 181.130 174.280 181.390 ;
        RECT 176.350 181.375 176.490 181.530 ;
        RECT 176.720 181.530 177.405 181.670 ;
        RECT 176.720 181.470 177.040 181.530 ;
        RECT 175.355 181.330 175.645 181.375 ;
        RECT 175.355 181.190 176.030 181.330 ;
        RECT 175.355 181.145 175.645 181.190 ;
        RECT 172.580 180.650 172.900 180.710 ;
        RECT 173.960 180.650 174.280 180.710 ;
        RECT 172.580 180.510 174.280 180.650 ;
        RECT 175.890 180.650 176.030 181.190 ;
        RECT 176.275 181.145 176.565 181.375 ;
        RECT 177.265 181.350 177.405 181.530 ;
        RECT 184.080 181.530 185.320 181.670 ;
        RECT 186.470 181.670 186.610 181.810 ;
        RECT 188.695 181.670 188.985 181.715 ;
        RECT 186.470 181.530 188.985 181.670 ;
        RECT 184.080 181.470 184.400 181.530 ;
        RECT 185.000 181.470 185.320 181.530 ;
        RECT 188.695 181.485 188.985 181.530 ;
        RECT 193.740 181.470 194.060 181.730 ;
        RECT 196.130 181.670 196.270 181.825 ;
        RECT 197.420 181.810 197.740 181.870 ;
        RECT 198.340 181.810 198.660 182.070 ;
        RECT 198.815 182.010 199.105 182.055 ;
        RECT 200.180 182.010 200.500 182.070 ;
        RECT 198.815 181.870 200.500 182.010 ;
        RECT 198.815 181.825 199.105 181.870 ;
        RECT 200.180 181.810 200.500 181.870 ;
        RECT 200.640 181.810 200.960 182.070 ;
        RECT 206.160 182.010 206.480 182.070 ;
        RECT 208.920 182.010 209.240 182.070 ;
        RECT 206.160 181.870 209.240 182.010 ;
        RECT 206.160 181.810 206.480 181.870 ;
        RECT 208.920 181.810 209.240 181.870 ;
        RECT 210.760 182.010 211.080 182.070 ;
        RECT 210.760 181.870 216.050 182.010 ;
        RECT 210.760 181.810 211.080 181.870 ;
        RECT 198.430 181.670 198.570 181.810 ;
        RECT 196.130 181.530 198.570 181.670 ;
        RECT 208.470 181.670 208.760 181.715 ;
        RECT 209.390 181.670 209.680 181.715 ;
        RECT 214.910 181.670 215.200 181.715 ;
        RECT 208.470 181.530 215.200 181.670 ;
        RECT 208.470 181.485 208.760 181.530 ;
        RECT 209.390 181.485 209.680 181.530 ;
        RECT 214.910 181.485 215.200 181.530 ;
        RECT 177.655 181.350 177.945 181.375 ;
        RECT 177.265 181.210 177.945 181.350 ;
        RECT 177.655 181.145 177.945 181.210 ;
        RECT 181.335 181.145 181.625 181.375 ;
        RECT 182.240 181.330 182.560 181.390 ;
        RECT 186.380 181.330 186.700 181.390 ;
        RECT 182.240 181.190 190.290 181.330 ;
        RECT 176.720 180.790 177.040 181.050 ;
        RECT 179.940 180.990 180.260 181.050 ;
        RECT 181.410 180.990 181.550 181.145 ;
        RECT 182.240 181.130 182.560 181.190 ;
        RECT 179.940 180.850 181.550 180.990 ;
        RECT 179.940 180.790 180.260 180.850 ;
        RECT 185.000 180.790 185.320 181.050 ;
        RECT 186.010 181.035 186.150 181.190 ;
        RECT 186.380 181.130 186.700 181.190 ;
        RECT 185.935 180.805 186.225 181.035 ;
        RECT 189.140 180.790 189.460 181.050 ;
        RECT 190.150 181.035 190.290 181.190 ;
        RECT 198.340 181.130 198.660 181.390 ;
        RECT 198.800 181.330 199.120 181.390 ;
        RECT 202.495 181.330 202.785 181.375 ;
        RECT 198.800 181.190 202.785 181.330 ;
        RECT 198.800 181.130 199.120 181.190 ;
        RECT 202.495 181.145 202.785 181.190 ;
        RECT 205.700 181.130 206.020 181.390 ;
        RECT 207.965 181.330 208.255 181.375 ;
        RECT 209.805 181.330 210.095 181.375 ;
        RECT 207.965 181.190 210.095 181.330 ;
        RECT 207.965 181.145 208.255 181.190 ;
        RECT 209.805 181.145 210.095 181.190 ;
        RECT 210.300 181.130 210.620 181.390 ;
        RECT 210.760 181.375 211.080 181.390 ;
        RECT 210.760 181.145 211.295 181.375 ;
        RECT 210.760 181.130 211.080 181.145 ;
        RECT 211.680 181.130 212.000 181.390 ;
        RECT 212.150 181.330 212.440 181.375 ;
        RECT 213.990 181.330 214.280 181.375 ;
        RECT 212.150 181.190 214.280 181.330 ;
        RECT 212.150 181.145 212.440 181.190 ;
        RECT 213.990 181.145 214.280 181.190 ;
        RECT 215.910 181.050 216.050 181.870 ;
        RECT 216.740 181.810 217.060 182.070 ;
        RECT 217.200 181.810 217.520 182.070 ;
        RECT 235.600 182.010 235.920 182.070 ;
        RECT 222.810 181.870 235.920 182.010 ;
        RECT 216.295 181.330 216.585 181.375 ;
        RECT 216.830 181.330 216.970 181.810 ;
        RECT 216.295 181.190 216.970 181.330 ;
        RECT 216.295 181.145 216.585 181.190 ;
        RECT 190.075 180.990 190.365 181.035 ;
        RECT 193.295 180.990 193.585 181.035 ;
        RECT 196.960 180.990 197.280 181.050 ;
        RECT 190.075 180.850 197.280 180.990 ;
        RECT 190.075 180.805 190.365 180.850 ;
        RECT 193.295 180.805 193.585 180.850 ;
        RECT 196.960 180.790 197.280 180.850 ;
        RECT 199.260 180.790 199.580 181.050 ;
        RECT 202.955 180.805 203.245 181.035 ;
        RECT 176.810 180.650 176.950 180.790 ;
        RECT 175.890 180.510 176.950 180.650 ;
        RECT 178.575 180.650 178.865 180.695 ;
        RECT 192.360 180.650 192.680 180.710 ;
        RECT 178.575 180.510 192.680 180.650 ;
        RECT 172.580 180.450 172.900 180.510 ;
        RECT 173.960 180.450 174.280 180.510 ;
        RECT 178.575 180.465 178.865 180.510 ;
        RECT 192.360 180.450 192.680 180.510 ;
        RECT 194.660 180.650 194.980 180.710 ;
        RECT 203.030 180.650 203.170 180.805 ;
        RECT 203.860 180.790 204.180 181.050 ;
        RECT 213.520 180.990 213.840 181.050 ;
        RECT 214.900 180.990 215.220 181.050 ;
        RECT 215.375 180.990 215.665 181.035 ;
        RECT 213.520 180.850 214.210 180.990 ;
        RECT 213.520 180.790 213.840 180.850 ;
        RECT 194.660 180.510 203.170 180.650 ;
        RECT 208.885 180.650 209.175 180.695 ;
        RECT 212.115 180.650 212.405 180.695 ;
        RECT 208.885 180.510 212.405 180.650 ;
        RECT 194.660 180.450 194.980 180.510 ;
        RECT 208.885 180.465 209.175 180.510 ;
        RECT 212.115 180.465 212.405 180.510 ;
        RECT 213.045 180.465 213.335 180.695 ;
        RECT 167.535 180.310 167.825 180.355 ;
        RECT 168.900 180.310 169.220 180.370 ;
        RECT 167.535 180.170 169.220 180.310 ;
        RECT 167.535 180.125 167.825 180.170 ;
        RECT 168.900 180.110 169.220 180.170 ;
        RECT 180.875 180.310 181.165 180.355 ;
        RECT 181.780 180.310 182.100 180.370 ;
        RECT 180.875 180.170 182.100 180.310 ;
        RECT 180.875 180.125 181.165 180.170 ;
        RECT 181.780 180.110 182.100 180.170 ;
        RECT 190.060 180.310 190.380 180.370 ;
        RECT 191.900 180.310 192.220 180.370 ;
        RECT 190.060 180.170 192.220 180.310 ;
        RECT 190.060 180.110 190.380 180.170 ;
        RECT 191.900 180.110 192.220 180.170 ;
        RECT 206.620 180.110 206.940 180.370 ;
        RECT 207.080 180.110 207.400 180.370 ;
        RECT 207.540 180.310 207.860 180.370 ;
        RECT 211.680 180.310 212.000 180.370 ;
        RECT 207.540 180.170 212.000 180.310 ;
        RECT 213.150 180.310 213.290 180.465 ;
        RECT 213.520 180.310 213.840 180.370 ;
        RECT 213.150 180.170 213.840 180.310 ;
        RECT 214.070 180.310 214.210 180.850 ;
        RECT 214.900 180.850 215.665 180.990 ;
        RECT 214.900 180.790 215.220 180.850 ;
        RECT 215.375 180.805 215.665 180.850 ;
        RECT 215.820 180.790 216.140 181.050 ;
        RECT 217.290 180.990 217.430 181.810 ;
        RECT 218.580 181.715 218.900 181.730 ;
        RECT 218.575 181.485 218.900 181.715 ;
        RECT 220.435 181.485 220.725 181.715 ;
        RECT 221.340 181.670 221.660 181.730 ;
        RECT 222.810 181.715 222.950 181.870 ;
        RECT 235.600 181.810 235.920 181.870 ;
        RECT 222.275 181.670 222.565 181.715 ;
        RECT 221.340 181.530 222.565 181.670 ;
        RECT 218.580 181.470 218.900 181.485 ;
        RECT 220.510 181.330 220.650 181.485 ;
        RECT 221.340 181.470 221.660 181.530 ;
        RECT 222.275 181.485 222.565 181.530 ;
        RECT 222.735 181.485 223.025 181.715 ;
        RECT 218.670 181.190 220.650 181.330 ;
        RECT 222.350 181.330 222.490 181.485 ;
        RECT 224.100 181.470 224.420 181.730 ;
        RECT 225.940 181.670 226.260 181.730 ;
        RECT 224.650 181.530 226.260 181.670 ;
        RECT 224.650 181.330 224.790 181.530 ;
        RECT 225.940 181.470 226.260 181.530 ;
        RECT 228.260 181.670 228.550 181.715 ;
        RECT 233.780 181.670 234.070 181.715 ;
        RECT 234.700 181.670 234.990 181.715 ;
        RECT 228.260 181.530 234.990 181.670 ;
        RECT 228.260 181.485 228.550 181.530 ;
        RECT 233.780 181.485 234.070 181.530 ;
        RECT 234.700 181.485 234.990 181.530 ;
        RECT 222.350 181.190 224.790 181.330 ;
        RECT 226.400 181.350 226.720 181.390 ;
        RECT 226.875 181.350 227.165 181.375 ;
        RECT 226.400 181.210 227.165 181.350 ;
        RECT 229.180 181.330 229.470 181.375 ;
        RECT 231.020 181.330 231.310 181.375 ;
        RECT 218.670 180.990 218.810 181.190 ;
        RECT 226.400 181.130 226.720 181.210 ;
        RECT 226.875 181.145 227.165 181.210 ;
        RECT 227.410 181.190 228.470 181.330 ;
        RECT 217.290 180.850 218.810 180.990 ;
        RECT 219.055 180.990 219.345 181.035 ;
        RECT 224.115 180.990 224.405 181.035 ;
        RECT 225.035 180.990 225.325 181.035 ;
        RECT 227.410 180.990 227.550 181.190 ;
        RECT 219.055 180.850 227.550 180.990 ;
        RECT 219.055 180.805 219.345 180.850 ;
        RECT 224.115 180.805 224.405 180.850 ;
        RECT 225.035 180.805 225.325 180.850 ;
        RECT 227.795 180.805 228.085 181.035 ;
        RECT 228.330 180.990 228.470 181.190 ;
        RECT 229.180 181.190 231.310 181.330 ;
        RECT 229.180 181.145 229.470 181.190 ;
        RECT 231.020 181.145 231.310 181.190 ;
        RECT 231.460 181.130 231.780 181.390 ;
        RECT 231.920 181.375 232.240 181.390 ;
        RECT 231.920 181.145 232.350 181.375 ;
        RECT 233.365 181.330 233.655 181.375 ;
        RECT 235.205 181.330 235.495 181.375 ;
        RECT 237.455 181.330 237.745 181.375 ;
        RECT 233.365 181.190 235.495 181.330 ;
        RECT 233.365 181.145 233.655 181.190 ;
        RECT 235.205 181.145 235.495 181.190 ;
        RECT 235.690 181.190 237.745 181.330 ;
        RECT 231.920 181.130 232.240 181.145 ;
        RECT 230.095 180.990 230.385 181.035 ;
        RECT 232.855 180.990 233.145 181.035 ;
        RECT 228.330 180.850 230.385 180.990 ;
        RECT 230.095 180.805 230.385 180.850 ;
        RECT 230.630 180.850 233.145 180.990 ;
        RECT 219.515 180.650 219.805 180.695 ;
        RECT 223.655 180.650 223.945 180.695 ;
        RECT 225.110 180.650 225.250 180.805 ;
        RECT 219.515 180.510 223.945 180.650 ;
        RECT 219.515 180.465 219.805 180.510 ;
        RECT 223.655 180.465 223.945 180.510 ;
        RECT 224.190 180.510 225.250 180.650 ;
        RECT 226.400 180.650 226.720 180.710 ;
        RECT 227.870 180.650 228.010 180.805 ;
        RECT 226.400 180.510 228.010 180.650 ;
        RECT 228.700 180.650 229.020 180.710 ;
        RECT 230.630 180.650 230.770 180.850 ;
        RECT 232.855 180.805 233.145 180.850 ;
        RECT 228.700 180.510 230.770 180.650 ;
        RECT 231.055 180.650 231.345 180.695 ;
        RECT 234.285 180.650 234.575 180.695 ;
        RECT 231.055 180.510 234.575 180.650 ;
        RECT 224.190 180.370 224.330 180.510 ;
        RECT 226.400 180.450 226.720 180.510 ;
        RECT 228.700 180.450 229.020 180.510 ;
        RECT 231.055 180.465 231.345 180.510 ;
        RECT 234.285 180.465 234.575 180.510 ;
        RECT 214.900 180.310 215.220 180.370 ;
        RECT 214.070 180.170 215.220 180.310 ;
        RECT 207.540 180.110 207.860 180.170 ;
        RECT 211.680 180.110 212.000 180.170 ;
        RECT 213.520 180.110 213.840 180.170 ;
        RECT 214.900 180.110 215.220 180.170 ;
        RECT 217.660 180.110 217.980 180.370 ;
        RECT 218.595 180.310 218.885 180.355 ;
        RECT 220.895 180.310 221.185 180.355 ;
        RECT 218.595 180.170 221.185 180.310 ;
        RECT 218.595 180.125 218.885 180.170 ;
        RECT 220.895 180.125 221.185 180.170 ;
        RECT 221.815 180.310 222.105 180.355 ;
        RECT 223.195 180.310 223.485 180.355 ;
        RECT 221.815 180.170 223.485 180.310 ;
        RECT 221.815 180.125 222.105 180.170 ;
        RECT 223.195 180.125 223.485 180.170 ;
        RECT 224.100 180.110 224.420 180.370 ;
        RECT 225.020 180.310 225.340 180.370 ;
        RECT 235.690 180.310 235.830 181.190 ;
        RECT 237.455 181.145 237.745 181.190 ;
        RECT 225.020 180.170 235.830 180.310 ;
        RECT 225.020 180.110 225.340 180.170 ;
        RECT 236.060 180.110 236.380 180.370 ;
        RECT 236.520 180.110 236.840 180.370 ;
        RECT 77.595 179.815 78.595 180.050 ;
        RECT 83.345 179.815 84.345 180.050 ;
        RECT 64.175 179.585 80.135 179.815 ;
        RECT 81.805 179.585 97.765 179.815 ;
        RECT 63.895 178.380 64.595 179.380 ;
        RECT 77.595 179.350 78.595 179.585 ;
        RECT 77.595 178.175 78.595 178.410 ;
        RECT 80.185 178.380 81.755 179.380 ;
        RECT 83.345 179.350 84.345 179.585 ;
        RECT 83.345 178.175 84.345 178.410 ;
        RECT 97.345 178.380 98.045 179.380 ;
        RECT 64.175 177.945 80.135 178.175 ;
        RECT 81.805 177.945 97.765 178.175 ;
        RECT 77.595 177.710 78.595 177.945 ;
        RECT 83.345 177.710 84.345 177.945 ;
        RECT 77.595 176.795 78.595 177.030 ;
        RECT 83.345 176.795 84.345 177.030 ;
        RECT 64.175 176.565 80.135 176.795 ;
        RECT 81.805 176.565 97.765 176.795 ;
        RECT 63.895 175.360 64.595 176.360 ;
        RECT 77.595 176.330 78.595 176.565 ;
        RECT 77.595 175.155 78.595 175.390 ;
        RECT 80.185 175.360 81.755 176.360 ;
        RECT 83.345 176.330 84.345 176.565 ;
        RECT 83.345 175.155 84.345 175.390 ;
        RECT 97.345 175.360 98.045 176.360 ;
        RECT 64.175 174.925 80.135 175.155 ;
        RECT 81.805 174.925 97.765 175.155 ;
        RECT 77.595 174.690 78.595 174.925 ;
        RECT 83.345 174.690 84.345 174.925 ;
        RECT 64.175 173.545 80.135 173.775 ;
        RECT 81.805 173.545 97.765 173.775 ;
        RECT 63.895 172.340 64.125 173.340 ;
        RECT 80.185 172.340 81.755 173.340 ;
        RECT 97.815 172.340 98.045 173.340 ;
        RECT 64.175 171.905 80.135 172.135 ;
        RECT 81.805 171.905 97.765 172.135 ;
        RECT 98.485 171.445 100.480 180.110 ;
        RECT 62.865 160.555 100.480 171.445 ;
        RECT 5.910 143.155 58.705 143.745 ;
        RECT 5.910 140.725 23.785 143.155 ;
        RECT 24.505 143.045 25.505 143.155 ;
        RECT 24.255 142.435 57.645 142.665 ;
        RECT 24.255 141.275 24.485 142.435 ;
        RECT 28.015 141.965 29.015 142.435 ;
        RECT 32.545 141.275 32.775 142.435 ;
        RECT 36.305 141.965 37.305 142.435 ;
        RECT 40.835 141.275 41.065 142.435 ;
        RECT 44.595 141.965 45.595 142.435 ;
        RECT 49.125 141.275 49.355 142.435 ;
        RECT 52.885 141.965 53.885 142.435 ;
        RECT 57.415 141.275 57.645 142.435 ;
        RECT 24.535 140.885 32.495 141.115 ;
        RECT 32.825 140.885 40.785 141.115 ;
        RECT 41.115 140.885 49.075 141.115 ;
        RECT 49.405 140.885 57.365 141.115 ;
        RECT 5.910 139.725 24.955 140.725 ;
        RECT 32.545 139.725 32.775 140.725 ;
        RECT 40.835 139.725 41.065 140.725 ;
        RECT 49.125 139.725 49.355 140.725 ;
        RECT 56.545 139.725 57.645 140.725 ;
        RECT 5.910 139.175 23.785 139.725 ;
        RECT 24.535 139.335 32.495 139.565 ;
        RECT 32.825 139.335 40.785 139.565 ;
        RECT 41.115 139.335 49.075 139.565 ;
        RECT 49.405 139.335 57.365 139.565 ;
        RECT 5.910 138.175 24.955 139.175 ;
        RECT 32.545 138.175 32.775 139.175 ;
        RECT 40.835 138.175 41.065 139.175 ;
        RECT 49.125 138.175 49.355 139.175 ;
        RECT 53.035 138.175 57.645 139.175 ;
        RECT 5.910 137.925 23.785 138.175 ;
        RECT 5.910 137.075 9.990 137.925 ;
        RECT 11.145 137.465 11.845 137.535 ;
        RECT 14.080 137.465 14.780 137.535 ;
        RECT 15.370 137.465 16.070 137.535 ;
        RECT 18.305 137.465 19.005 137.535 ;
        RECT 11.015 137.235 11.975 137.465 ;
        RECT 13.950 137.235 14.910 137.465 ;
        RECT 15.240 137.235 16.200 137.465 ;
        RECT 18.175 137.235 19.135 137.465 ;
        RECT 5.910 136.075 10.965 137.075 ;
        RECT 12.025 136.925 12.255 137.075 ;
        RECT 11.990 136.225 12.290 136.925 ;
        RECT 12.025 136.075 12.255 136.225 ;
        RECT 5.910 135.225 9.990 136.075 ;
        RECT 13.670 135.825 13.900 137.075 ;
        RECT 14.960 136.925 15.190 137.075 ;
        RECT 16.250 136.925 16.480 137.075 ;
        RECT 14.925 136.225 15.225 136.925 ;
        RECT 16.215 136.225 16.515 136.925 ;
        RECT 14.960 136.075 15.190 136.225 ;
        RECT 16.250 136.075 16.480 136.225 ;
        RECT 13.435 135.525 14.135 135.825 ;
        RECT 17.895 135.225 18.125 137.075 ;
        RECT 19.185 136.775 19.415 137.075 ;
        RECT 19.150 136.075 19.450 136.775 ;
        RECT 20.160 135.745 23.785 137.925 ;
        RECT 24.535 137.785 32.495 138.015 ;
        RECT 32.825 137.785 40.785 138.015 ;
        RECT 41.115 137.785 49.075 138.015 ;
        RECT 49.405 137.785 57.365 138.015 ;
        RECT 24.255 136.465 24.485 137.625 ;
        RECT 28.015 136.465 29.015 136.935 ;
        RECT 32.545 136.465 32.775 137.625 ;
        RECT 36.305 136.465 37.305 136.935 ;
        RECT 40.835 136.465 41.065 137.625 ;
        RECT 44.595 136.465 45.595 136.935 ;
        RECT 49.125 136.465 49.355 137.625 ;
        RECT 52.885 136.465 53.885 136.935 ;
        RECT 57.415 136.465 57.645 137.625 ;
        RECT 24.255 136.235 57.645 136.465 ;
        RECT 24.505 135.745 25.505 135.855 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 20.160 135.225 58.705 135.745 ;
        RECT 5.910 132.225 58.705 135.225 ;
        RECT 62.865 139.455 69.970 160.555 ;
        RECT 71.220 157.040 89.820 159.315 ;
        RECT 71.220 142.990 73.495 157.040 ;
        RECT 76.385 157.030 77.215 157.040 ;
        RECT 80.105 157.030 80.935 157.040 ;
        RECT 83.825 157.030 84.655 157.040 ;
        RECT 74.940 154.420 86.100 155.595 ;
        RECT 74.940 153.050 76.115 154.420 ;
        RECT 76.385 153.310 77.215 154.140 ;
        RECT 77.485 153.050 79.835 154.420 ;
        RECT 80.105 153.310 80.935 154.140 ;
        RECT 81.205 153.050 83.555 154.420 ;
        RECT 83.825 153.310 84.655 154.140 ;
        RECT 84.925 153.050 86.100 154.420 ;
        RECT 74.940 150.700 86.100 153.050 ;
        RECT 74.940 149.330 76.115 150.700 ;
        RECT 76.385 149.590 77.215 150.420 ;
        RECT 77.485 149.330 79.835 150.700 ;
        RECT 80.105 149.590 80.935 150.420 ;
        RECT 81.205 149.330 83.555 150.700 ;
        RECT 83.825 149.590 84.655 150.420 ;
        RECT 84.925 149.330 86.100 150.700 ;
        RECT 74.940 146.980 86.100 149.330 ;
        RECT 74.940 145.610 76.115 146.980 ;
        RECT 76.385 145.870 77.215 146.700 ;
        RECT 77.485 145.610 79.835 146.980 ;
        RECT 80.105 145.870 80.935 146.700 ;
        RECT 81.205 145.610 83.555 146.980 ;
        RECT 83.825 145.870 84.655 146.700 ;
        RECT 84.925 145.610 86.100 146.980 ;
        RECT 74.940 144.435 86.100 145.610 ;
        RECT 87.545 142.990 89.820 157.040 ;
        RECT 71.220 140.715 89.820 142.990 ;
        RECT 91.070 139.455 100.480 160.555 ;
        RECT 101.935 176.325 152.755 178.210 ;
        RECT 101.935 174.870 114.420 176.325 ;
        RECT 115.200 175.635 118.030 176.165 ;
        RECT 119.820 175.635 122.650 176.165 ;
        RECT 124.440 175.635 127.270 176.165 ;
        RECT 129.060 175.635 131.890 176.165 ;
        RECT 133.680 175.635 136.510 176.165 ;
        RECT 138.300 175.635 141.130 176.165 ;
        RECT 142.920 175.635 145.750 176.165 ;
        RECT 147.540 175.635 150.370 176.165 ;
        RECT 114.920 174.870 115.150 175.475 ;
        RECT 101.935 172.215 115.185 174.870 ;
        RECT 101.935 162.685 103.025 172.215 ;
        RECT 103.715 171.610 104.675 171.840 ;
        RECT 105.005 171.610 105.965 171.840 ;
        RECT 103.435 170.840 103.665 171.450 ;
        RECT 103.400 168.540 103.700 170.840 ;
        RECT 103.435 163.450 103.665 168.540 ;
        RECT 104.725 167.140 104.955 171.450 ;
        RECT 106.015 170.840 106.245 171.450 ;
        RECT 105.980 168.540 106.280 170.840 ;
        RECT 104.690 164.840 104.990 167.140 ;
        RECT 104.725 163.450 104.955 164.840 ;
        RECT 106.015 163.450 106.245 168.540 ;
        RECT 103.715 163.060 104.675 163.290 ;
        RECT 105.005 163.060 105.965 163.290 ;
        RECT 103.715 162.990 104.415 163.060 ;
        RECT 105.265 162.990 105.965 163.060 ;
        RECT 106.655 162.685 107.055 172.215 ;
        RECT 110.685 172.070 115.185 172.215 ;
        RECT 107.745 171.610 108.705 171.840 ;
        RECT 109.035 171.610 109.995 171.840 ;
        RECT 107.465 170.840 107.695 171.450 ;
        RECT 107.430 168.540 107.730 170.840 ;
        RECT 107.465 163.450 107.695 168.540 ;
        RECT 108.755 167.140 108.985 171.450 ;
        RECT 110.045 170.840 110.275 171.450 ;
        RECT 110.010 168.540 110.310 170.840 ;
        RECT 108.720 164.840 109.020 167.140 ;
        RECT 108.755 163.450 108.985 164.840 ;
        RECT 110.045 163.450 110.275 168.540 ;
        RECT 110.685 166.625 114.420 172.070 ;
        RECT 114.920 167.475 115.150 172.070 ;
        RECT 115.710 170.895 115.940 175.475 ;
        RECT 116.500 174.870 116.730 175.475 ;
        RECT 116.465 172.070 116.765 174.870 ;
        RECT 115.675 168.095 115.975 170.895 ;
        RECT 115.710 167.475 115.940 168.095 ;
        RECT 116.500 167.475 116.730 172.070 ;
        RECT 117.290 170.895 117.520 175.475 ;
        RECT 118.080 174.870 118.310 175.475 ;
        RECT 119.540 174.870 119.770 175.475 ;
        RECT 118.045 172.070 118.345 174.870 ;
        RECT 119.505 172.070 119.805 174.870 ;
        RECT 117.255 168.095 117.555 170.895 ;
        RECT 117.290 167.475 117.520 168.095 ;
        RECT 118.080 167.475 118.310 172.070 ;
        RECT 119.540 167.475 119.770 172.070 ;
        RECT 120.330 170.895 120.560 175.475 ;
        RECT 121.120 174.870 121.350 175.475 ;
        RECT 121.085 172.070 121.385 174.870 ;
        RECT 120.295 168.095 120.595 170.895 ;
        RECT 120.330 167.475 120.560 168.095 ;
        RECT 121.120 167.475 121.350 172.070 ;
        RECT 121.910 170.895 122.140 175.475 ;
        RECT 122.700 174.870 122.930 175.475 ;
        RECT 124.160 174.870 124.390 175.475 ;
        RECT 122.665 172.070 122.965 174.870 ;
        RECT 124.125 172.070 124.425 174.870 ;
        RECT 121.875 168.095 122.175 170.895 ;
        RECT 121.910 167.475 122.140 168.095 ;
        RECT 122.700 167.475 122.930 172.070 ;
        RECT 124.160 167.475 124.390 172.070 ;
        RECT 124.950 170.895 125.180 175.475 ;
        RECT 125.740 174.870 125.970 175.475 ;
        RECT 125.705 172.070 126.005 174.870 ;
        RECT 124.915 168.095 125.215 170.895 ;
        RECT 124.950 167.475 125.180 168.095 ;
        RECT 125.740 167.475 125.970 172.070 ;
        RECT 126.530 170.895 126.760 175.475 ;
        RECT 127.320 174.870 127.550 175.475 ;
        RECT 128.780 174.870 129.010 175.475 ;
        RECT 127.285 172.070 127.585 174.870 ;
        RECT 128.745 172.070 129.045 174.870 ;
        RECT 126.495 168.095 126.795 170.895 ;
        RECT 126.530 167.475 126.760 168.095 ;
        RECT 127.320 167.475 127.550 172.070 ;
        RECT 128.780 167.475 129.010 172.070 ;
        RECT 129.570 170.895 129.800 175.475 ;
        RECT 130.360 174.870 130.590 175.475 ;
        RECT 130.325 172.070 130.625 174.870 ;
        RECT 129.535 168.095 129.835 170.895 ;
        RECT 129.570 167.475 129.800 168.095 ;
        RECT 130.360 167.475 130.590 172.070 ;
        RECT 131.150 170.895 131.380 175.475 ;
        RECT 131.940 174.870 132.170 175.475 ;
        RECT 133.400 174.870 133.630 175.475 ;
        RECT 131.905 172.070 132.205 174.870 ;
        RECT 133.365 172.070 133.665 174.870 ;
        RECT 131.115 168.095 131.415 170.895 ;
        RECT 131.150 167.475 131.380 168.095 ;
        RECT 131.940 167.475 132.170 172.070 ;
        RECT 133.400 167.475 133.630 172.070 ;
        RECT 134.190 170.895 134.420 175.475 ;
        RECT 134.980 174.870 135.210 175.475 ;
        RECT 134.945 172.070 135.245 174.870 ;
        RECT 134.155 168.095 134.455 170.895 ;
        RECT 134.190 167.475 134.420 168.095 ;
        RECT 134.980 167.475 135.210 172.070 ;
        RECT 135.770 170.895 136.000 175.475 ;
        RECT 136.560 174.870 136.790 175.475 ;
        RECT 138.020 174.870 138.250 175.475 ;
        RECT 136.525 172.070 136.825 174.870 ;
        RECT 137.985 172.070 138.285 174.870 ;
        RECT 135.735 168.095 136.035 170.895 ;
        RECT 135.770 167.475 136.000 168.095 ;
        RECT 136.560 167.475 136.790 172.070 ;
        RECT 138.020 167.475 138.250 172.070 ;
        RECT 138.810 170.895 139.040 175.475 ;
        RECT 139.600 174.870 139.830 175.475 ;
        RECT 139.565 172.070 139.865 174.870 ;
        RECT 138.775 168.095 139.075 170.895 ;
        RECT 138.810 167.475 139.040 168.095 ;
        RECT 139.600 167.475 139.830 172.070 ;
        RECT 140.390 170.895 140.620 175.475 ;
        RECT 141.180 174.870 141.410 175.475 ;
        RECT 142.640 174.870 142.870 175.475 ;
        RECT 141.145 172.070 141.445 174.870 ;
        RECT 142.605 172.070 142.905 174.870 ;
        RECT 140.355 168.095 140.655 170.895 ;
        RECT 140.390 167.475 140.620 168.095 ;
        RECT 141.180 167.475 141.410 172.070 ;
        RECT 142.640 167.475 142.870 172.070 ;
        RECT 143.430 170.895 143.660 175.475 ;
        RECT 144.220 174.870 144.450 175.475 ;
        RECT 144.185 172.070 144.485 174.870 ;
        RECT 143.395 168.095 143.695 170.895 ;
        RECT 143.430 167.475 143.660 168.095 ;
        RECT 144.220 167.475 144.450 172.070 ;
        RECT 145.010 170.895 145.240 175.475 ;
        RECT 145.800 174.870 146.030 175.475 ;
        RECT 147.260 174.870 147.490 175.475 ;
        RECT 145.765 172.070 146.065 174.870 ;
        RECT 147.225 172.070 147.525 174.870 ;
        RECT 144.975 168.095 145.275 170.895 ;
        RECT 145.010 167.475 145.240 168.095 ;
        RECT 145.800 167.475 146.030 172.070 ;
        RECT 147.260 167.475 147.490 172.070 ;
        RECT 148.050 170.895 148.280 175.475 ;
        RECT 148.840 174.870 149.070 175.475 ;
        RECT 148.805 172.070 149.105 174.870 ;
        RECT 148.015 168.095 148.315 170.895 ;
        RECT 148.050 167.475 148.280 168.095 ;
        RECT 148.840 167.475 149.070 172.070 ;
        RECT 149.630 170.895 149.860 175.475 ;
        RECT 150.420 174.870 150.650 175.475 ;
        RECT 150.385 172.070 150.685 174.870 ;
        RECT 149.595 168.095 149.895 170.895 ;
        RECT 149.630 167.475 149.860 168.095 ;
        RECT 150.420 167.475 150.650 172.070 ;
        RECT 115.200 167.085 115.660 167.315 ;
        RECT 115.990 167.085 116.450 167.315 ;
        RECT 116.780 167.085 117.240 167.315 ;
        RECT 117.570 167.085 118.030 167.315 ;
        RECT 119.820 167.085 120.280 167.315 ;
        RECT 120.610 167.085 121.070 167.315 ;
        RECT 121.400 167.085 121.860 167.315 ;
        RECT 122.190 167.085 122.650 167.315 ;
        RECT 124.440 167.085 124.900 167.315 ;
        RECT 125.230 167.085 125.690 167.315 ;
        RECT 126.020 167.085 126.480 167.315 ;
        RECT 126.810 167.085 127.270 167.315 ;
        RECT 129.060 167.085 129.520 167.315 ;
        RECT 129.850 167.085 130.310 167.315 ;
        RECT 130.640 167.085 131.100 167.315 ;
        RECT 131.430 167.085 131.890 167.315 ;
        RECT 133.680 167.085 134.140 167.315 ;
        RECT 134.470 167.085 134.930 167.315 ;
        RECT 135.260 167.085 135.720 167.315 ;
        RECT 136.050 167.085 136.510 167.315 ;
        RECT 138.300 167.085 138.760 167.315 ;
        RECT 139.090 167.085 139.550 167.315 ;
        RECT 139.880 167.085 140.340 167.315 ;
        RECT 140.670 167.085 141.130 167.315 ;
        RECT 142.920 167.085 143.380 167.315 ;
        RECT 143.710 167.085 144.170 167.315 ;
        RECT 144.500 167.085 144.960 167.315 ;
        RECT 145.290 167.085 145.750 167.315 ;
        RECT 147.540 167.085 148.000 167.315 ;
        RECT 148.330 167.085 148.790 167.315 ;
        RECT 149.120 167.085 149.580 167.315 ;
        RECT 149.910 167.085 150.370 167.315 ;
        RECT 151.150 166.625 152.755 176.325 ;
        RECT 110.685 166.035 152.755 166.625 ;
        RECT 107.745 163.060 108.705 163.290 ;
        RECT 109.035 163.060 109.995 163.290 ;
        RECT 107.745 162.990 108.445 163.060 ;
        RECT 109.295 162.990 109.995 163.060 ;
        RECT 110.685 162.685 114.420 166.035 ;
        RECT 134.745 165.030 135.445 165.080 ;
        RECT 146.905 165.030 147.605 165.080 ;
        RECT 134.745 164.430 147.605 165.030 ;
        RECT 134.745 164.380 135.445 164.430 ;
        RECT 146.905 164.380 147.605 164.430 ;
        RECT 133.735 163.740 134.435 163.790 ;
        RECT 143.985 163.740 144.685 163.790 ;
        RECT 133.735 163.140 144.685 163.740 ;
        RECT 133.735 163.090 134.435 163.140 ;
        RECT 143.985 163.090 144.685 163.140 ;
        RECT 101.935 162.285 114.420 162.685 ;
        RECT 101.935 158.755 103.025 162.285 ;
        RECT 103.435 160.445 103.665 161.520 ;
        RECT 103.400 159.745 103.700 160.445 ;
        RECT 103.435 159.520 103.665 159.745 ;
        RECT 104.725 159.520 104.955 162.285 ;
        RECT 106.015 160.445 106.245 161.520 ;
        RECT 105.980 159.745 106.280 160.445 ;
        RECT 106.015 159.520 106.245 159.745 ;
        RECT 103.715 159.130 104.675 159.360 ;
        RECT 105.005 159.130 105.965 159.360 ;
        RECT 103.845 159.060 104.545 159.130 ;
        RECT 105.135 159.060 105.835 159.130 ;
        RECT 106.655 158.755 107.055 162.285 ;
        RECT 107.465 160.445 107.695 161.520 ;
        RECT 107.430 159.745 107.730 160.445 ;
        RECT 107.465 159.520 107.695 159.745 ;
        RECT 108.755 159.520 108.985 162.285 ;
        RECT 110.045 160.445 110.275 161.520 ;
        RECT 110.010 159.745 110.310 160.445 ;
        RECT 110.045 159.520 110.275 159.745 ;
        RECT 107.745 159.130 108.705 159.360 ;
        RECT 109.035 159.130 109.995 159.360 ;
        RECT 107.875 159.060 108.575 159.130 ;
        RECT 109.165 159.060 109.865 159.130 ;
        RECT 110.685 158.755 114.420 162.285 ;
        RECT 136.825 162.330 137.525 162.400 ;
        RECT 143.985 162.330 144.685 162.400 ;
        RECT 136.825 161.730 144.685 162.330 ;
        RECT 136.825 161.700 137.525 161.730 ;
        RECT 143.985 161.700 144.685 161.730 ;
        RECT 134.745 160.160 135.445 160.210 ;
        RECT 145.575 160.160 146.275 160.210 ;
        RECT 134.745 159.560 146.275 160.160 ;
        RECT 134.745 159.510 135.445 159.560 ;
        RECT 145.575 159.510 146.275 159.560 ;
        RECT 101.935 157.850 114.420 158.755 ;
        RECT 141.665 159.150 142.365 159.200 ;
        RECT 148.605 159.150 149.305 159.200 ;
        RECT 141.665 158.550 149.305 159.150 ;
        RECT 141.665 158.500 142.365 158.550 ;
        RECT 148.605 158.500 149.305 158.550 ;
        RECT 153.960 158.060 155.900 180.110 ;
        RECT 165.150 179.490 239.210 179.970 ;
        RECT 168.440 179.090 168.760 179.350 ;
        RECT 169.835 179.290 170.125 179.335 ;
        RECT 170.740 179.290 171.060 179.350 ;
        RECT 168.990 179.150 171.060 179.290 ;
        RECT 168.990 178.610 169.130 179.150 ;
        RECT 169.835 179.105 170.125 179.150 ;
        RECT 170.740 179.090 171.060 179.150 ;
        RECT 173.975 179.290 174.265 179.335 ;
        RECT 175.340 179.290 175.660 179.350 ;
        RECT 173.975 179.150 175.660 179.290 ;
        RECT 173.975 179.105 174.265 179.150 ;
        RECT 175.340 179.090 175.660 179.150 ;
        RECT 175.800 179.290 176.120 179.350 ;
        RECT 178.575 179.290 178.865 179.335 ;
        RECT 175.800 179.150 178.865 179.290 ;
        RECT 175.800 179.090 176.120 179.150 ;
        RECT 178.575 179.105 178.865 179.150 ;
        RECT 179.495 179.105 179.785 179.335 ;
        RECT 180.860 179.290 181.180 179.350 ;
        RECT 182.715 179.290 183.005 179.335 ;
        RECT 180.860 179.150 183.005 179.290 ;
        RECT 169.360 178.950 169.680 179.010 ;
        RECT 177.640 178.950 177.960 179.010 ;
        RECT 179.570 178.950 179.710 179.105 ;
        RECT 180.860 179.090 181.180 179.150 ;
        RECT 182.715 179.105 183.005 179.150 ;
        RECT 184.540 179.090 184.860 179.350 ;
        RECT 185.000 179.290 185.320 179.350 ;
        RECT 186.855 179.290 187.145 179.335 ;
        RECT 185.000 179.150 187.145 179.290 ;
        RECT 185.000 179.090 185.320 179.150 ;
        RECT 186.855 179.105 187.145 179.150 ;
        RECT 188.235 179.290 188.525 179.335 ;
        RECT 189.140 179.290 189.460 179.350 ;
        RECT 188.235 179.150 189.460 179.290 ;
        RECT 188.235 179.105 188.525 179.150 ;
        RECT 189.140 179.090 189.460 179.150 ;
        RECT 189.600 179.090 189.920 179.350 ;
        RECT 190.535 179.105 190.825 179.335 ;
        RECT 191.440 179.290 191.760 179.350 ;
        RECT 192.835 179.290 193.125 179.335 ;
        RECT 191.440 179.150 193.125 179.290 ;
        RECT 169.360 178.810 174.650 178.950 ;
        RECT 169.360 178.750 169.680 178.810 ;
        RECT 168.990 178.470 171.890 178.610 ;
        RECT 167.520 178.070 167.840 178.330 ;
        RECT 168.900 178.270 169.220 178.330 ;
        RECT 169.375 178.270 169.665 178.315 ;
        RECT 168.900 178.130 169.665 178.270 ;
        RECT 168.900 178.070 169.220 178.130 ;
        RECT 169.375 178.085 169.665 178.130 ;
        RECT 169.820 178.270 170.140 178.330 ;
        RECT 171.750 178.315 171.890 178.470 ;
        RECT 172.580 178.410 172.900 178.670 ;
        RECT 170.755 178.270 171.045 178.315 ;
        RECT 169.820 178.130 171.045 178.270 ;
        RECT 169.450 177.930 169.590 178.085 ;
        RECT 169.820 178.070 170.140 178.130 ;
        RECT 170.755 178.085 171.045 178.130 ;
        RECT 171.675 178.085 171.965 178.315 ;
        RECT 172.670 178.270 172.810 178.410 ;
        RECT 173.055 178.270 173.345 178.315 ;
        RECT 172.670 178.130 173.345 178.270 ;
        RECT 174.510 178.270 174.650 178.810 ;
        RECT 177.640 178.810 179.710 178.950 ;
        RECT 177.640 178.750 177.960 178.810 ;
        RECT 181.780 178.750 182.100 179.010 ;
        RECT 182.255 178.950 182.545 178.995 ;
        RECT 182.255 178.810 182.930 178.950 ;
        RECT 182.255 178.765 182.545 178.810 ;
        RECT 174.895 178.610 175.185 178.655 ;
        RECT 176.720 178.610 177.040 178.670 ;
        RECT 181.870 178.610 182.010 178.750 ;
        RECT 182.790 178.670 182.930 178.810 ;
        RECT 174.895 178.470 182.010 178.610 ;
        RECT 174.895 178.425 175.185 178.470 ;
        RECT 176.720 178.410 177.040 178.470 ;
        RECT 182.700 178.410 183.020 178.670 ;
        RECT 184.630 178.610 184.770 179.090 ;
        RECT 189.690 178.950 189.830 179.090 ;
        RECT 185.090 178.810 189.830 178.950 ;
        RECT 190.610 178.950 190.750 179.105 ;
        RECT 191.440 179.090 191.760 179.150 ;
        RECT 192.835 179.105 193.125 179.150 ;
        RECT 193.295 179.290 193.585 179.335 ;
        RECT 193.740 179.290 194.060 179.350 ;
        RECT 193.295 179.150 194.060 179.290 ;
        RECT 193.295 179.105 193.585 179.150 ;
        RECT 193.740 179.090 194.060 179.150 ;
        RECT 194.200 179.290 194.520 179.350 ;
        RECT 196.055 179.290 196.345 179.335 ;
        RECT 199.260 179.290 199.580 179.350 ;
        RECT 194.200 179.150 196.345 179.290 ;
        RECT 194.200 179.090 194.520 179.150 ;
        RECT 196.055 179.105 196.345 179.150 ;
        RECT 198.890 179.150 199.580 179.290 ;
        RECT 194.660 178.950 194.980 179.010 ;
        RECT 190.610 178.810 194.980 178.950 ;
        RECT 185.090 178.655 185.230 178.810 ;
        RECT 194.660 178.750 194.980 178.810 ;
        RECT 195.580 178.750 195.900 179.010 ;
        RECT 197.420 178.950 197.740 179.010 ;
        RECT 198.890 178.950 199.030 179.150 ;
        RECT 199.260 179.090 199.580 179.150 ;
        RECT 202.940 179.290 203.260 179.350 ;
        RECT 203.415 179.290 203.705 179.335 ;
        RECT 202.940 179.150 203.705 179.290 ;
        RECT 202.940 179.090 203.260 179.150 ;
        RECT 203.415 179.105 203.705 179.150 ;
        RECT 204.320 179.290 204.640 179.350 ;
        RECT 207.095 179.290 207.385 179.335 ;
        RECT 215.820 179.290 216.140 179.350 ;
        RECT 236.520 179.290 236.840 179.350 ;
        RECT 204.320 179.150 207.385 179.290 ;
        RECT 204.320 179.090 204.640 179.150 ;
        RECT 207.095 179.105 207.385 179.150 ;
        RECT 208.550 179.150 215.590 179.290 ;
        RECT 197.420 178.810 199.030 178.950 ;
        RECT 197.420 178.750 197.740 178.810 ;
        RECT 184.170 178.470 184.770 178.610 ;
        RECT 179.940 178.270 180.260 178.330 ;
        RECT 180.875 178.270 181.165 178.315 ;
        RECT 174.510 178.130 179.710 178.270 ;
        RECT 173.055 178.085 173.345 178.130 ;
        RECT 176.275 177.930 176.565 177.975 ;
        RECT 169.450 177.790 176.565 177.930 ;
        RECT 179.570 177.930 179.710 178.130 ;
        RECT 179.940 178.130 181.165 178.270 ;
        RECT 179.940 178.070 180.260 178.130 ;
        RECT 180.875 178.085 181.165 178.130 ;
        RECT 181.335 178.270 181.625 178.315 ;
        RECT 181.780 178.270 182.100 178.330 ;
        RECT 181.335 178.130 182.100 178.270 ;
        RECT 181.335 178.085 181.625 178.130 ;
        RECT 181.780 178.070 182.100 178.130 ;
        RECT 182.240 177.930 182.560 177.990 ;
        RECT 179.570 177.790 182.560 177.930 ;
        RECT 176.275 177.745 176.565 177.790 ;
        RECT 176.350 177.590 176.490 177.745 ;
        RECT 182.240 177.730 182.560 177.790 ;
        RECT 180.860 177.590 181.180 177.650 ;
        RECT 176.350 177.450 181.180 177.590 ;
        RECT 184.170 177.590 184.310 178.470 ;
        RECT 185.015 178.425 185.305 178.655 ;
        RECT 185.935 178.610 186.225 178.655 ;
        RECT 186.380 178.610 186.700 178.670 ;
        RECT 185.935 178.470 186.700 178.610 ;
        RECT 185.935 178.425 186.225 178.470 ;
        RECT 186.380 178.410 186.700 178.470 ;
        RECT 190.060 178.610 190.380 178.670 ;
        RECT 193.280 178.610 193.600 178.670 ;
        RECT 198.890 178.655 199.030 178.810 ;
        RECT 205.715 178.950 206.005 178.995 ;
        RECT 208.550 178.950 208.690 179.150 ;
        RECT 205.715 178.810 208.690 178.950 ;
        RECT 208.885 178.950 209.175 178.995 ;
        RECT 212.115 178.950 212.405 178.995 ;
        RECT 215.450 178.950 215.590 179.150 ;
        RECT 215.820 179.150 236.840 179.290 ;
        RECT 215.820 179.090 216.140 179.150 ;
        RECT 236.520 179.090 236.840 179.150 ;
        RECT 218.580 178.950 218.900 179.010 ;
        RECT 208.885 178.810 212.405 178.950 ;
        RECT 205.715 178.765 206.005 178.810 ;
        RECT 208.885 178.765 209.175 178.810 ;
        RECT 212.115 178.765 212.405 178.810 ;
        RECT 212.690 178.810 215.130 178.950 ;
        RECT 215.450 178.810 218.900 178.950 ;
        RECT 190.060 178.470 193.600 178.610 ;
        RECT 190.060 178.410 190.380 178.470 ;
        RECT 193.280 178.410 193.600 178.470 ;
        RECT 195.210 178.470 198.595 178.610 ;
        RECT 184.540 178.070 184.860 178.330 ;
        RECT 187.775 178.085 188.065 178.315 ;
        RECT 189.155 178.085 189.445 178.315 ;
        RECT 184.630 177.930 184.770 178.070 ;
        RECT 186.380 177.930 186.700 177.990 ;
        RECT 184.630 177.790 186.700 177.930 ;
        RECT 186.380 177.730 186.700 177.790 ;
        RECT 184.555 177.590 184.845 177.635 ;
        RECT 184.170 177.450 184.845 177.590 ;
        RECT 187.850 177.590 187.990 178.085 ;
        RECT 189.230 177.930 189.370 178.085 ;
        RECT 189.600 178.070 189.920 178.330 ;
        RECT 191.900 178.070 192.220 178.330 ;
        RECT 194.200 178.070 194.520 178.330 ;
        RECT 194.675 178.270 194.965 178.315 ;
        RECT 195.210 178.270 195.350 178.470 ;
        RECT 194.675 178.130 195.350 178.270 ;
        RECT 194.675 178.085 194.965 178.130 ;
        RECT 195.580 178.070 195.900 178.330 ;
        RECT 198.455 178.270 198.595 178.470 ;
        RECT 198.815 178.425 199.105 178.655 ;
        RECT 206.620 178.610 206.940 178.670 ;
        RECT 212.690 178.610 212.830 178.810 ;
        RECT 206.620 178.470 212.830 178.610 ;
        RECT 213.075 178.610 213.365 178.655 ;
        RECT 213.520 178.610 213.840 178.670 ;
        RECT 214.990 178.610 215.130 178.810 ;
        RECT 218.580 178.750 218.900 178.810 ;
        RECT 223.195 178.950 223.485 178.995 ;
        RECT 223.640 178.950 223.960 179.010 ;
        RECT 223.195 178.810 223.960 178.950 ;
        RECT 223.195 178.765 223.485 178.810 ;
        RECT 215.375 178.610 215.665 178.655 ;
        RECT 223.270 178.610 223.410 178.765 ;
        RECT 223.640 178.750 223.960 178.810 ;
        RECT 224.155 178.950 224.445 178.995 ;
        RECT 227.385 178.950 227.675 178.995 ;
        RECT 224.155 178.810 227.675 178.950 ;
        RECT 224.155 178.765 224.445 178.810 ;
        RECT 227.385 178.765 227.675 178.810 ;
        RECT 228.240 178.950 228.560 179.010 ;
        RECT 229.175 178.950 229.465 178.995 ;
        RECT 228.240 178.810 229.465 178.950 ;
        RECT 228.240 178.750 228.560 178.810 ;
        RECT 229.175 178.765 229.465 178.810 ;
        RECT 232.380 178.750 232.700 179.010 ;
        RECT 233.760 178.950 234.080 179.010 ;
        RECT 235.615 178.950 235.905 178.995 ;
        RECT 233.760 178.810 235.905 178.950 ;
        RECT 233.760 178.750 234.080 178.810 ;
        RECT 235.615 178.765 235.905 178.810 ;
        RECT 213.075 178.470 214.670 178.610 ;
        RECT 214.990 178.470 215.665 178.610 ;
        RECT 206.620 178.410 206.940 178.470 ;
        RECT 213.075 178.425 213.365 178.470 ;
        RECT 213.520 178.410 213.840 178.470 ;
        RECT 200.640 178.270 200.960 178.330 ;
        RECT 198.455 178.130 200.960 178.270 ;
        RECT 200.640 178.070 200.960 178.130 ;
        RECT 201.115 178.085 201.405 178.315 ;
        RECT 195.670 177.930 195.810 178.070 ;
        RECT 198.355 177.930 198.645 177.975 ;
        RECT 189.230 177.790 195.350 177.930 ;
        RECT 195.670 177.790 198.645 177.930 ;
        RECT 190.060 177.590 190.380 177.650 ;
        RECT 187.850 177.450 190.380 177.590 ;
        RECT 195.210 177.590 195.350 177.790 ;
        RECT 198.355 177.745 198.645 177.790 ;
        RECT 199.260 177.730 199.580 177.990 ;
        RECT 201.190 177.930 201.330 178.085 ;
        RECT 202.480 178.070 202.800 178.330 ;
        RECT 204.780 178.070 205.100 178.330 ;
        RECT 207.965 178.270 208.255 178.315 ;
        RECT 209.805 178.270 210.095 178.315 ;
        RECT 207.965 178.130 210.095 178.270 ;
        RECT 207.965 178.085 208.255 178.130 ;
        RECT 209.805 178.085 210.095 178.130 ;
        RECT 210.300 178.070 210.620 178.330 ;
        RECT 211.220 178.315 211.540 178.330 ;
        RECT 211.110 178.085 211.540 178.315 ;
        RECT 211.220 178.070 211.540 178.085 ;
        RECT 211.680 178.070 212.000 178.330 ;
        RECT 212.150 178.270 212.440 178.315 ;
        RECT 213.990 178.270 214.280 178.315 ;
        RECT 212.150 178.130 214.280 178.270 ;
        RECT 214.530 178.270 214.670 178.470 ;
        RECT 215.375 178.425 215.665 178.470 ;
        RECT 215.910 178.470 223.410 178.610 ;
        RECT 225.265 178.610 225.555 178.655 ;
        RECT 232.470 178.610 232.610 178.750 ;
        RECT 225.265 178.470 232.610 178.610 ;
        RECT 215.910 178.270 216.050 178.470 ;
        RECT 225.265 178.425 225.555 178.470 ;
        RECT 232.840 178.410 233.160 178.670 ;
        RECT 214.530 178.130 216.050 178.270 ;
        RECT 212.150 178.085 212.440 178.130 ;
        RECT 213.990 178.085 214.280 178.130 ;
        RECT 216.280 178.070 216.600 178.330 ;
        RECT 217.200 178.070 217.520 178.330 ;
        RECT 218.595 178.085 218.885 178.315 ;
        RECT 206.160 177.930 206.480 177.990 ;
        RECT 201.190 177.790 206.480 177.930 ;
        RECT 206.160 177.730 206.480 177.790 ;
        RECT 208.470 177.930 208.760 177.975 ;
        RECT 209.390 177.930 209.680 177.975 ;
        RECT 214.910 177.930 215.200 177.975 ;
        RECT 208.470 177.790 215.200 177.930 ;
        RECT 208.470 177.745 208.760 177.790 ;
        RECT 209.390 177.745 209.680 177.790 ;
        RECT 214.910 177.745 215.200 177.790 ;
        RECT 215.360 177.930 215.680 177.990 ;
        RECT 218.670 177.930 218.810 178.085 ;
        RECT 219.040 178.070 219.360 178.330 ;
        RECT 219.500 178.270 219.820 178.330 ;
        RECT 219.975 178.270 220.265 178.315 ;
        RECT 219.500 178.130 220.265 178.270 ;
        RECT 219.500 178.070 219.820 178.130 ;
        RECT 219.975 178.085 220.265 178.130 ;
        RECT 220.895 178.085 221.185 178.315 ;
        RECT 222.280 178.270 222.570 178.315 ;
        RECT 224.120 178.270 224.410 178.315 ;
        RECT 222.280 178.130 224.410 178.270 ;
        RECT 222.280 178.085 222.570 178.130 ;
        RECT 224.120 178.085 224.410 178.130 ;
        RECT 215.360 177.790 218.810 177.930 ;
        RECT 215.360 177.730 215.680 177.790 ;
        RECT 196.960 177.590 197.280 177.650 ;
        RECT 195.210 177.450 197.280 177.590 ;
        RECT 180.860 177.390 181.180 177.450 ;
        RECT 184.555 177.405 184.845 177.450 ;
        RECT 190.060 177.390 190.380 177.450 ;
        RECT 196.960 177.390 197.280 177.450 ;
        RECT 197.895 177.590 198.185 177.635 ;
        RECT 199.350 177.590 199.490 177.730 ;
        RECT 197.895 177.450 199.490 177.590 ;
        RECT 202.035 177.590 202.325 177.635 ;
        RECT 210.300 177.590 210.620 177.650 ;
        RECT 202.035 177.450 210.620 177.590 ;
        RECT 197.895 177.405 198.185 177.450 ;
        RECT 202.035 177.405 202.325 177.450 ;
        RECT 210.300 177.390 210.620 177.450 ;
        RECT 211.680 177.590 212.000 177.650 ;
        RECT 213.980 177.590 214.300 177.650 ;
        RECT 211.680 177.450 214.300 177.590 ;
        RECT 211.680 177.390 212.000 177.450 ;
        RECT 213.980 177.390 214.300 177.450 ;
        RECT 218.135 177.590 218.425 177.635 ;
        RECT 219.130 177.590 219.270 178.070 ;
        RECT 218.135 177.450 219.270 177.590 ;
        RECT 219.515 177.590 219.805 177.635 ;
        RECT 220.970 177.590 221.110 178.085 ;
        RECT 224.560 178.070 224.880 178.330 ;
        RECT 225.940 178.070 226.260 178.330 ;
        RECT 226.465 178.270 226.755 178.315 ;
        RECT 228.305 178.270 228.595 178.315 ;
        RECT 226.465 178.130 228.595 178.270 ;
        RECT 226.465 178.085 226.755 178.130 ;
        RECT 228.305 178.085 228.595 178.130 ;
        RECT 229.160 178.270 229.480 178.330 ;
        RECT 231.015 178.270 231.305 178.315 ;
        RECT 231.460 178.270 231.780 178.330 ;
        RECT 229.160 178.130 230.770 178.270 ;
        RECT 229.160 178.070 229.480 178.130 ;
        RECT 221.360 177.930 221.650 177.975 ;
        RECT 226.880 177.930 227.170 177.975 ;
        RECT 227.800 177.930 228.090 177.975 ;
        RECT 221.360 177.790 228.090 177.930 ;
        RECT 221.360 177.745 221.650 177.790 ;
        RECT 226.880 177.745 227.170 177.790 ;
        RECT 227.800 177.745 228.090 177.790 ;
        RECT 228.330 177.790 230.310 177.930 ;
        RECT 219.515 177.450 221.110 177.590 ;
        RECT 221.800 177.590 222.120 177.650 ;
        RECT 228.330 177.590 228.470 177.790 ;
        RECT 230.170 177.635 230.310 177.790 ;
        RECT 221.800 177.450 228.470 177.590 ;
        RECT 218.135 177.405 218.425 177.450 ;
        RECT 219.515 177.405 219.805 177.450 ;
        RECT 221.800 177.390 222.120 177.450 ;
        RECT 230.095 177.405 230.385 177.635 ;
        RECT 230.630 177.590 230.770 178.130 ;
        RECT 231.015 178.130 231.780 178.270 ;
        RECT 231.015 178.085 231.305 178.130 ;
        RECT 231.460 178.070 231.780 178.130 ;
        RECT 232.380 178.070 232.700 178.330 ;
        RECT 232.930 177.635 233.070 178.410 ;
        RECT 233.760 178.070 234.080 178.330 ;
        RECT 235.140 178.070 235.460 178.330 ;
        RECT 236.520 178.070 236.840 178.330 ;
        RECT 231.475 177.590 231.765 177.635 ;
        RECT 230.630 177.450 231.765 177.590 ;
        RECT 231.475 177.405 231.765 177.450 ;
        RECT 232.855 177.405 233.145 177.635 ;
        RECT 234.220 177.390 234.540 177.650 ;
        RECT 165.150 176.770 239.990 177.250 ;
        RECT 167.980 176.570 168.300 176.630 ;
        RECT 178.100 176.570 178.420 176.630 ;
        RECT 167.980 176.430 178.420 176.570 ;
        RECT 167.980 176.370 168.300 176.430 ;
        RECT 178.100 176.370 178.420 176.430 ;
        RECT 180.860 176.370 181.180 176.630 ;
        RECT 183.620 176.570 183.940 176.630 ;
        RECT 186.380 176.570 186.700 176.630 ;
        RECT 183.620 176.430 186.700 176.570 ;
        RECT 183.620 176.370 183.940 176.430 ;
        RECT 186.380 176.370 186.700 176.430 ;
        RECT 190.060 176.570 190.380 176.630 ;
        RECT 195.580 176.570 195.900 176.630 ;
        RECT 190.060 176.430 195.900 176.570 ;
        RECT 190.060 176.370 190.380 176.430 ;
        RECT 195.580 176.370 195.900 176.430 ;
        RECT 200.180 176.570 200.500 176.630 ;
        RECT 201.100 176.570 201.420 176.630 ;
        RECT 200.180 176.430 201.420 176.570 ;
        RECT 200.180 176.370 200.500 176.430 ;
        RECT 201.100 176.370 201.420 176.430 ;
        RECT 202.940 176.570 203.260 176.630 ;
        RECT 203.860 176.570 204.180 176.630 ;
        RECT 202.940 176.430 204.180 176.570 ;
        RECT 202.940 176.370 203.260 176.430 ;
        RECT 203.860 176.370 204.180 176.430 ;
        RECT 210.300 176.370 210.620 176.630 ;
        RECT 211.220 176.370 211.540 176.630 ;
        RECT 213.980 176.570 214.300 176.630 ;
        RECT 214.900 176.570 215.220 176.630 ;
        RECT 213.980 176.430 215.220 176.570 ;
        RECT 213.980 176.370 214.300 176.430 ;
        RECT 214.900 176.370 215.220 176.430 ;
        RECT 221.340 176.570 221.660 176.630 ;
        RECT 223.180 176.570 223.500 176.630 ;
        RECT 221.340 176.430 223.500 176.570 ;
        RECT 221.340 176.370 221.660 176.430 ;
        RECT 223.180 176.370 223.500 176.430 ;
        RECT 225.020 176.570 225.340 176.630 ;
        RECT 233.300 176.570 233.620 176.630 ;
        RECT 225.020 176.430 233.620 176.570 ;
        RECT 225.020 176.370 225.340 176.430 ;
        RECT 233.300 176.370 233.620 176.430 ;
        RECT 234.220 176.370 234.540 176.630 ;
        RECT 166.600 176.230 166.920 176.290 ;
        RECT 176.260 176.230 176.580 176.290 ;
        RECT 166.600 176.090 176.580 176.230 ;
        RECT 166.600 176.030 166.920 176.090 ;
        RECT 176.260 176.030 176.580 176.090 ;
        RECT 180.950 175.890 181.090 176.370 ;
        RECT 181.780 176.230 182.100 176.290 ;
        RECT 193.740 176.230 194.060 176.290 ;
        RECT 181.780 176.090 194.060 176.230 ;
        RECT 181.780 176.030 182.100 176.090 ;
        RECT 193.740 176.030 194.060 176.090 ;
        RECT 194.660 176.230 194.980 176.290 ;
        RECT 199.260 176.230 199.580 176.290 ;
        RECT 194.660 176.090 199.580 176.230 ;
        RECT 194.660 176.030 194.980 176.090 ;
        RECT 199.260 176.030 199.580 176.090 ;
        RECT 191.900 175.890 192.220 175.950 ;
        RECT 198.340 175.890 198.660 175.950 ;
        RECT 180.950 175.750 191.670 175.890 ;
        RECT 167.520 175.550 167.840 175.610 ;
        RECT 190.980 175.550 191.300 175.610 ;
        RECT 167.520 175.410 191.300 175.550 ;
        RECT 191.530 175.550 191.670 175.750 ;
        RECT 191.900 175.750 198.660 175.890 ;
        RECT 191.900 175.690 192.220 175.750 ;
        RECT 198.340 175.690 198.660 175.750 ;
        RECT 197.420 175.550 197.740 175.610 ;
        RECT 191.530 175.410 197.740 175.550 ;
        RECT 167.520 175.350 167.840 175.410 ;
        RECT 190.980 175.350 191.300 175.410 ;
        RECT 197.420 175.350 197.740 175.410 ;
        RECT 210.390 175.210 210.530 176.370 ;
        RECT 211.310 175.890 211.450 176.370 ;
        RECT 216.740 176.230 217.060 176.290 ;
        RECT 231.460 176.230 231.780 176.290 ;
        RECT 216.740 176.090 231.780 176.230 ;
        RECT 216.740 176.030 217.060 176.090 ;
        RECT 231.460 176.030 231.780 176.090 ;
        RECT 234.310 175.890 234.450 176.370 ;
        RECT 211.310 175.750 234.450 175.890 ;
        RECT 222.260 175.550 222.580 175.610 ;
        RECT 236.520 175.550 236.840 175.610 ;
        RECT 222.260 175.410 236.840 175.550 ;
        RECT 222.260 175.350 222.580 175.410 ;
        RECT 236.520 175.350 236.840 175.410 ;
        RECT 225.940 175.210 226.260 175.270 ;
        RECT 210.390 175.070 226.260 175.210 ;
        RECT 225.940 175.010 226.260 175.070 ;
        RECT 226.860 175.210 227.180 175.270 ;
        RECT 237.900 175.210 238.220 175.270 ;
        RECT 226.860 175.070 238.220 175.210 ;
        RECT 226.860 175.010 227.180 175.070 ;
        RECT 237.900 175.010 238.220 175.070 ;
        RECT 220.420 174.870 220.740 174.930 ;
        RECT 235.140 174.870 235.460 174.930 ;
        RECT 220.420 174.730 235.460 174.870 ;
        RECT 220.420 174.670 220.740 174.730 ;
        RECT 235.140 174.670 235.460 174.730 ;
        RECT 115.985 156.185 155.900 158.060 ;
        RECT 115.985 156.060 116.575 156.185 ;
        RECT 102.625 155.660 116.575 156.060 ;
        RECT 102.625 152.040 103.025 155.660 ;
        RECT 103.715 155.055 104.675 155.385 ;
        RECT 105.005 155.055 105.965 155.385 ;
        RECT 103.435 153.515 103.665 154.850 ;
        RECT 103.400 152.815 103.700 153.515 ;
        RECT 104.725 152.040 104.955 154.850 ;
        RECT 106.015 154.585 106.245 154.850 ;
        RECT 105.980 153.885 106.280 154.585 ;
        RECT 106.015 152.850 106.245 153.885 ;
        RECT 106.655 152.040 107.055 155.660 ;
        RECT 107.745 155.055 108.705 155.385 ;
        RECT 109.035 155.055 109.995 155.385 ;
        RECT 107.465 153.515 107.695 154.850 ;
        RECT 107.430 152.815 107.730 153.515 ;
        RECT 108.755 152.040 108.985 154.850 ;
        RECT 110.045 154.585 110.275 154.850 ;
        RECT 110.010 153.885 110.310 154.585 ;
        RECT 110.045 152.850 110.275 153.885 ;
        RECT 110.685 152.040 116.575 155.660 ;
        RECT 102.625 151.550 116.575 152.040 ;
        RECT 102.625 142.020 103.025 151.550 ;
        RECT 103.715 151.035 104.675 151.365 ;
        RECT 105.005 151.035 105.965 151.365 ;
        RECT 103.435 145.785 103.665 150.830 ;
        RECT 104.725 149.485 104.955 150.830 ;
        RECT 104.690 147.185 104.990 149.485 ;
        RECT 103.400 143.485 103.700 145.785 ;
        RECT 103.435 142.830 103.665 143.485 ;
        RECT 104.725 142.830 104.955 147.185 ;
        RECT 106.015 145.785 106.245 150.830 ;
        RECT 105.980 143.485 106.280 145.785 ;
        RECT 106.015 142.830 106.245 143.485 ;
        RECT 103.715 142.395 104.675 142.625 ;
        RECT 105.005 142.395 105.965 142.625 ;
        RECT 106.655 142.020 107.055 151.550 ;
        RECT 107.745 151.035 108.705 151.365 ;
        RECT 109.035 151.035 109.995 151.365 ;
        RECT 107.465 145.785 107.695 150.830 ;
        RECT 108.755 149.485 108.985 150.830 ;
        RECT 108.720 147.185 109.020 149.485 ;
        RECT 107.430 143.485 107.730 145.785 ;
        RECT 107.465 142.830 107.695 143.485 ;
        RECT 108.755 142.830 108.985 147.185 ;
        RECT 110.045 145.785 110.275 150.830 ;
        RECT 110.010 143.485 110.310 145.785 ;
        RECT 110.045 142.830 110.275 143.485 ;
        RECT 107.745 142.395 108.705 142.625 ;
        RECT 109.035 142.395 109.995 142.625 ;
        RECT 110.685 142.020 116.575 151.550 ;
        RECT 117.160 142.145 119.265 155.605 ;
        RECT 122.405 146.245 124.510 155.605 ;
        RECT 125.090 146.825 127.195 155.605 ;
        RECT 130.335 146.825 132.440 155.605 ;
        RECT 133.020 154.960 135.125 155.660 ;
        RECT 133.020 152.675 135.125 154.435 ;
        RECT 138.265 153.845 140.370 155.605 ;
        RECT 133.020 151.450 135.125 152.150 ;
        RECT 138.265 151.505 140.370 153.265 ;
        RECT 140.950 152.675 143.055 156.185 ;
        RECT 146.195 152.675 148.300 156.185 ;
        RECT 140.950 151.460 143.055 152.160 ;
        RECT 133.020 150.280 135.125 150.980 ;
        RECT 133.020 149.110 135.125 149.810 ;
        RECT 138.265 149.165 140.370 150.925 ;
        RECT 140.950 149.165 143.055 150.925 ;
        RECT 146.195 150.335 148.300 152.095 ;
        RECT 133.020 146.825 135.125 148.585 ;
        RECT 138.265 146.825 140.370 148.585 ;
        RECT 140.950 146.825 143.055 148.585 ;
        RECT 146.195 147.995 148.300 149.755 ;
        RECT 122.405 142.145 127.195 146.245 ;
        RECT 130.335 142.145 132.440 146.245 ;
        RECT 133.020 142.145 135.125 146.245 ;
        RECT 138.265 142.145 140.370 146.245 ;
        RECT 140.950 144.485 143.055 146.245 ;
        RECT 146.195 145.655 148.300 147.415 ;
        RECT 140.950 143.290 143.055 143.990 ;
        RECT 146.195 143.315 148.300 145.075 ;
        RECT 140.950 142.040 143.055 142.740 ;
        RECT 146.195 142.080 148.300 142.780 ;
        RECT 102.625 141.620 116.575 142.020 ;
        RECT 62.865 130.990 100.480 139.455 ;
        RECT 111.085 141.565 116.575 141.620 ;
        RECT 148.885 141.565 155.900 156.185 ;
        RECT 111.085 137.690 155.900 141.565 ;
        RECT 111.085 130.990 135.120 137.690 ;
        RECT 62.865 127.485 135.120 130.990 ;
        RECT 138.080 134.100 145.960 137.690 ;
        RECT 138.080 130.310 138.670 134.100 ;
        RECT 139.615 133.640 140.315 133.760 ;
        RECT 140.905 133.640 141.605 133.760 ;
        RECT 139.485 133.410 140.445 133.640 ;
        RECT 140.775 133.410 141.735 133.640 ;
        RECT 139.205 132.990 139.435 133.205 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 139.205 131.205 139.435 131.390 ;
        RECT 140.495 130.310 140.725 133.205 ;
        RECT 141.785 132.990 142.015 133.205 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 143.315 132.640 143.545 133.205 ;
        RECT 143.280 131.940 143.580 132.640 ;
        RECT 141.785 131.205 142.015 131.390 ;
        RECT 143.315 131.205 143.545 131.940 ;
        RECT 144.605 131.205 144.835 134.100 ;
        RECT 143.595 130.770 144.555 131.000 ;
        RECT 143.725 130.700 144.425 130.770 ;
        RECT 145.370 130.310 145.960 134.100 ;
        RECT 138.080 129.720 145.960 130.310 ;
        RECT 4.100 124.285 135.120 127.485 ;
        RECT 4.100 44.835 4.900 124.285 ;
        RECT 8.665 123.695 70.175 124.285 ;
        RECT 8.665 122.800 10.615 123.695 ;
        RECT 11.335 123.005 13.295 123.235 ;
        RECT 13.625 123.005 15.585 123.235 ;
        RECT 17.255 123.005 19.215 123.305 ;
        RECT 19.545 123.005 21.505 123.305 ;
        RECT 23.175 123.005 25.135 123.305 ;
        RECT 25.465 123.005 27.425 123.305 ;
        RECT 29.095 123.005 31.055 123.305 ;
        RECT 31.385 123.005 33.345 123.305 ;
        RECT 35.015 123.005 36.975 123.305 ;
        RECT 37.305 123.005 39.265 123.305 ;
        RECT 40.935 123.005 42.895 123.305 ;
        RECT 43.225 123.005 45.185 123.305 ;
        RECT 46.855 123.005 48.815 123.305 ;
        RECT 49.145 123.005 51.105 123.305 ;
        RECT 52.775 123.005 54.735 123.305 ;
        RECT 55.065 123.005 57.025 123.305 ;
        RECT 58.695 123.005 60.655 123.305 ;
        RECT 60.985 123.005 62.945 123.305 ;
        RECT 64.615 123.005 66.575 123.235 ;
        RECT 66.905 123.005 68.865 123.235 ;
        RECT 69.585 122.800 70.175 123.695 ;
        RECT 8.665 117.050 11.285 122.800 ;
        RECT 13.345 117.050 13.575 122.800 ;
        RECT 15.635 117.050 15.865 122.800 ;
        RECT 16.975 117.050 17.205 122.800 ;
        RECT 19.265 122.050 19.495 122.800 ;
        RECT 19.030 120.550 19.730 122.050 ;
        RECT 8.665 115.550 11.520 117.050 ;
        RECT 13.110 115.550 13.810 117.050 ;
        RECT 15.400 115.550 16.100 117.050 ;
        RECT 16.740 115.550 17.440 117.050 ;
        RECT 8.665 114.595 11.285 115.550 ;
        RECT 13.345 114.595 13.575 115.550 ;
        RECT 15.635 114.595 15.865 115.550 ;
        RECT 16.975 114.800 17.205 115.550 ;
        RECT 19.265 114.800 19.495 120.550 ;
        RECT 21.555 117.050 21.785 122.800 ;
        RECT 22.895 117.050 23.125 122.800 ;
        RECT 25.185 119.550 25.415 122.800 ;
        RECT 24.950 118.050 25.650 119.550 ;
        RECT 21.320 115.550 22.020 117.050 ;
        RECT 22.660 115.550 23.360 117.050 ;
        RECT 21.555 114.800 21.785 115.550 ;
        RECT 22.895 114.800 23.125 115.550 ;
        RECT 25.185 114.800 25.415 118.050 ;
        RECT 27.475 117.050 27.705 122.800 ;
        RECT 28.815 117.050 29.045 122.800 ;
        RECT 27.240 115.550 27.940 117.050 ;
        RECT 28.580 115.550 29.280 117.050 ;
        RECT 27.475 114.800 27.705 115.550 ;
        RECT 28.815 114.800 29.045 115.550 ;
        RECT 31.105 114.595 31.335 122.800 ;
        RECT 33.395 117.050 33.625 122.800 ;
        RECT 34.735 117.050 34.965 122.800 ;
        RECT 37.025 122.050 37.255 122.800 ;
        RECT 36.790 120.550 37.490 122.050 ;
        RECT 33.160 115.550 33.860 117.050 ;
        RECT 34.500 115.550 35.200 117.050 ;
        RECT 33.395 114.800 33.625 115.550 ;
        RECT 34.735 114.800 34.965 115.550 ;
        RECT 37.025 114.800 37.255 120.550 ;
        RECT 39.315 117.050 39.545 122.800 ;
        RECT 40.655 117.050 40.885 122.800 ;
        RECT 42.945 122.050 43.175 122.800 ;
        RECT 42.710 120.550 43.410 122.050 ;
        RECT 39.080 115.550 39.780 117.050 ;
        RECT 40.420 115.550 41.120 117.050 ;
        RECT 39.315 114.800 39.545 115.550 ;
        RECT 40.655 114.800 40.885 115.550 ;
        RECT 42.945 114.800 43.175 120.550 ;
        RECT 45.235 117.050 45.465 122.800 ;
        RECT 46.575 117.050 46.805 122.800 ;
        RECT 45.000 115.550 45.700 117.050 ;
        RECT 46.340 115.550 47.040 117.050 ;
        RECT 45.235 114.800 45.465 115.550 ;
        RECT 46.575 114.800 46.805 115.550 ;
        RECT 48.865 114.595 49.095 122.800 ;
        RECT 51.155 117.050 51.385 122.800 ;
        RECT 52.495 117.050 52.725 122.800 ;
        RECT 54.785 119.550 55.015 122.800 ;
        RECT 54.550 118.050 55.250 119.550 ;
        RECT 50.920 115.550 51.620 117.050 ;
        RECT 52.260 115.550 52.960 117.050 ;
        RECT 51.155 114.800 51.385 115.550 ;
        RECT 52.495 114.800 52.725 115.550 ;
        RECT 54.785 114.800 55.015 118.050 ;
        RECT 57.075 117.050 57.305 122.800 ;
        RECT 58.415 117.050 58.645 122.800 ;
        RECT 60.705 122.050 60.935 122.800 ;
        RECT 60.470 120.550 61.170 122.050 ;
        RECT 56.840 115.550 57.540 117.050 ;
        RECT 58.180 115.550 58.880 117.050 ;
        RECT 57.075 114.800 57.305 115.550 ;
        RECT 58.415 114.800 58.645 115.550 ;
        RECT 60.705 114.800 60.935 120.550 ;
        RECT 62.995 117.050 63.225 122.800 ;
        RECT 64.335 117.050 64.565 122.800 ;
        RECT 66.625 117.050 66.855 122.800 ;
        RECT 68.915 117.050 70.175 122.800 ;
        RECT 62.760 115.550 63.460 117.050 ;
        RECT 64.100 115.550 64.800 117.050 ;
        RECT 66.390 115.550 67.090 117.050 ;
        RECT 68.680 115.550 70.175 117.050 ;
        RECT 62.995 114.800 63.225 115.550 ;
        RECT 64.335 114.595 64.565 115.550 ;
        RECT 66.625 114.595 66.855 115.550 ;
        RECT 68.915 114.595 70.175 115.550 ;
        RECT 8.665 114.365 15.865 114.595 ;
        RECT 8.665 113.215 10.615 114.365 ;
        RECT 17.255 114.295 19.215 114.595 ;
        RECT 19.545 114.295 21.505 114.595 ;
        RECT 23.175 114.295 25.135 114.595 ;
        RECT 25.465 114.295 27.425 114.595 ;
        RECT 29.095 114.365 33.345 114.595 ;
        RECT 29.095 114.295 31.055 114.365 ;
        RECT 31.385 114.295 33.345 114.365 ;
        RECT 35.015 114.295 36.975 114.595 ;
        RECT 37.305 114.295 39.265 114.595 ;
        RECT 40.935 114.295 42.895 114.595 ;
        RECT 43.225 114.295 45.185 114.595 ;
        RECT 46.855 114.365 51.105 114.595 ;
        RECT 46.855 114.295 48.815 114.365 ;
        RECT 49.145 114.295 51.105 114.365 ;
        RECT 52.775 114.295 54.735 114.595 ;
        RECT 55.065 114.295 57.025 114.595 ;
        RECT 58.695 114.295 60.655 114.595 ;
        RECT 60.985 114.295 62.945 114.595 ;
        RECT 64.335 114.365 70.175 114.595 ;
        RECT 8.665 112.985 15.865 113.215 ;
        RECT 17.255 112.985 19.215 113.285 ;
        RECT 19.545 112.985 21.505 113.285 ;
        RECT 23.175 112.985 25.135 113.285 ;
        RECT 25.465 112.985 27.425 113.285 ;
        RECT 29.095 113.215 31.055 113.285 ;
        RECT 31.385 113.215 33.345 113.285 ;
        RECT 29.095 112.985 33.345 113.215 ;
        RECT 35.015 112.985 36.975 113.285 ;
        RECT 37.305 112.985 39.265 113.285 ;
        RECT 40.935 112.985 42.895 113.285 ;
        RECT 43.225 112.985 45.185 113.285 ;
        RECT 46.855 113.215 48.815 113.285 ;
        RECT 49.145 113.215 51.105 113.285 ;
        RECT 46.855 112.985 51.105 113.215 ;
        RECT 52.775 112.985 54.735 113.285 ;
        RECT 55.065 112.985 57.025 113.285 ;
        RECT 58.695 112.985 60.655 113.285 ;
        RECT 60.985 112.985 62.945 113.285 ;
        RECT 69.585 113.215 70.175 114.365 ;
        RECT 64.335 112.985 70.175 113.215 ;
        RECT 8.665 112.030 11.285 112.985 ;
        RECT 13.345 112.030 13.575 112.985 ;
        RECT 15.635 112.030 15.865 112.985 ;
        RECT 16.975 112.030 17.205 112.780 ;
        RECT 8.665 110.530 11.520 112.030 ;
        RECT 13.110 110.530 13.810 112.030 ;
        RECT 15.400 110.530 16.100 112.030 ;
        RECT 16.740 110.530 17.440 112.030 ;
        RECT 8.665 104.780 11.285 110.530 ;
        RECT 13.345 104.780 13.575 110.530 ;
        RECT 15.635 104.780 15.865 110.530 ;
        RECT 16.975 104.780 17.205 110.530 ;
        RECT 19.265 107.030 19.495 112.780 ;
        RECT 21.555 112.030 21.785 112.780 ;
        RECT 22.895 112.030 23.125 112.780 ;
        RECT 21.320 110.530 22.020 112.030 ;
        RECT 22.660 110.530 23.360 112.030 ;
        RECT 19.030 105.530 19.730 107.030 ;
        RECT 19.265 104.780 19.495 105.530 ;
        RECT 21.555 104.780 21.785 110.530 ;
        RECT 22.895 104.780 23.125 110.530 ;
        RECT 25.185 109.530 25.415 112.780 ;
        RECT 27.475 112.030 27.705 112.780 ;
        RECT 28.815 112.030 29.045 112.780 ;
        RECT 27.240 110.530 27.940 112.030 ;
        RECT 28.580 110.530 29.280 112.030 ;
        RECT 24.950 108.030 25.650 109.530 ;
        RECT 25.185 104.780 25.415 108.030 ;
        RECT 27.475 104.780 27.705 110.530 ;
        RECT 28.815 104.780 29.045 110.530 ;
        RECT 31.105 104.780 31.335 112.985 ;
        RECT 33.395 112.030 33.625 112.780 ;
        RECT 34.735 112.030 34.965 112.780 ;
        RECT 33.160 110.530 33.860 112.030 ;
        RECT 34.500 110.530 35.200 112.030 ;
        RECT 33.395 104.780 33.625 110.530 ;
        RECT 34.735 104.780 34.965 110.530 ;
        RECT 37.025 107.030 37.255 112.780 ;
        RECT 39.315 112.030 39.545 112.780 ;
        RECT 40.655 112.030 40.885 112.780 ;
        RECT 39.080 110.530 39.780 112.030 ;
        RECT 40.420 110.530 41.120 112.030 ;
        RECT 36.790 105.530 37.490 107.030 ;
        RECT 37.025 104.780 37.255 105.530 ;
        RECT 39.315 104.780 39.545 110.530 ;
        RECT 40.655 104.780 40.885 110.530 ;
        RECT 42.945 107.030 43.175 112.780 ;
        RECT 45.235 112.030 45.465 112.780 ;
        RECT 46.575 112.030 46.805 112.780 ;
        RECT 45.000 110.530 45.700 112.030 ;
        RECT 46.340 110.530 47.040 112.030 ;
        RECT 42.710 105.530 43.410 107.030 ;
        RECT 42.945 104.780 43.175 105.530 ;
        RECT 45.235 104.780 45.465 110.530 ;
        RECT 46.575 104.780 46.805 110.530 ;
        RECT 48.865 104.780 49.095 112.985 ;
        RECT 51.155 112.030 51.385 112.780 ;
        RECT 52.495 112.030 52.725 112.780 ;
        RECT 50.920 110.530 51.620 112.030 ;
        RECT 52.260 110.530 52.960 112.030 ;
        RECT 51.155 104.780 51.385 110.530 ;
        RECT 52.495 104.780 52.725 110.530 ;
        RECT 54.785 109.530 55.015 112.780 ;
        RECT 57.075 112.030 57.305 112.780 ;
        RECT 58.415 112.030 58.645 112.780 ;
        RECT 56.840 110.530 57.540 112.030 ;
        RECT 58.180 110.530 58.880 112.030 ;
        RECT 54.550 108.030 55.250 109.530 ;
        RECT 54.785 104.780 55.015 108.030 ;
        RECT 57.075 104.780 57.305 110.530 ;
        RECT 58.415 104.780 58.645 110.530 ;
        RECT 60.705 107.030 60.935 112.780 ;
        RECT 62.995 112.030 63.225 112.780 ;
        RECT 64.335 112.030 64.565 112.985 ;
        RECT 66.625 112.030 66.855 112.985 ;
        RECT 68.915 112.030 70.175 112.985 ;
        RECT 62.760 110.530 63.460 112.030 ;
        RECT 64.100 110.530 64.800 112.030 ;
        RECT 66.390 110.530 67.090 112.030 ;
        RECT 68.680 110.530 70.175 112.030 ;
        RECT 60.470 105.530 61.170 107.030 ;
        RECT 60.705 104.780 60.935 105.530 ;
        RECT 62.995 104.780 63.225 110.530 ;
        RECT 64.335 104.780 64.565 110.530 ;
        RECT 66.625 104.780 66.855 110.530 ;
        RECT 68.915 104.780 70.175 110.530 ;
        RECT 8.665 103.885 10.615 104.780 ;
        RECT 11.335 104.345 13.295 104.575 ;
        RECT 13.625 104.345 15.585 104.575 ;
        RECT 17.255 104.275 19.215 104.575 ;
        RECT 19.545 104.275 21.505 104.575 ;
        RECT 23.175 104.275 25.135 104.575 ;
        RECT 25.465 104.275 27.425 104.575 ;
        RECT 29.095 104.275 31.055 104.575 ;
        RECT 31.385 104.275 33.345 104.575 ;
        RECT 35.015 104.275 36.975 104.575 ;
        RECT 37.305 104.275 39.265 104.575 ;
        RECT 40.935 104.275 42.895 104.575 ;
        RECT 43.225 104.275 45.185 104.575 ;
        RECT 46.855 104.275 48.815 104.575 ;
        RECT 49.145 104.275 51.105 104.575 ;
        RECT 52.775 104.275 54.735 104.575 ;
        RECT 55.065 104.275 57.025 104.575 ;
        RECT 58.695 104.275 60.655 104.575 ;
        RECT 60.985 104.275 62.945 104.575 ;
        RECT 64.615 104.345 66.575 104.575 ;
        RECT 66.905 104.345 68.865 104.575 ;
        RECT 69.585 103.885 70.175 104.780 ;
        RECT 8.665 102.705 70.175 103.885 ;
        RECT 71.775 123.695 114.165 124.285 ;
        RECT 71.775 103.885 72.365 123.695 ;
        RECT 72.805 122.800 77.615 123.695 ;
        RECT 79.005 123.005 80.965 123.305 ;
        RECT 81.295 123.005 83.255 123.305 ;
        RECT 84.925 123.005 86.885 123.305 ;
        RECT 87.215 123.005 89.175 123.305 ;
        RECT 90.845 123.005 95.095 123.305 ;
        RECT 96.765 123.005 98.725 123.305 ;
        RECT 99.055 123.005 101.015 123.305 ;
        RECT 102.685 123.005 104.645 123.305 ;
        RECT 104.975 123.005 106.935 123.305 ;
        RECT 72.805 114.800 73.035 122.800 ;
        RECT 75.095 114.800 75.325 122.800 ;
        RECT 77.385 114.800 77.615 122.800 ;
        RECT 78.725 120.650 78.955 122.800 ;
        RECT 78.490 119.950 79.190 120.650 ;
        RECT 78.725 114.800 78.955 119.950 ;
        RECT 81.015 119.150 81.245 122.800 ;
        RECT 83.305 120.650 83.535 122.800 ;
        RECT 83.070 119.950 83.770 120.650 ;
        RECT 80.780 118.450 81.480 119.150 ;
        RECT 81.015 114.800 81.245 118.450 ;
        RECT 83.305 114.800 83.535 119.950 ;
        RECT 84.645 116.150 84.875 122.800 ;
        RECT 86.935 117.650 87.165 122.800 ;
        RECT 86.700 116.950 87.400 117.650 ;
        RECT 84.410 115.450 85.110 116.150 ;
        RECT 84.645 114.800 84.875 115.450 ;
        RECT 86.935 114.800 87.165 116.950 ;
        RECT 89.225 116.150 89.455 122.800 ;
        RECT 90.565 122.150 90.795 122.800 ;
        RECT 90.330 121.450 91.030 122.150 ;
        RECT 88.990 115.450 89.690 116.150 ;
        RECT 89.225 114.800 89.455 115.450 ;
        RECT 90.565 114.800 90.795 121.450 ;
        RECT 92.855 114.800 93.085 123.005 ;
        RECT 108.325 122.800 113.135 123.695 ;
        RECT 95.145 122.150 95.375 122.800 ;
        RECT 94.910 121.450 95.610 122.150 ;
        RECT 95.145 114.800 95.375 121.450 ;
        RECT 96.485 116.150 96.715 122.800 ;
        RECT 98.775 117.650 99.005 122.800 ;
        RECT 98.540 116.950 99.240 117.650 ;
        RECT 96.250 115.450 96.950 116.150 ;
        RECT 96.485 114.800 96.715 115.450 ;
        RECT 98.775 114.800 99.005 116.950 ;
        RECT 101.065 116.150 101.295 122.800 ;
        RECT 102.405 120.650 102.635 122.800 ;
        RECT 102.170 119.950 102.870 120.650 ;
        RECT 100.830 115.450 101.530 116.150 ;
        RECT 101.065 114.800 101.295 115.450 ;
        RECT 102.405 114.800 102.635 119.950 ;
        RECT 104.695 119.150 104.925 122.800 ;
        RECT 106.985 120.650 107.215 122.800 ;
        RECT 106.750 119.950 107.450 120.650 ;
        RECT 104.460 118.450 105.160 119.150 ;
        RECT 104.695 114.800 104.925 118.450 ;
        RECT 106.985 114.800 107.215 119.950 ;
        RECT 108.325 114.800 108.555 122.800 ;
        RECT 110.615 114.800 110.845 122.800 ;
        RECT 112.905 114.800 113.135 122.800 ;
        RECT 73.085 114.365 75.045 114.595 ;
        RECT 75.375 114.365 77.335 114.595 ;
        RECT 79.005 114.295 80.965 114.595 ;
        RECT 81.295 114.295 83.255 114.595 ;
        RECT 84.925 114.295 86.885 114.595 ;
        RECT 87.215 114.295 89.175 114.595 ;
        RECT 90.845 114.295 92.805 114.595 ;
        RECT 93.135 114.295 95.095 114.595 ;
        RECT 96.765 114.295 98.725 114.595 ;
        RECT 99.055 114.295 101.015 114.595 ;
        RECT 102.685 114.295 104.645 114.595 ;
        RECT 104.975 114.295 106.935 114.595 ;
        RECT 108.605 114.365 110.565 114.595 ;
        RECT 110.895 114.365 112.855 114.595 ;
        RECT 73.085 112.985 75.045 113.215 ;
        RECT 75.375 112.985 77.335 113.215 ;
        RECT 79.005 112.985 80.965 113.285 ;
        RECT 81.295 112.985 83.255 113.285 ;
        RECT 84.925 112.985 86.885 113.285 ;
        RECT 87.215 112.985 89.175 113.285 ;
        RECT 90.845 112.985 92.805 113.285 ;
        RECT 93.135 112.985 95.095 113.285 ;
        RECT 96.765 112.985 98.725 113.285 ;
        RECT 99.055 112.985 101.015 113.285 ;
        RECT 102.685 112.985 104.645 113.285 ;
        RECT 104.975 112.985 106.935 113.285 ;
        RECT 108.605 112.985 110.565 113.215 ;
        RECT 110.895 112.985 112.855 113.215 ;
        RECT 72.805 104.780 73.035 112.780 ;
        RECT 75.095 104.780 75.325 112.780 ;
        RECT 77.385 104.780 77.615 112.780 ;
        RECT 78.725 107.630 78.955 112.780 ;
        RECT 81.015 109.130 81.245 112.780 ;
        RECT 80.780 108.430 81.480 109.130 ;
        RECT 78.490 106.930 79.190 107.630 ;
        RECT 78.725 104.780 78.955 106.930 ;
        RECT 81.015 104.780 81.245 108.430 ;
        RECT 83.305 107.630 83.535 112.780 ;
        RECT 84.645 112.130 84.875 112.780 ;
        RECT 84.410 111.430 85.110 112.130 ;
        RECT 83.070 106.930 83.770 107.630 ;
        RECT 83.305 104.780 83.535 106.930 ;
        RECT 84.645 104.780 84.875 111.430 ;
        RECT 86.935 110.630 87.165 112.780 ;
        RECT 89.225 112.130 89.455 112.780 ;
        RECT 88.990 111.430 89.690 112.130 ;
        RECT 86.700 109.930 87.400 110.630 ;
        RECT 86.935 104.780 87.165 109.930 ;
        RECT 89.225 104.780 89.455 111.430 ;
        RECT 90.565 106.130 90.795 112.780 ;
        RECT 90.330 105.430 91.030 106.130 ;
        RECT 90.565 104.780 90.795 105.430 ;
        RECT 72.805 103.885 77.615 104.780 ;
        RECT 92.855 104.575 93.085 112.780 ;
        RECT 95.145 106.130 95.375 112.780 ;
        RECT 96.485 112.130 96.715 112.780 ;
        RECT 96.250 111.430 96.950 112.130 ;
        RECT 94.910 105.430 95.610 106.130 ;
        RECT 95.145 104.780 95.375 105.430 ;
        RECT 96.485 104.780 96.715 111.430 ;
        RECT 98.775 110.630 99.005 112.780 ;
        RECT 101.065 112.130 101.295 112.780 ;
        RECT 100.830 111.430 101.530 112.130 ;
        RECT 98.540 109.930 99.240 110.630 ;
        RECT 98.775 104.780 99.005 109.930 ;
        RECT 101.065 104.780 101.295 111.430 ;
        RECT 102.405 107.630 102.635 112.780 ;
        RECT 104.695 109.130 104.925 112.780 ;
        RECT 104.460 108.430 105.160 109.130 ;
        RECT 102.170 106.930 102.870 107.630 ;
        RECT 102.405 104.780 102.635 106.930 ;
        RECT 104.695 104.780 104.925 108.430 ;
        RECT 106.985 107.630 107.215 112.780 ;
        RECT 106.750 106.930 107.450 107.630 ;
        RECT 106.985 104.780 107.215 106.930 ;
        RECT 108.325 104.780 108.555 112.780 ;
        RECT 110.615 104.780 110.845 112.780 ;
        RECT 112.905 104.780 113.135 112.780 ;
        RECT 79.005 104.275 80.965 104.575 ;
        RECT 81.295 104.275 83.255 104.575 ;
        RECT 84.925 104.275 86.885 104.575 ;
        RECT 87.215 104.275 89.175 104.575 ;
        RECT 90.845 104.275 95.095 104.575 ;
        RECT 96.765 104.275 98.725 104.575 ;
        RECT 99.055 104.275 101.015 104.575 ;
        RECT 102.685 104.275 104.645 104.575 ;
        RECT 104.975 104.275 106.935 104.575 ;
        RECT 108.325 103.885 113.135 104.780 ;
        RECT 113.575 103.885 114.165 123.695 ;
        RECT 128.935 123.505 135.120 124.285 ;
        RECT 138.080 128.380 145.960 128.970 ;
        RECT 138.080 124.680 138.670 128.380 ;
        RECT 139.205 127.290 139.435 127.530 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.205 125.530 139.435 125.690 ;
        RECT 140.495 125.530 140.725 128.380 ;
        RECT 143.725 127.920 144.425 127.990 ;
        RECT 143.595 127.690 144.555 127.920 ;
        RECT 141.785 127.290 142.015 127.530 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 143.315 126.865 143.545 127.530 ;
        RECT 143.280 126.165 143.580 126.865 ;
        RECT 141.785 125.530 142.015 125.690 ;
        RECT 143.315 125.370 143.545 126.165 ;
        RECT 139.390 125.140 143.545 125.370 ;
        RECT 144.605 124.680 144.835 127.530 ;
        RECT 145.370 124.680 145.960 128.380 ;
        RECT 138.080 124.090 145.960 124.680 ;
        RECT 71.775 102.705 114.165 103.885 ;
        RECT 115.905 122.915 135.120 123.505 ;
        RECT 115.905 122.475 116.495 122.915 ;
        RECT 115.905 122.245 118.390 122.475 ;
        RECT 115.905 114.185 117.185 122.245 ;
        RECT 118.595 114.235 118.825 122.195 ;
        RECT 119.975 118.645 120.205 122.195 ;
        RECT 120.410 122.010 121.410 122.710 ;
        RECT 121.615 118.645 121.845 122.195 ;
        RECT 119.975 117.075 121.845 118.645 ;
        RECT 115.905 113.955 118.390 114.185 ;
        RECT 115.905 112.845 116.495 113.955 ;
        RECT 115.905 112.615 118.390 112.845 ;
        RECT 115.905 104.555 117.185 112.615 ;
        RECT 118.595 104.605 118.825 112.565 ;
        RECT 119.975 109.685 120.205 117.075 ;
        RECT 121.615 114.235 121.845 117.075 ;
        RECT 122.995 118.645 123.225 122.195 ;
        RECT 123.430 122.010 124.430 122.710 ;
        RECT 128.345 122.475 135.120 122.915 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 126.450 122.245 135.120 122.475 ;
        RECT 124.635 118.645 124.865 122.195 ;
        RECT 122.995 117.075 124.865 118.645 ;
        RECT 122.995 114.235 123.225 117.075 ;
        RECT 120.410 112.615 121.410 114.185 ;
        RECT 123.430 112.615 124.430 114.185 ;
        RECT 121.615 109.685 121.845 112.565 ;
        RECT 119.975 108.115 121.845 109.685 ;
        RECT 119.975 104.605 120.205 108.115 ;
        RECT 115.905 104.325 118.390 104.555 ;
        RECT 115.905 103.885 116.495 104.325 ;
        RECT 120.410 104.090 121.410 104.790 ;
        RECT 121.615 104.605 121.845 108.115 ;
        RECT 122.995 109.685 123.225 112.565 ;
        RECT 124.635 109.685 124.865 117.075 ;
        RECT 126.015 114.235 126.245 122.195 ;
        RECT 127.655 114.185 135.120 122.245 ;
        RECT 126.450 113.955 135.120 114.185 ;
        RECT 128.345 112.845 135.120 113.955 ;
        RECT 126.450 112.615 135.120 112.845 ;
        RECT 122.995 108.115 124.865 109.685 ;
        RECT 122.995 104.605 123.225 108.115 ;
        RECT 123.430 104.090 124.430 104.790 ;
        RECT 124.635 104.605 124.865 108.115 ;
        RECT 126.015 104.605 126.245 112.565 ;
        RECT 127.655 107.765 135.120 112.615 ;
        RECT 136.295 108.925 142.995 109.515 ;
        RECT 127.655 104.835 138.400 107.765 ;
        RECT 127.655 104.555 135.710 104.835 ;
        RECT 126.450 104.325 135.710 104.555 ;
        RECT 128.345 103.885 135.710 104.325 ;
        RECT 115.905 102.705 135.710 103.885 ;
        RECT 8.665 102.115 135.710 102.705 ;
        RECT 136.295 102.495 138.400 104.255 ;
        RECT 8.665 44.835 10.615 102.115 ;
        RECT 4.100 42.225 10.615 44.835 ;
        RECT 11.055 101.425 29.605 102.115 ;
        RECT 11.055 93.015 11.285 101.425 ;
        RECT 13.345 93.015 13.575 101.425 ;
        RECT 15.635 93.015 15.865 101.425 ;
        RECT 17.925 93.015 18.155 101.425 ;
        RECT 20.215 93.015 20.445 101.425 ;
        RECT 22.505 93.015 22.735 101.425 ;
        RECT 24.795 93.015 25.025 101.425 ;
        RECT 27.085 93.015 27.315 101.425 ;
        RECT 29.375 93.015 29.605 101.425 ;
        RECT 30.715 101.425 49.265 102.115 ;
        RECT 30.715 93.220 30.945 101.425 ;
        RECT 33.005 93.220 33.235 101.425 ;
        RECT 35.295 93.220 35.525 101.425 ;
        RECT 37.585 93.220 37.815 101.425 ;
        RECT 39.875 93.220 40.105 101.425 ;
        RECT 42.165 93.220 42.395 101.425 ;
        RECT 44.455 93.220 44.685 101.425 ;
        RECT 46.745 93.220 46.975 101.425 ;
        RECT 49.035 93.220 49.265 101.425 ;
        RECT 50.375 101.425 68.925 102.115 ;
        RECT 50.375 93.220 50.605 101.425 ;
        RECT 52.665 93.220 52.895 101.425 ;
        RECT 54.955 93.220 55.185 101.425 ;
        RECT 57.245 93.220 57.475 101.425 ;
        RECT 59.535 93.220 59.765 101.425 ;
        RECT 61.825 93.220 62.055 101.425 ;
        RECT 64.115 93.220 64.345 101.425 ;
        RECT 66.405 93.220 66.635 101.425 ;
        RECT 68.695 93.220 68.925 101.425 ;
        RECT 70.035 101.425 88.585 102.115 ;
        RECT 70.035 93.220 70.265 101.425 ;
        RECT 72.325 93.220 72.555 101.425 ;
        RECT 74.615 93.220 74.845 101.425 ;
        RECT 76.905 93.220 77.135 101.425 ;
        RECT 79.195 93.220 79.425 101.425 ;
        RECT 81.485 93.220 81.715 101.425 ;
        RECT 83.775 93.220 84.005 101.425 ;
        RECT 86.065 93.220 86.295 101.425 ;
        RECT 88.355 93.220 88.585 101.425 ;
        RECT 89.695 101.425 108.245 102.115 ;
        RECT 89.695 93.220 89.925 101.425 ;
        RECT 91.985 93.220 92.215 101.425 ;
        RECT 94.275 93.220 94.505 101.425 ;
        RECT 96.565 93.220 96.795 101.425 ;
        RECT 98.855 93.220 99.085 101.425 ;
        RECT 101.145 93.220 101.375 101.425 ;
        RECT 103.435 93.220 103.665 101.425 ;
        RECT 105.725 93.220 105.955 101.425 ;
        RECT 108.015 93.220 108.245 101.425 ;
        RECT 109.355 101.425 127.905 102.115 ;
        RECT 109.355 93.015 109.585 101.425 ;
        RECT 111.645 93.015 111.875 101.425 ;
        RECT 113.935 93.015 114.165 101.425 ;
        RECT 116.225 93.015 116.455 101.425 ;
        RECT 118.515 93.015 118.745 101.425 ;
        RECT 120.805 93.015 121.035 101.425 ;
        RECT 123.095 93.015 123.325 101.425 ;
        RECT 125.385 93.015 125.615 101.425 ;
        RECT 127.675 93.015 127.905 101.425 ;
        RECT 11.055 91.405 29.605 93.015 ;
        RECT 30.995 92.785 32.955 93.015 ;
        RECT 33.285 92.785 35.245 93.015 ;
        RECT 35.575 92.785 37.535 93.015 ;
        RECT 37.865 92.785 39.825 93.015 ;
        RECT 40.155 92.785 42.115 93.015 ;
        RECT 42.445 92.785 44.405 93.015 ;
        RECT 44.735 92.785 46.695 93.015 ;
        RECT 47.025 92.785 48.985 93.015 ;
        RECT 50.655 92.785 52.615 93.015 ;
        RECT 52.945 92.785 54.905 93.015 ;
        RECT 55.235 92.785 57.195 93.015 ;
        RECT 57.525 92.785 59.485 93.015 ;
        RECT 59.815 92.785 61.775 93.015 ;
        RECT 62.105 92.785 64.065 93.015 ;
        RECT 64.395 92.785 66.355 93.015 ;
        RECT 66.685 92.785 68.645 93.015 ;
        RECT 70.315 92.785 72.275 93.015 ;
        RECT 72.605 92.785 74.565 93.015 ;
        RECT 74.895 92.785 76.855 93.015 ;
        RECT 77.185 92.785 79.145 93.015 ;
        RECT 79.475 92.785 81.435 93.015 ;
        RECT 81.765 92.785 83.725 93.015 ;
        RECT 84.055 92.785 86.015 93.015 ;
        RECT 86.345 92.785 88.305 93.015 ;
        RECT 89.975 92.785 91.935 93.015 ;
        RECT 92.265 92.785 94.225 93.015 ;
        RECT 94.555 92.785 96.515 93.015 ;
        RECT 96.845 92.785 98.805 93.015 ;
        RECT 99.135 92.785 101.095 93.015 ;
        RECT 101.425 92.785 103.385 93.015 ;
        RECT 103.715 92.785 105.675 93.015 ;
        RECT 106.005 92.785 107.965 93.015 ;
        RECT 30.995 91.405 32.955 91.635 ;
        RECT 11.055 82.995 11.285 91.405 ;
        RECT 13.345 82.995 13.575 91.405 ;
        RECT 15.635 82.995 15.865 91.405 ;
        RECT 17.925 82.995 18.155 91.405 ;
        RECT 20.215 82.995 20.445 91.405 ;
        RECT 22.505 82.995 22.735 91.405 ;
        RECT 24.795 82.995 25.025 91.405 ;
        RECT 27.085 82.995 27.315 91.405 ;
        RECT 29.375 82.995 29.605 91.405 ;
        RECT 33.285 91.345 35.245 91.875 ;
        RECT 35.575 91.345 37.535 91.875 ;
        RECT 37.865 91.405 39.825 91.635 ;
        RECT 40.155 91.405 42.115 91.635 ;
        RECT 42.445 91.345 44.405 91.875 ;
        RECT 44.735 91.345 46.695 91.875 ;
        RECT 47.025 91.405 48.985 91.635 ;
        RECT 50.655 91.345 52.615 91.875 ;
        RECT 52.945 91.405 54.905 91.635 ;
        RECT 55.235 91.405 57.195 91.635 ;
        RECT 57.525 91.345 59.485 91.875 ;
        RECT 59.815 91.345 61.775 91.875 ;
        RECT 62.105 91.405 64.065 91.635 ;
        RECT 64.395 91.405 66.355 91.635 ;
        RECT 66.685 91.345 68.645 91.875 ;
        RECT 70.315 91.345 72.275 91.875 ;
        RECT 72.605 91.405 74.565 91.635 ;
        RECT 74.895 91.405 76.855 91.635 ;
        RECT 77.185 91.345 79.145 91.875 ;
        RECT 79.475 91.345 81.435 91.875 ;
        RECT 81.765 91.405 83.725 91.635 ;
        RECT 84.055 91.405 86.015 91.635 ;
        RECT 86.345 91.345 88.305 91.875 ;
        RECT 89.975 91.405 91.935 91.635 ;
        RECT 92.265 91.345 94.225 91.875 ;
        RECT 94.555 91.345 96.515 91.875 ;
        RECT 96.845 91.405 98.805 91.635 ;
        RECT 99.135 91.405 101.095 91.635 ;
        RECT 101.425 91.345 103.385 91.875 ;
        RECT 103.715 91.345 105.675 91.875 ;
        RECT 106.005 91.405 107.965 91.635 ;
        RECT 109.355 91.405 127.905 93.015 ;
        RECT 30.715 84.590 30.945 91.200 ;
        RECT 33.005 88.540 33.235 91.200 ;
        RECT 35.295 91.090 35.525 91.200 ;
        RECT 35.260 89.690 35.560 91.090 ;
        RECT 32.970 85.740 33.270 88.540 ;
        RECT 30.680 83.190 30.980 84.590 ;
        RECT 33.005 83.200 33.235 85.740 ;
        RECT 35.295 83.200 35.525 89.690 ;
        RECT 37.585 88.540 37.815 91.200 ;
        RECT 37.550 85.740 37.850 88.540 ;
        RECT 37.585 83.200 37.815 85.740 ;
        RECT 39.875 84.590 40.105 91.200 ;
        RECT 42.165 88.540 42.395 91.200 ;
        RECT 44.455 91.090 44.685 91.200 ;
        RECT 44.420 89.690 44.720 91.090 ;
        RECT 42.130 85.740 42.430 88.540 ;
        RECT 39.840 83.190 40.140 84.590 ;
        RECT 42.165 83.200 42.395 85.740 ;
        RECT 44.455 83.200 44.685 89.690 ;
        RECT 46.745 88.540 46.975 91.200 ;
        RECT 46.710 85.740 47.010 88.540 ;
        RECT 46.745 83.200 46.975 85.740 ;
        RECT 49.035 84.590 49.265 91.200 ;
        RECT 50.375 91.090 50.605 91.200 ;
        RECT 50.340 89.690 50.640 91.090 ;
        RECT 49.000 83.190 49.300 84.590 ;
        RECT 50.375 83.200 50.605 89.690 ;
        RECT 52.665 88.540 52.895 91.200 ;
        RECT 52.630 85.740 52.930 88.540 ;
        RECT 52.665 83.200 52.895 85.740 ;
        RECT 54.955 84.590 55.185 91.200 ;
        RECT 57.245 88.540 57.475 91.200 ;
        RECT 59.535 91.090 59.765 91.200 ;
        RECT 59.500 89.690 59.800 91.090 ;
        RECT 57.210 85.740 57.510 88.540 ;
        RECT 54.920 83.190 55.220 84.590 ;
        RECT 57.245 83.200 57.475 85.740 ;
        RECT 59.535 83.200 59.765 89.690 ;
        RECT 61.825 88.540 62.055 91.200 ;
        RECT 61.790 85.740 62.090 88.540 ;
        RECT 61.825 83.200 62.055 85.740 ;
        RECT 64.115 84.590 64.345 91.200 ;
        RECT 66.405 88.540 66.635 91.200 ;
        RECT 68.695 91.090 68.925 91.200 ;
        RECT 70.035 91.090 70.265 91.200 ;
        RECT 68.660 89.690 68.960 91.090 ;
        RECT 70.000 89.690 70.300 91.090 ;
        RECT 66.370 85.740 66.670 88.540 ;
        RECT 64.080 83.190 64.380 84.590 ;
        RECT 66.405 83.200 66.635 85.740 ;
        RECT 68.695 83.200 68.925 89.690 ;
        RECT 70.035 83.200 70.265 89.690 ;
        RECT 72.325 88.540 72.555 91.200 ;
        RECT 72.290 85.740 72.590 88.540 ;
        RECT 72.325 83.200 72.555 85.740 ;
        RECT 74.615 84.590 74.845 91.200 ;
        RECT 76.905 88.540 77.135 91.200 ;
        RECT 79.195 91.090 79.425 91.200 ;
        RECT 79.160 89.690 79.460 91.090 ;
        RECT 76.870 85.740 77.170 88.540 ;
        RECT 74.580 83.190 74.880 84.590 ;
        RECT 76.905 83.200 77.135 85.740 ;
        RECT 79.195 83.200 79.425 89.690 ;
        RECT 81.485 88.540 81.715 91.200 ;
        RECT 81.450 85.740 81.750 88.540 ;
        RECT 81.485 83.200 81.715 85.740 ;
        RECT 83.775 84.590 84.005 91.200 ;
        RECT 86.065 88.540 86.295 91.200 ;
        RECT 88.355 91.090 88.585 91.200 ;
        RECT 88.320 89.690 88.620 91.090 ;
        RECT 86.030 85.740 86.330 88.540 ;
        RECT 83.740 83.190 84.040 84.590 ;
        RECT 86.065 83.200 86.295 85.740 ;
        RECT 88.355 83.200 88.585 89.690 ;
        RECT 89.695 84.590 89.925 91.200 ;
        RECT 91.985 88.540 92.215 91.200 ;
        RECT 94.275 91.090 94.505 91.200 ;
        RECT 94.240 89.690 94.540 91.090 ;
        RECT 91.950 85.740 92.250 88.540 ;
        RECT 89.660 83.190 89.960 84.590 ;
        RECT 91.985 83.200 92.215 85.740 ;
        RECT 94.275 83.200 94.505 89.690 ;
        RECT 96.565 88.540 96.795 91.200 ;
        RECT 96.530 85.740 96.830 88.540 ;
        RECT 96.565 83.200 96.795 85.740 ;
        RECT 98.855 84.590 99.085 91.200 ;
        RECT 101.145 88.540 101.375 91.200 ;
        RECT 103.435 91.090 103.665 91.200 ;
        RECT 103.400 89.690 103.700 91.090 ;
        RECT 101.110 85.740 101.410 88.540 ;
        RECT 98.820 83.190 99.120 84.590 ;
        RECT 101.145 83.200 101.375 85.740 ;
        RECT 103.435 83.200 103.665 89.690 ;
        RECT 105.725 88.540 105.955 91.200 ;
        RECT 105.690 85.740 105.990 88.540 ;
        RECT 105.725 83.200 105.955 85.740 ;
        RECT 108.015 84.590 108.245 91.200 ;
        RECT 107.980 83.190 108.280 84.590 ;
        RECT 109.355 82.995 109.585 91.405 ;
        RECT 111.645 82.995 111.875 91.405 ;
        RECT 113.935 82.995 114.165 91.405 ;
        RECT 116.225 82.995 116.455 91.405 ;
        RECT 118.515 82.995 118.745 91.405 ;
        RECT 120.805 82.995 121.035 91.405 ;
        RECT 123.095 82.995 123.325 91.405 ;
        RECT 125.385 82.995 125.615 91.405 ;
        RECT 127.675 82.995 127.905 91.405 ;
        RECT 11.055 81.385 29.605 82.995 ;
        RECT 30.995 82.405 32.955 82.995 ;
        RECT 33.285 82.765 35.245 82.995 ;
        RECT 35.575 82.765 37.535 82.995 ;
        RECT 37.865 82.405 39.825 82.995 ;
        RECT 40.155 82.405 42.115 82.995 ;
        RECT 42.445 82.765 44.405 82.995 ;
        RECT 44.735 82.765 46.695 82.995 ;
        RECT 47.025 82.405 48.985 82.995 ;
        RECT 50.655 82.765 52.615 82.995 ;
        RECT 52.945 82.405 54.905 82.995 ;
        RECT 55.235 82.405 57.195 82.995 ;
        RECT 57.525 82.765 59.485 82.995 ;
        RECT 59.815 82.765 61.775 82.995 ;
        RECT 62.105 82.405 64.065 82.995 ;
        RECT 64.395 82.405 66.355 82.995 ;
        RECT 66.685 82.765 68.645 82.995 ;
        RECT 70.315 82.765 72.275 82.995 ;
        RECT 72.605 82.405 74.565 82.995 ;
        RECT 74.895 82.405 76.855 82.995 ;
        RECT 77.185 82.765 79.145 82.995 ;
        RECT 79.475 82.765 81.435 82.995 ;
        RECT 81.765 82.405 83.725 82.995 ;
        RECT 84.055 82.405 86.015 82.995 ;
        RECT 86.345 82.765 88.305 82.995 ;
        RECT 89.975 82.405 91.935 82.995 ;
        RECT 92.265 82.765 94.225 82.995 ;
        RECT 94.555 82.765 96.515 82.995 ;
        RECT 96.845 82.405 98.805 82.995 ;
        RECT 99.135 82.405 101.095 82.995 ;
        RECT 101.425 82.765 103.385 82.995 ;
        RECT 103.715 82.765 105.675 82.995 ;
        RECT 106.005 82.405 107.965 82.995 ;
        RECT 30.995 81.385 32.955 81.615 ;
        RECT 11.055 72.975 11.285 81.385 ;
        RECT 13.345 72.975 13.575 81.385 ;
        RECT 15.635 72.975 15.865 81.385 ;
        RECT 17.925 72.975 18.155 81.385 ;
        RECT 20.215 72.975 20.445 81.385 ;
        RECT 22.505 72.975 22.735 81.385 ;
        RECT 24.795 72.975 25.025 81.385 ;
        RECT 27.085 72.975 27.315 81.385 ;
        RECT 29.375 72.975 29.605 81.385 ;
        RECT 33.285 81.325 35.245 81.855 ;
        RECT 35.575 81.325 37.535 81.855 ;
        RECT 37.865 81.385 39.825 81.615 ;
        RECT 40.155 81.385 42.115 81.615 ;
        RECT 42.445 81.325 44.405 81.855 ;
        RECT 44.735 81.325 46.695 81.855 ;
        RECT 47.025 81.385 48.985 81.615 ;
        RECT 50.655 81.325 52.615 81.855 ;
        RECT 52.945 81.385 54.905 81.615 ;
        RECT 55.235 81.385 57.195 81.615 ;
        RECT 57.525 81.325 59.485 81.855 ;
        RECT 59.815 81.325 61.775 81.855 ;
        RECT 62.105 81.385 64.065 81.615 ;
        RECT 64.395 81.385 66.355 81.615 ;
        RECT 66.685 81.325 68.645 81.855 ;
        RECT 70.315 81.325 72.275 81.855 ;
        RECT 72.605 81.385 74.565 81.615 ;
        RECT 74.895 81.385 76.855 81.615 ;
        RECT 77.185 81.325 79.145 81.855 ;
        RECT 79.475 81.325 81.435 81.855 ;
        RECT 81.765 81.385 83.725 81.615 ;
        RECT 84.055 81.385 86.015 81.615 ;
        RECT 86.345 81.325 88.305 81.855 ;
        RECT 89.975 81.385 91.935 81.615 ;
        RECT 92.265 81.325 94.225 81.855 ;
        RECT 94.555 81.325 96.515 81.855 ;
        RECT 96.845 81.385 98.805 81.615 ;
        RECT 99.135 81.385 101.095 81.615 ;
        RECT 101.425 81.325 103.385 81.855 ;
        RECT 103.715 81.325 105.675 81.855 ;
        RECT 106.005 81.385 107.965 81.615 ;
        RECT 109.355 81.385 127.905 82.995 ;
        RECT 30.715 81.070 30.945 81.180 ;
        RECT 30.680 79.670 30.980 81.070 ;
        RECT 30.715 73.180 30.945 79.670 ;
        RECT 33.005 78.520 33.235 81.180 ;
        RECT 32.970 75.720 33.270 78.520 ;
        RECT 33.005 73.180 33.235 75.720 ;
        RECT 35.295 74.570 35.525 81.180 ;
        RECT 37.585 78.520 37.815 81.180 ;
        RECT 39.875 81.070 40.105 81.180 ;
        RECT 39.840 79.670 40.140 81.070 ;
        RECT 37.550 75.720 37.850 78.520 ;
        RECT 35.260 73.170 35.560 74.570 ;
        RECT 37.585 73.180 37.815 75.720 ;
        RECT 39.875 73.180 40.105 79.670 ;
        RECT 42.165 78.520 42.395 81.180 ;
        RECT 42.130 75.720 42.430 78.520 ;
        RECT 42.165 73.180 42.395 75.720 ;
        RECT 44.455 74.570 44.685 81.180 ;
        RECT 46.745 78.520 46.975 81.180 ;
        RECT 49.035 81.070 49.265 81.180 ;
        RECT 49.000 79.670 49.300 81.070 ;
        RECT 46.710 75.720 47.010 78.520 ;
        RECT 44.420 73.170 44.720 74.570 ;
        RECT 46.745 73.180 46.975 75.720 ;
        RECT 49.035 73.180 49.265 79.670 ;
        RECT 50.375 74.570 50.605 81.180 ;
        RECT 52.665 78.520 52.895 81.180 ;
        RECT 54.955 81.070 55.185 81.180 ;
        RECT 54.920 79.670 55.220 81.070 ;
        RECT 52.630 75.720 52.930 78.520 ;
        RECT 50.340 73.170 50.640 74.570 ;
        RECT 52.665 73.180 52.895 75.720 ;
        RECT 54.955 73.180 55.185 79.670 ;
        RECT 57.245 78.520 57.475 81.180 ;
        RECT 57.210 75.720 57.510 78.520 ;
        RECT 57.245 73.180 57.475 75.720 ;
        RECT 59.535 74.570 59.765 81.180 ;
        RECT 61.825 78.520 62.055 81.180 ;
        RECT 64.115 81.070 64.345 81.180 ;
        RECT 64.080 79.670 64.380 81.070 ;
        RECT 61.790 75.720 62.090 78.520 ;
        RECT 59.500 73.170 59.800 74.570 ;
        RECT 61.825 73.180 62.055 75.720 ;
        RECT 64.115 73.180 64.345 79.670 ;
        RECT 66.405 78.520 66.635 81.180 ;
        RECT 66.370 75.720 66.670 78.520 ;
        RECT 66.405 73.180 66.635 75.720 ;
        RECT 68.695 74.570 68.925 81.180 ;
        RECT 70.035 74.570 70.265 81.180 ;
        RECT 72.325 78.520 72.555 81.180 ;
        RECT 74.615 81.070 74.845 81.180 ;
        RECT 74.580 79.670 74.880 81.070 ;
        RECT 72.290 75.720 72.590 78.520 ;
        RECT 68.660 73.170 68.960 74.570 ;
        RECT 70.000 73.170 70.300 74.570 ;
        RECT 72.325 73.180 72.555 75.720 ;
        RECT 74.615 73.180 74.845 79.670 ;
        RECT 76.905 78.520 77.135 81.180 ;
        RECT 76.870 75.720 77.170 78.520 ;
        RECT 76.905 73.180 77.135 75.720 ;
        RECT 79.195 74.570 79.425 81.180 ;
        RECT 81.485 78.520 81.715 81.180 ;
        RECT 83.775 81.070 84.005 81.180 ;
        RECT 83.740 79.670 84.040 81.070 ;
        RECT 81.450 75.720 81.750 78.520 ;
        RECT 79.160 73.170 79.460 74.570 ;
        RECT 81.485 73.180 81.715 75.720 ;
        RECT 83.775 73.180 84.005 79.670 ;
        RECT 86.065 78.520 86.295 81.180 ;
        RECT 86.030 75.720 86.330 78.520 ;
        RECT 86.065 73.180 86.295 75.720 ;
        RECT 88.355 74.570 88.585 81.180 ;
        RECT 89.695 81.070 89.925 81.180 ;
        RECT 89.660 79.670 89.960 81.070 ;
        RECT 88.320 73.170 88.620 74.570 ;
        RECT 89.695 73.180 89.925 79.670 ;
        RECT 91.985 78.520 92.215 81.180 ;
        RECT 91.950 75.720 92.250 78.520 ;
        RECT 91.985 73.180 92.215 75.720 ;
        RECT 94.275 74.570 94.505 81.180 ;
        RECT 96.565 78.520 96.795 81.180 ;
        RECT 98.855 81.070 99.085 81.180 ;
        RECT 98.820 79.670 99.120 81.070 ;
        RECT 96.530 75.720 96.830 78.520 ;
        RECT 94.240 73.170 94.540 74.570 ;
        RECT 96.565 73.180 96.795 75.720 ;
        RECT 98.855 73.180 99.085 79.670 ;
        RECT 101.145 78.520 101.375 81.180 ;
        RECT 101.110 75.720 101.410 78.520 ;
        RECT 101.145 73.180 101.375 75.720 ;
        RECT 103.435 74.570 103.665 81.180 ;
        RECT 105.725 78.520 105.955 81.180 ;
        RECT 108.015 81.070 108.245 81.180 ;
        RECT 107.980 79.670 108.280 81.070 ;
        RECT 105.690 75.720 105.990 78.520 ;
        RECT 103.400 73.170 103.700 74.570 ;
        RECT 105.725 73.180 105.955 75.720 ;
        RECT 108.015 73.180 108.245 79.670 ;
        RECT 109.355 72.975 109.585 81.385 ;
        RECT 111.645 72.975 111.875 81.385 ;
        RECT 113.935 72.975 114.165 81.385 ;
        RECT 116.225 72.975 116.455 81.385 ;
        RECT 118.515 72.975 118.745 81.385 ;
        RECT 120.805 72.975 121.035 81.385 ;
        RECT 123.095 72.975 123.325 81.385 ;
        RECT 125.385 72.975 125.615 81.385 ;
        RECT 127.675 72.975 127.905 81.385 ;
        RECT 11.055 71.365 29.605 72.975 ;
        RECT 30.995 72.385 32.955 72.975 ;
        RECT 33.285 72.745 35.245 72.975 ;
        RECT 35.575 72.745 37.535 72.975 ;
        RECT 37.865 72.385 39.825 72.975 ;
        RECT 40.155 72.385 42.115 72.975 ;
        RECT 42.445 72.745 44.405 72.975 ;
        RECT 44.735 72.745 46.695 72.975 ;
        RECT 47.025 72.385 48.985 72.975 ;
        RECT 50.655 72.745 52.615 72.975 ;
        RECT 52.945 72.385 54.905 72.975 ;
        RECT 55.235 72.385 57.195 72.975 ;
        RECT 57.525 72.745 59.485 72.975 ;
        RECT 59.815 72.745 61.775 72.975 ;
        RECT 62.105 72.385 64.065 72.975 ;
        RECT 64.395 72.385 66.355 72.975 ;
        RECT 66.685 72.745 68.645 72.975 ;
        RECT 70.315 72.745 72.275 72.975 ;
        RECT 72.605 72.385 74.565 72.975 ;
        RECT 74.895 72.385 76.855 72.975 ;
        RECT 77.185 72.745 79.145 72.975 ;
        RECT 79.475 72.745 81.435 72.975 ;
        RECT 81.765 72.385 83.725 72.975 ;
        RECT 84.055 72.385 86.015 72.975 ;
        RECT 86.345 72.745 88.305 72.975 ;
        RECT 89.975 72.385 91.935 72.975 ;
        RECT 92.265 72.745 94.225 72.975 ;
        RECT 94.555 72.745 96.515 72.975 ;
        RECT 96.845 72.385 98.805 72.975 ;
        RECT 99.135 72.385 101.095 72.975 ;
        RECT 101.425 72.745 103.385 72.975 ;
        RECT 103.715 72.745 105.675 72.975 ;
        RECT 106.005 72.385 107.965 72.975 ;
        RECT 11.055 62.955 11.285 71.365 ;
        RECT 13.345 62.955 13.575 71.365 ;
        RECT 15.635 62.955 15.865 71.365 ;
        RECT 17.925 62.955 18.155 71.365 ;
        RECT 20.215 62.955 20.445 71.365 ;
        RECT 22.505 62.955 22.735 71.365 ;
        RECT 24.795 62.955 25.025 71.365 ;
        RECT 27.085 62.955 27.315 71.365 ;
        RECT 29.375 62.955 29.605 71.365 ;
        RECT 30.995 71.305 32.955 71.835 ;
        RECT 33.285 71.365 35.245 71.595 ;
        RECT 35.575 71.365 37.535 71.595 ;
        RECT 37.865 71.305 39.825 71.835 ;
        RECT 40.155 71.305 42.115 71.835 ;
        RECT 42.445 71.365 44.405 71.595 ;
        RECT 44.735 71.365 46.695 71.595 ;
        RECT 47.025 71.305 48.985 71.835 ;
        RECT 50.655 71.365 52.615 71.595 ;
        RECT 52.945 71.305 54.905 71.835 ;
        RECT 55.235 71.305 57.195 71.835 ;
        RECT 57.525 71.365 59.485 71.595 ;
        RECT 59.815 71.365 61.775 71.595 ;
        RECT 62.105 71.305 64.065 71.835 ;
        RECT 64.395 71.305 66.355 71.835 ;
        RECT 66.685 71.365 68.645 71.595 ;
        RECT 70.315 71.365 72.275 71.595 ;
        RECT 72.605 71.305 74.565 71.835 ;
        RECT 74.895 71.305 76.855 71.835 ;
        RECT 77.185 71.365 79.145 71.595 ;
        RECT 79.475 71.365 81.435 71.595 ;
        RECT 81.765 71.305 83.725 71.835 ;
        RECT 84.055 71.305 86.015 71.835 ;
        RECT 86.345 71.365 88.305 71.595 ;
        RECT 89.975 71.305 91.935 71.835 ;
        RECT 92.265 71.365 94.225 71.595 ;
        RECT 94.555 71.365 96.515 71.595 ;
        RECT 96.845 71.305 98.805 71.835 ;
        RECT 99.135 71.305 101.095 71.835 ;
        RECT 101.425 71.365 103.385 71.595 ;
        RECT 103.715 71.365 105.675 71.595 ;
        RECT 106.005 71.305 107.965 71.835 ;
        RECT 109.355 71.365 127.905 72.975 ;
        RECT 30.715 71.050 30.945 71.160 ;
        RECT 30.680 69.650 30.980 71.050 ;
        RECT 30.715 63.160 30.945 69.650 ;
        RECT 33.005 68.500 33.235 71.160 ;
        RECT 32.970 65.700 33.270 68.500 ;
        RECT 33.005 63.160 33.235 65.700 ;
        RECT 35.295 64.550 35.525 71.160 ;
        RECT 37.585 68.500 37.815 71.160 ;
        RECT 39.875 71.050 40.105 71.160 ;
        RECT 39.840 69.650 40.140 71.050 ;
        RECT 37.550 65.700 37.850 68.500 ;
        RECT 35.260 63.150 35.560 64.550 ;
        RECT 37.585 63.160 37.815 65.700 ;
        RECT 39.875 63.160 40.105 69.650 ;
        RECT 42.165 68.500 42.395 71.160 ;
        RECT 42.130 65.700 42.430 68.500 ;
        RECT 42.165 63.160 42.395 65.700 ;
        RECT 44.455 64.550 44.685 71.160 ;
        RECT 46.745 68.500 46.975 71.160 ;
        RECT 49.035 71.050 49.265 71.160 ;
        RECT 49.000 69.650 49.300 71.050 ;
        RECT 46.710 65.700 47.010 68.500 ;
        RECT 44.420 63.150 44.720 64.550 ;
        RECT 46.745 63.160 46.975 65.700 ;
        RECT 49.035 63.160 49.265 69.650 ;
        RECT 50.375 64.550 50.605 71.160 ;
        RECT 52.665 68.500 52.895 71.160 ;
        RECT 54.955 71.050 55.185 71.160 ;
        RECT 54.920 69.650 55.220 71.050 ;
        RECT 52.630 65.700 52.930 68.500 ;
        RECT 50.340 63.150 50.640 64.550 ;
        RECT 52.665 63.160 52.895 65.700 ;
        RECT 54.955 63.160 55.185 69.650 ;
        RECT 57.245 68.500 57.475 71.160 ;
        RECT 57.210 65.700 57.510 68.500 ;
        RECT 57.245 63.160 57.475 65.700 ;
        RECT 59.535 64.550 59.765 71.160 ;
        RECT 61.825 68.500 62.055 71.160 ;
        RECT 64.115 71.050 64.345 71.160 ;
        RECT 64.080 69.650 64.380 71.050 ;
        RECT 61.790 65.700 62.090 68.500 ;
        RECT 59.500 63.150 59.800 64.550 ;
        RECT 61.825 63.160 62.055 65.700 ;
        RECT 64.115 63.160 64.345 69.650 ;
        RECT 66.405 68.500 66.635 71.160 ;
        RECT 66.370 65.700 66.670 68.500 ;
        RECT 66.405 63.160 66.635 65.700 ;
        RECT 68.695 64.550 68.925 71.160 ;
        RECT 70.035 64.550 70.265 71.160 ;
        RECT 72.325 68.500 72.555 71.160 ;
        RECT 74.615 71.050 74.845 71.160 ;
        RECT 74.580 69.650 74.880 71.050 ;
        RECT 72.290 65.700 72.590 68.500 ;
        RECT 68.660 63.150 68.960 64.550 ;
        RECT 70.000 63.150 70.300 64.550 ;
        RECT 72.325 63.160 72.555 65.700 ;
        RECT 74.615 63.160 74.845 69.650 ;
        RECT 76.905 68.500 77.135 71.160 ;
        RECT 76.870 65.700 77.170 68.500 ;
        RECT 76.905 63.160 77.135 65.700 ;
        RECT 79.195 64.550 79.425 71.160 ;
        RECT 81.485 68.500 81.715 71.160 ;
        RECT 83.775 71.050 84.005 71.160 ;
        RECT 83.740 69.650 84.040 71.050 ;
        RECT 81.450 65.700 81.750 68.500 ;
        RECT 79.160 63.150 79.460 64.550 ;
        RECT 81.485 63.160 81.715 65.700 ;
        RECT 83.775 63.160 84.005 69.650 ;
        RECT 86.065 68.500 86.295 71.160 ;
        RECT 86.030 65.700 86.330 68.500 ;
        RECT 86.065 63.160 86.295 65.700 ;
        RECT 88.355 64.550 88.585 71.160 ;
        RECT 89.695 71.050 89.925 71.160 ;
        RECT 89.660 69.650 89.960 71.050 ;
        RECT 88.320 63.150 88.620 64.550 ;
        RECT 89.695 63.160 89.925 69.650 ;
        RECT 91.985 68.500 92.215 71.160 ;
        RECT 91.950 65.700 92.250 68.500 ;
        RECT 91.985 63.160 92.215 65.700 ;
        RECT 94.275 64.550 94.505 71.160 ;
        RECT 96.565 68.500 96.795 71.160 ;
        RECT 98.855 71.050 99.085 71.160 ;
        RECT 98.820 69.650 99.120 71.050 ;
        RECT 96.530 65.700 96.830 68.500 ;
        RECT 94.240 63.150 94.540 64.550 ;
        RECT 96.565 63.160 96.795 65.700 ;
        RECT 98.855 63.160 99.085 69.650 ;
        RECT 101.145 68.500 101.375 71.160 ;
        RECT 101.110 65.700 101.410 68.500 ;
        RECT 101.145 63.160 101.375 65.700 ;
        RECT 103.435 64.550 103.665 71.160 ;
        RECT 105.725 68.500 105.955 71.160 ;
        RECT 108.015 71.050 108.245 71.160 ;
        RECT 107.980 69.650 108.280 71.050 ;
        RECT 105.690 65.700 105.990 68.500 ;
        RECT 103.400 63.150 103.700 64.550 ;
        RECT 105.725 63.160 105.955 65.700 ;
        RECT 108.015 63.160 108.245 69.650 ;
        RECT 109.355 62.955 109.585 71.365 ;
        RECT 111.645 62.955 111.875 71.365 ;
        RECT 113.935 62.955 114.165 71.365 ;
        RECT 116.225 62.955 116.455 71.365 ;
        RECT 118.515 62.955 118.745 71.365 ;
        RECT 120.805 62.955 121.035 71.365 ;
        RECT 123.095 62.955 123.325 71.365 ;
        RECT 125.385 62.955 125.615 71.365 ;
        RECT 127.675 62.955 127.905 71.365 ;
        RECT 11.055 61.345 29.605 62.955 ;
        RECT 30.995 62.725 32.955 62.955 ;
        RECT 33.285 62.365 35.245 62.955 ;
        RECT 35.575 62.365 37.535 62.955 ;
        RECT 37.865 62.725 39.825 62.955 ;
        RECT 40.155 62.725 42.115 62.955 ;
        RECT 42.445 62.365 44.405 62.955 ;
        RECT 44.735 62.365 46.695 62.955 ;
        RECT 47.025 62.725 48.985 62.955 ;
        RECT 50.655 62.365 52.615 62.955 ;
        RECT 52.945 62.725 54.905 62.955 ;
        RECT 55.235 62.725 57.195 62.955 ;
        RECT 57.525 62.365 59.485 62.955 ;
        RECT 59.815 62.365 61.775 62.955 ;
        RECT 62.105 62.725 64.065 62.955 ;
        RECT 64.395 62.725 66.355 62.955 ;
        RECT 66.685 62.365 68.645 62.955 ;
        RECT 70.315 62.365 72.275 62.955 ;
        RECT 72.605 62.725 74.565 62.955 ;
        RECT 74.895 62.725 76.855 62.955 ;
        RECT 77.185 62.365 79.145 62.955 ;
        RECT 79.475 62.365 81.435 62.955 ;
        RECT 81.765 62.725 83.725 62.955 ;
        RECT 84.055 62.725 86.015 62.955 ;
        RECT 86.345 62.365 88.305 62.955 ;
        RECT 89.975 62.725 91.935 62.955 ;
        RECT 92.265 62.365 94.225 62.955 ;
        RECT 94.555 62.365 96.515 62.955 ;
        RECT 96.845 62.725 98.805 62.955 ;
        RECT 99.135 62.725 101.095 62.955 ;
        RECT 101.425 62.365 103.385 62.955 ;
        RECT 103.715 62.365 105.675 62.955 ;
        RECT 106.005 62.725 107.965 62.955 ;
        RECT 11.055 52.935 11.285 61.345 ;
        RECT 13.345 52.935 13.575 61.345 ;
        RECT 15.635 52.935 15.865 61.345 ;
        RECT 17.925 52.935 18.155 61.345 ;
        RECT 20.215 52.935 20.445 61.345 ;
        RECT 22.505 52.935 22.735 61.345 ;
        RECT 24.795 52.935 25.025 61.345 ;
        RECT 27.085 52.935 27.315 61.345 ;
        RECT 29.375 52.935 29.605 61.345 ;
        RECT 30.995 61.285 32.955 61.815 ;
        RECT 33.285 61.345 35.245 61.575 ;
        RECT 35.575 61.345 37.535 61.575 ;
        RECT 37.865 61.285 39.825 61.815 ;
        RECT 40.155 61.285 42.115 61.815 ;
        RECT 42.445 61.345 44.405 61.575 ;
        RECT 44.735 61.345 46.695 61.575 ;
        RECT 47.025 61.285 48.985 61.815 ;
        RECT 50.655 61.345 52.615 61.575 ;
        RECT 52.945 61.285 54.905 61.815 ;
        RECT 55.235 61.285 57.195 61.815 ;
        RECT 57.525 61.345 59.485 61.575 ;
        RECT 59.815 61.345 61.775 61.575 ;
        RECT 62.105 61.285 64.065 61.815 ;
        RECT 64.395 61.285 66.355 61.815 ;
        RECT 66.685 61.345 68.645 61.575 ;
        RECT 70.315 61.345 72.275 61.575 ;
        RECT 72.605 61.285 74.565 61.815 ;
        RECT 74.895 61.285 76.855 61.815 ;
        RECT 77.185 61.345 79.145 61.575 ;
        RECT 79.475 61.345 81.435 61.575 ;
        RECT 81.765 61.285 83.725 61.815 ;
        RECT 84.055 61.285 86.015 61.815 ;
        RECT 86.345 61.345 88.305 61.575 ;
        RECT 89.975 61.285 91.935 61.815 ;
        RECT 92.265 61.345 94.225 61.575 ;
        RECT 94.555 61.345 96.515 61.575 ;
        RECT 96.845 61.285 98.805 61.815 ;
        RECT 99.135 61.285 101.095 61.815 ;
        RECT 101.425 61.345 103.385 61.575 ;
        RECT 103.715 61.345 105.675 61.575 ;
        RECT 106.005 61.285 107.965 61.815 ;
        RECT 109.355 61.345 127.905 62.955 ;
        RECT 30.715 54.530 30.945 61.140 ;
        RECT 33.005 58.480 33.235 61.140 ;
        RECT 35.295 61.030 35.525 61.140 ;
        RECT 35.260 59.630 35.560 61.030 ;
        RECT 32.970 55.680 33.270 58.480 ;
        RECT 30.680 53.130 30.980 54.530 ;
        RECT 33.005 53.140 33.235 55.680 ;
        RECT 35.295 53.140 35.525 59.630 ;
        RECT 37.585 58.480 37.815 61.140 ;
        RECT 37.550 55.680 37.850 58.480 ;
        RECT 37.585 53.140 37.815 55.680 ;
        RECT 39.875 54.530 40.105 61.140 ;
        RECT 42.165 58.480 42.395 61.140 ;
        RECT 44.455 61.030 44.685 61.140 ;
        RECT 44.420 59.630 44.720 61.030 ;
        RECT 42.130 55.680 42.430 58.480 ;
        RECT 39.840 53.130 40.140 54.530 ;
        RECT 42.165 53.140 42.395 55.680 ;
        RECT 44.455 53.140 44.685 59.630 ;
        RECT 46.745 58.480 46.975 61.140 ;
        RECT 46.710 55.680 47.010 58.480 ;
        RECT 46.745 53.140 46.975 55.680 ;
        RECT 49.035 54.530 49.265 61.140 ;
        RECT 50.375 61.030 50.605 61.140 ;
        RECT 50.340 59.630 50.640 61.030 ;
        RECT 49.000 53.130 49.300 54.530 ;
        RECT 50.375 53.140 50.605 59.630 ;
        RECT 52.665 58.480 52.895 61.140 ;
        RECT 52.630 55.680 52.930 58.480 ;
        RECT 52.665 53.140 52.895 55.680 ;
        RECT 54.955 54.530 55.185 61.140 ;
        RECT 57.245 58.480 57.475 61.140 ;
        RECT 59.535 61.030 59.765 61.140 ;
        RECT 59.500 59.630 59.800 61.030 ;
        RECT 57.210 55.680 57.510 58.480 ;
        RECT 54.920 53.130 55.220 54.530 ;
        RECT 57.245 53.140 57.475 55.680 ;
        RECT 59.535 53.140 59.765 59.630 ;
        RECT 61.825 58.480 62.055 61.140 ;
        RECT 61.790 55.680 62.090 58.480 ;
        RECT 61.825 53.140 62.055 55.680 ;
        RECT 64.115 54.530 64.345 61.140 ;
        RECT 66.405 58.480 66.635 61.140 ;
        RECT 68.695 61.030 68.925 61.140 ;
        RECT 70.035 61.030 70.265 61.140 ;
        RECT 68.660 59.630 68.960 61.030 ;
        RECT 70.000 59.630 70.300 61.030 ;
        RECT 66.370 55.680 66.670 58.480 ;
        RECT 64.080 53.130 64.380 54.530 ;
        RECT 66.405 53.140 66.635 55.680 ;
        RECT 68.695 53.140 68.925 59.630 ;
        RECT 70.035 53.140 70.265 59.630 ;
        RECT 72.325 58.480 72.555 61.140 ;
        RECT 72.290 55.680 72.590 58.480 ;
        RECT 72.325 53.140 72.555 55.680 ;
        RECT 74.615 54.530 74.845 61.140 ;
        RECT 76.905 58.480 77.135 61.140 ;
        RECT 79.195 61.030 79.425 61.140 ;
        RECT 79.160 59.630 79.460 61.030 ;
        RECT 76.870 55.680 77.170 58.480 ;
        RECT 74.580 53.130 74.880 54.530 ;
        RECT 76.905 53.140 77.135 55.680 ;
        RECT 79.195 53.140 79.425 59.630 ;
        RECT 81.485 58.480 81.715 61.140 ;
        RECT 81.450 55.680 81.750 58.480 ;
        RECT 81.485 53.140 81.715 55.680 ;
        RECT 83.775 54.530 84.005 61.140 ;
        RECT 86.065 58.480 86.295 61.140 ;
        RECT 88.355 61.030 88.585 61.140 ;
        RECT 88.320 59.630 88.620 61.030 ;
        RECT 86.030 55.680 86.330 58.480 ;
        RECT 83.740 53.130 84.040 54.530 ;
        RECT 86.065 53.140 86.295 55.680 ;
        RECT 88.355 53.140 88.585 59.630 ;
        RECT 89.695 54.530 89.925 61.140 ;
        RECT 91.985 58.480 92.215 61.140 ;
        RECT 94.275 61.030 94.505 61.140 ;
        RECT 94.240 59.630 94.540 61.030 ;
        RECT 91.950 55.680 92.250 58.480 ;
        RECT 89.660 53.130 89.960 54.530 ;
        RECT 91.985 53.140 92.215 55.680 ;
        RECT 94.275 53.140 94.505 59.630 ;
        RECT 96.565 58.480 96.795 61.140 ;
        RECT 96.530 55.680 96.830 58.480 ;
        RECT 96.565 53.140 96.795 55.680 ;
        RECT 98.855 54.530 99.085 61.140 ;
        RECT 101.145 58.480 101.375 61.140 ;
        RECT 103.435 61.030 103.665 61.140 ;
        RECT 103.400 59.630 103.700 61.030 ;
        RECT 101.110 55.680 101.410 58.480 ;
        RECT 98.820 53.130 99.120 54.530 ;
        RECT 101.145 53.140 101.375 55.680 ;
        RECT 103.435 53.140 103.665 59.630 ;
        RECT 105.725 58.480 105.955 61.140 ;
        RECT 105.690 55.680 105.990 58.480 ;
        RECT 105.725 53.140 105.955 55.680 ;
        RECT 108.015 54.530 108.245 61.140 ;
        RECT 107.980 53.130 108.280 54.530 ;
        RECT 109.355 52.935 109.585 61.345 ;
        RECT 111.645 52.935 111.875 61.345 ;
        RECT 113.935 52.935 114.165 61.345 ;
        RECT 116.225 52.935 116.455 61.345 ;
        RECT 118.515 52.935 118.745 61.345 ;
        RECT 120.805 52.935 121.035 61.345 ;
        RECT 123.095 52.935 123.325 61.345 ;
        RECT 125.385 52.935 125.615 61.345 ;
        RECT 127.675 52.935 127.905 61.345 ;
        RECT 11.055 51.325 29.605 52.935 ;
        RECT 30.995 52.705 32.955 52.935 ;
        RECT 33.285 52.345 35.245 52.935 ;
        RECT 35.575 52.345 37.535 52.935 ;
        RECT 37.865 52.705 39.825 52.935 ;
        RECT 40.155 52.705 42.115 52.935 ;
        RECT 42.445 52.345 44.405 52.935 ;
        RECT 44.735 52.345 46.695 52.935 ;
        RECT 47.025 52.705 48.985 52.935 ;
        RECT 50.655 52.345 52.615 52.935 ;
        RECT 52.945 52.705 54.905 52.935 ;
        RECT 55.235 52.705 57.195 52.935 ;
        RECT 57.525 52.345 59.485 52.935 ;
        RECT 59.815 52.345 61.775 52.935 ;
        RECT 62.105 52.705 64.065 52.935 ;
        RECT 64.395 52.705 66.355 52.935 ;
        RECT 66.685 52.345 68.645 52.935 ;
        RECT 70.315 52.345 72.275 52.935 ;
        RECT 72.605 52.705 74.565 52.935 ;
        RECT 74.895 52.705 76.855 52.935 ;
        RECT 77.185 52.345 79.145 52.935 ;
        RECT 79.475 52.345 81.435 52.935 ;
        RECT 81.765 52.705 83.725 52.935 ;
        RECT 84.055 52.705 86.015 52.935 ;
        RECT 86.345 52.345 88.305 52.935 ;
        RECT 89.975 52.705 91.935 52.935 ;
        RECT 92.265 52.345 94.225 52.935 ;
        RECT 94.555 52.345 96.515 52.935 ;
        RECT 96.845 52.705 98.805 52.935 ;
        RECT 99.135 52.705 101.095 52.935 ;
        RECT 101.425 52.345 103.385 52.935 ;
        RECT 103.715 52.345 105.675 52.935 ;
        RECT 106.005 52.705 107.965 52.935 ;
        RECT 30.995 51.325 32.955 51.555 ;
        RECT 33.285 51.325 35.245 51.555 ;
        RECT 35.575 51.325 37.535 51.555 ;
        RECT 37.865 51.325 39.825 51.555 ;
        RECT 40.155 51.325 42.115 51.555 ;
        RECT 42.445 51.325 44.405 51.555 ;
        RECT 44.735 51.325 46.695 51.555 ;
        RECT 47.025 51.325 48.985 51.555 ;
        RECT 50.655 51.325 52.615 51.555 ;
        RECT 52.945 51.325 54.905 51.555 ;
        RECT 55.235 51.325 57.195 51.555 ;
        RECT 57.525 51.325 59.485 51.555 ;
        RECT 59.815 51.325 61.775 51.555 ;
        RECT 62.105 51.325 64.065 51.555 ;
        RECT 64.395 51.325 66.355 51.555 ;
        RECT 66.685 51.325 68.645 51.555 ;
        RECT 70.315 51.325 72.275 51.555 ;
        RECT 72.605 51.325 74.565 51.555 ;
        RECT 74.895 51.325 76.855 51.555 ;
        RECT 77.185 51.325 79.145 51.555 ;
        RECT 79.475 51.325 81.435 51.555 ;
        RECT 81.765 51.325 83.725 51.555 ;
        RECT 84.055 51.325 86.015 51.555 ;
        RECT 86.345 51.325 88.305 51.555 ;
        RECT 89.975 51.325 91.935 51.555 ;
        RECT 92.265 51.325 94.225 51.555 ;
        RECT 94.555 51.325 96.515 51.555 ;
        RECT 96.845 51.325 98.805 51.555 ;
        RECT 99.135 51.325 101.095 51.555 ;
        RECT 101.425 51.325 103.385 51.555 ;
        RECT 103.715 51.325 105.675 51.555 ;
        RECT 106.005 51.325 107.965 51.555 ;
        RECT 109.355 51.325 127.905 52.935 ;
        RECT 11.055 42.915 11.285 51.325 ;
        RECT 13.345 42.915 13.575 51.325 ;
        RECT 15.635 42.915 15.865 51.325 ;
        RECT 17.925 42.915 18.155 51.325 ;
        RECT 20.215 42.915 20.445 51.325 ;
        RECT 22.505 42.915 22.735 51.325 ;
        RECT 24.795 42.915 25.025 51.325 ;
        RECT 27.085 42.915 27.315 51.325 ;
        RECT 29.375 42.915 29.605 51.325 ;
        RECT 11.055 42.225 29.605 42.915 ;
        RECT 30.715 42.915 30.945 51.120 ;
        RECT 33.005 42.915 33.235 51.120 ;
        RECT 35.295 42.915 35.525 51.120 ;
        RECT 37.585 42.915 37.815 51.120 ;
        RECT 39.875 42.915 40.105 51.120 ;
        RECT 42.165 42.915 42.395 51.120 ;
        RECT 44.455 42.915 44.685 51.120 ;
        RECT 46.745 42.915 46.975 51.120 ;
        RECT 49.035 42.915 49.265 51.120 ;
        RECT 30.715 42.225 49.265 42.915 ;
        RECT 50.375 42.915 50.605 51.120 ;
        RECT 52.665 42.915 52.895 51.120 ;
        RECT 54.955 42.915 55.185 51.120 ;
        RECT 57.245 42.915 57.475 51.120 ;
        RECT 59.535 42.915 59.765 51.120 ;
        RECT 61.825 42.915 62.055 51.120 ;
        RECT 64.115 42.915 64.345 51.120 ;
        RECT 66.405 42.915 66.635 51.120 ;
        RECT 68.695 42.915 68.925 51.120 ;
        RECT 50.375 42.225 68.925 42.915 ;
        RECT 70.035 42.915 70.265 51.120 ;
        RECT 72.325 42.915 72.555 51.120 ;
        RECT 74.615 42.915 74.845 51.120 ;
        RECT 76.905 42.915 77.135 51.120 ;
        RECT 79.195 42.915 79.425 51.120 ;
        RECT 81.485 42.915 81.715 51.120 ;
        RECT 83.775 42.915 84.005 51.120 ;
        RECT 86.065 42.915 86.295 51.120 ;
        RECT 88.355 42.915 88.585 51.120 ;
        RECT 70.035 42.225 88.585 42.915 ;
        RECT 89.695 42.915 89.925 51.120 ;
        RECT 91.985 42.915 92.215 51.120 ;
        RECT 94.275 42.915 94.505 51.120 ;
        RECT 96.565 42.915 96.795 51.120 ;
        RECT 98.855 42.915 99.085 51.120 ;
        RECT 101.145 42.915 101.375 51.120 ;
        RECT 103.435 42.915 103.665 51.120 ;
        RECT 105.725 42.915 105.955 51.120 ;
        RECT 108.015 42.915 108.245 51.120 ;
        RECT 89.695 42.225 108.245 42.915 ;
        RECT 109.355 42.915 109.585 51.325 ;
        RECT 111.645 42.915 111.875 51.325 ;
        RECT 113.935 42.915 114.165 51.325 ;
        RECT 116.225 42.915 116.455 51.325 ;
        RECT 118.515 42.915 118.745 51.325 ;
        RECT 120.805 42.915 121.035 51.325 ;
        RECT 123.095 42.915 123.325 51.325 ;
        RECT 125.385 42.915 125.615 51.325 ;
        RECT 127.675 42.915 127.905 51.325 ;
        RECT 109.355 42.225 127.905 42.915 ;
        RECT 128.345 42.225 135.710 102.115 ;
        RECT 136.295 100.155 138.400 101.915 ;
        RECT 136.295 97.815 138.400 99.575 ;
        RECT 136.295 95.475 138.400 97.235 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 141.695 93.725 142.995 108.925 ;
        RECT 149.570 107.765 155.900 137.690 ;
        RECT 246.345 108.365 246.665 108.425 ;
        RECT 280.845 108.365 281.165 108.425 ;
        RECT 297.865 108.365 298.185 108.425 ;
        RECT 246.345 108.225 298.185 108.365 ;
        RECT 246.345 108.165 246.665 108.225 ;
        RECT 280.845 108.165 281.165 108.225 ;
        RECT 297.865 108.165 298.185 108.225 ;
        RECT 146.290 104.835 155.900 107.765 ;
        RECT 224.265 107.685 224.585 107.745 ;
        RECT 267.965 107.685 268.285 107.745 ;
        RECT 288.205 107.685 288.525 107.745 ;
        RECT 300.165 107.685 300.485 107.745 ;
        RECT 224.265 107.545 283.605 107.685 ;
        RECT 224.265 107.485 224.585 107.545 ;
        RECT 267.965 107.485 268.285 107.545 ;
        RECT 218.745 107.345 219.065 107.405 ;
        RECT 252.785 107.345 253.105 107.405 ;
        RECT 218.745 107.205 253.105 107.345 ;
        RECT 218.745 107.145 219.065 107.205 ;
        RECT 252.785 107.145 253.105 107.205 ;
        RECT 265.205 107.345 265.525 107.405 ;
        RECT 276.245 107.345 276.565 107.405 ;
        RECT 265.205 107.205 276.565 107.345 ;
        RECT 283.465 107.345 283.605 107.545 ;
        RECT 288.205 107.545 300.485 107.685 ;
        RECT 288.205 107.485 288.525 107.545 ;
        RECT 300.165 107.485 300.485 107.545 ;
        RECT 290.045 107.345 290.365 107.405 ;
        RECT 283.465 107.205 290.365 107.345 ;
        RECT 265.205 107.145 265.525 107.205 ;
        RECT 276.245 107.145 276.565 107.205 ;
        RECT 290.045 107.145 290.365 107.205 ;
        RECT 221.045 107.005 221.365 107.065 ;
        RECT 223.805 107.005 224.125 107.065 ;
        RECT 221.045 106.865 224.125 107.005 ;
        RECT 221.045 106.805 221.365 106.865 ;
        RECT 223.805 106.805 224.125 106.865 ;
        RECT 241.745 107.005 242.065 107.065 ;
        RECT 267.045 107.005 267.365 107.065 ;
        RECT 241.745 106.865 267.365 107.005 ;
        RECT 241.745 106.805 242.065 106.865 ;
        RECT 267.045 106.805 267.365 106.865 ;
        RECT 274.405 107.005 274.725 107.065 ;
        RECT 283.145 107.005 283.465 107.065 ;
        RECT 274.405 106.865 283.465 107.005 ;
        RECT 274.405 106.805 274.725 106.865 ;
        RECT 283.145 106.805 283.465 106.865 ;
        RECT 292.805 107.005 293.125 107.065 ;
        RECT 302.465 107.005 302.785 107.065 ;
        RECT 292.805 106.865 302.785 107.005 ;
        RECT 292.805 106.805 293.125 106.865 ;
        RECT 302.465 106.805 302.785 106.865 ;
        RECT 162.095 106.185 311.935 106.665 ;
        RECT 164.005 105.985 164.325 106.045 ;
        RECT 164.480 105.985 164.770 106.030 ;
        RECT 164.005 105.845 164.770 105.985 ;
        RECT 164.005 105.785 164.325 105.845 ;
        RECT 164.480 105.800 164.770 105.845 ;
        RECT 166.305 105.985 166.625 106.045 ;
        RECT 168.160 105.985 168.450 106.030 ;
        RECT 166.305 105.845 168.450 105.985 ;
        RECT 166.305 105.785 166.625 105.845 ;
        RECT 168.160 105.800 168.450 105.845 ;
        RECT 170.905 105.785 171.225 106.045 ;
        RECT 172.760 105.985 173.050 106.030 ;
        RECT 173.205 105.985 173.525 106.045 ;
        RECT 172.760 105.845 173.525 105.985 ;
        RECT 172.760 105.800 173.050 105.845 ;
        RECT 173.205 105.785 173.525 105.845 ;
        RECT 176.900 105.985 177.190 106.030 ;
        RECT 177.805 105.985 178.125 106.045 ;
        RECT 176.900 105.845 178.125 105.985 ;
        RECT 176.900 105.800 177.190 105.845 ;
        RECT 177.805 105.785 178.125 105.845 ;
        RECT 180.105 105.785 180.425 106.045 ;
        RECT 183.340 105.985 183.630 106.030 ;
        RECT 184.705 105.985 185.025 106.045 ;
        RECT 183.340 105.845 185.025 105.985 ;
        RECT 183.340 105.800 183.630 105.845 ;
        RECT 184.705 105.785 185.025 105.845 ;
        RECT 187.005 105.985 187.325 106.045 ;
        RECT 188.860 105.985 189.150 106.030 ;
        RECT 187.005 105.845 189.150 105.985 ;
        RECT 187.005 105.785 187.325 105.845 ;
        RECT 188.860 105.800 189.150 105.845 ;
        RECT 193.000 105.985 193.290 106.030 ;
        RECT 193.905 105.985 194.225 106.045 ;
        RECT 193.000 105.845 194.225 105.985 ;
        RECT 193.000 105.800 193.290 105.845 ;
        RECT 193.905 105.785 194.225 105.845 ;
        RECT 196.205 105.785 196.525 106.045 ;
        RECT 197.600 105.985 197.890 106.030 ;
        RECT 198.045 105.985 198.365 106.045 ;
        RECT 197.600 105.845 198.365 105.985 ;
        RECT 197.600 105.800 197.890 105.845 ;
        RECT 198.045 105.785 198.365 105.845 ;
        RECT 200.805 105.985 201.125 106.045 ;
        RECT 201.740 105.985 202.030 106.030 ;
        RECT 200.805 105.845 202.030 105.985 ;
        RECT 200.805 105.785 201.125 105.845 ;
        RECT 201.740 105.800 202.030 105.845 ;
        RECT 205.880 105.985 206.170 106.030 ;
        RECT 207.705 105.985 208.025 106.045 ;
        RECT 205.880 105.845 208.025 105.985 ;
        RECT 205.880 105.800 206.170 105.845 ;
        RECT 207.705 105.785 208.025 105.845 ;
        RECT 209.100 105.985 209.390 106.030 ;
        RECT 211.385 105.985 211.705 106.045 ;
        RECT 209.100 105.845 211.705 105.985 ;
        RECT 209.100 105.800 209.390 105.845 ;
        RECT 211.385 105.785 211.705 105.845 ;
        RECT 212.305 105.785 212.625 106.045 ;
        RECT 214.605 105.785 214.925 106.045 ;
        RECT 218.745 105.785 219.065 106.045 ;
        RECT 219.220 105.985 219.510 106.030 ;
        RECT 221.045 105.985 221.365 106.045 ;
        RECT 219.220 105.845 221.365 105.985 ;
        RECT 219.220 105.800 219.510 105.845 ;
        RECT 221.045 105.785 221.365 105.845 ;
        RECT 221.505 105.985 221.825 106.045 ;
        RECT 221.980 105.985 222.270 106.030 ;
        RECT 221.505 105.845 222.270 105.985 ;
        RECT 221.505 105.785 221.825 105.845 ;
        RECT 221.980 105.800 222.270 105.845 ;
        RECT 223.820 105.985 224.110 106.030 ;
        RECT 226.105 105.985 226.425 106.045 ;
        RECT 223.820 105.845 226.425 105.985 ;
        RECT 223.820 105.800 224.110 105.845 ;
        RECT 226.105 105.785 226.425 105.845 ;
        RECT 227.960 105.985 228.250 106.030 ;
        RECT 228.405 105.985 228.725 106.045 ;
        RECT 227.960 105.845 228.725 105.985 ;
        RECT 227.960 105.800 228.250 105.845 ;
        RECT 228.405 105.785 228.725 105.845 ;
        RECT 231.180 105.985 231.470 106.030 ;
        RECT 233.005 105.985 233.325 106.045 ;
        RECT 231.180 105.845 233.325 105.985 ;
        RECT 231.180 105.800 231.470 105.845 ;
        RECT 233.005 105.785 233.325 105.845 ;
        RECT 235.305 105.985 235.625 106.045 ;
        RECT 235.780 105.985 236.070 106.030 ;
        RECT 235.305 105.845 236.070 105.985 ;
        RECT 235.305 105.785 235.625 105.845 ;
        RECT 235.780 105.800 236.070 105.845 ;
        RECT 238.540 105.985 238.830 106.030 ;
        RECT 239.905 105.985 240.225 106.045 ;
        RECT 238.540 105.845 240.225 105.985 ;
        RECT 238.540 105.800 238.830 105.845 ;
        RECT 239.905 105.785 240.225 105.845 ;
        RECT 242.205 105.985 242.525 106.045 ;
        RECT 248.660 105.985 248.950 106.030 ;
        RECT 242.205 105.845 248.950 105.985 ;
        RECT 242.205 105.785 242.525 105.845 ;
        RECT 248.660 105.800 248.950 105.845 ;
        RECT 253.705 105.985 254.025 106.045 ;
        RECT 256.020 105.985 256.310 106.030 ;
        RECT 253.705 105.845 256.310 105.985 ;
        RECT 253.705 105.785 254.025 105.845 ;
        RECT 256.020 105.800 256.310 105.845 ;
        RECT 260.605 105.985 260.925 106.045 ;
        RECT 261.540 105.985 261.830 106.030 ;
        RECT 260.605 105.845 261.830 105.985 ;
        RECT 260.605 105.785 260.925 105.845 ;
        RECT 261.540 105.800 261.830 105.845 ;
        RECT 262.905 105.785 263.225 106.045 ;
        RECT 267.505 105.985 267.825 106.045 ;
        RECT 268.900 105.985 269.190 106.030 ;
        RECT 267.505 105.845 269.190 105.985 ;
        RECT 267.505 105.785 267.825 105.845 ;
        RECT 268.900 105.800 269.190 105.845 ;
        RECT 269.805 105.985 270.125 106.045 ;
        RECT 271.660 105.985 271.950 106.030 ;
        RECT 269.805 105.845 271.950 105.985 ;
        RECT 269.805 105.785 270.125 105.845 ;
        RECT 271.660 105.800 271.950 105.845 ;
        RECT 274.420 105.800 274.710 106.030 ;
        RECT 169.540 105.645 169.830 105.690 ;
        RECT 181.945 105.645 182.265 105.705 ;
        RECT 169.540 105.505 182.265 105.645 ;
        RECT 169.540 105.460 169.830 105.505 ;
        RECT 181.945 105.445 182.265 105.505 ;
        RECT 194.380 105.645 194.670 105.690 ;
        RECT 196.665 105.645 196.985 105.705 ;
        RECT 194.380 105.505 196.985 105.645 ;
        RECT 194.380 105.460 194.670 105.505 ;
        RECT 196.665 105.445 196.985 105.505 ;
        RECT 197.125 105.645 197.445 105.705 ;
        RECT 199.885 105.645 200.205 105.705 ;
        RECT 218.835 105.645 218.975 105.785 ;
        RECT 244.505 105.645 244.825 105.705 ;
        RECT 252.800 105.645 253.090 105.690 ;
        RECT 197.125 105.505 199.195 105.645 ;
        RECT 197.125 105.445 197.445 105.505 ;
        RECT 165.400 105.305 165.690 105.350 ;
        RECT 171.840 105.305 172.130 105.350 ;
        RECT 165.400 105.165 167.455 105.305 ;
        RECT 165.400 105.120 165.690 105.165 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 146.290 101.325 148.395 103.085 ;
        RECT 146.290 98.985 148.395 100.745 ;
        RECT 146.290 96.645 148.395 98.405 ;
        RECT 146.290 94.305 148.395 96.065 ;
        RECT 136.295 91.965 138.400 93.725 ;
        RECT 141.695 93.135 148.395 93.725 ;
        RECT 146.290 91.965 148.395 92.555 ;
        RECT 136.295 90.795 143.395 91.385 ;
        RECT 136.295 89.625 138.400 90.215 ;
        RECT 146.290 89.625 148.395 91.385 ;
        RECT 136.295 87.285 138.400 89.045 ;
        RECT 146.290 88.455 148.395 89.045 ;
        RECT 146.290 87.285 148.395 87.875 ;
        RECT 136.295 86.115 138.400 86.705 ;
        RECT 136.295 84.945 138.400 85.535 ;
        RECT 146.290 84.945 148.395 86.705 ;
        RECT 136.295 82.605 138.400 84.365 ;
        RECT 146.290 83.775 148.395 84.365 ;
        RECT 146.290 82.605 148.395 83.195 ;
        RECT 136.295 81.435 141.260 82.025 ;
        RECT 143.790 81.435 148.395 82.025 ;
        RECT 136.295 80.265 138.400 80.855 ;
        RECT 136.295 79.095 138.400 79.685 ;
        RECT 136.295 76.755 138.400 78.515 ;
        RECT 136.295 75.585 138.400 76.175 ;
        RECT 136.295 74.415 138.400 75.005 ;
        RECT 136.295 72.075 138.400 73.835 ;
        RECT 136.295 70.905 138.400 71.495 ;
        RECT 136.295 69.735 138.400 70.325 ;
        RECT 136.295 67.395 138.400 69.155 ;
        RECT 136.295 66.225 138.400 66.815 ;
        RECT 136.295 65.055 138.400 65.645 ;
        RECT 136.295 62.715 138.400 64.475 ;
        RECT 143.790 62.135 145.190 81.435 ;
        RECT 146.290 79.095 148.395 80.855 ;
        RECT 146.290 77.925 148.395 78.515 ;
        RECT 146.290 76.755 148.395 77.345 ;
        RECT 146.290 74.415 148.395 76.175 ;
        RECT 146.290 73.245 148.395 73.835 ;
        RECT 146.290 72.075 148.395 72.665 ;
        RECT 146.290 69.735 148.395 71.495 ;
        RECT 146.290 68.565 148.395 69.155 ;
        RECT 146.290 67.395 148.395 67.985 ;
        RECT 146.290 65.055 148.395 66.815 ;
        RECT 146.290 63.885 148.395 64.475 ;
        RECT 146.290 62.715 148.395 63.305 ;
        RECT 136.295 61.545 140.910 62.135 ;
        RECT 143.790 61.545 148.395 62.135 ;
        RECT 136.295 60.375 138.400 60.965 ;
        RECT 136.295 59.205 138.400 59.795 ;
        RECT 136.295 56.865 138.400 58.625 ;
        RECT 136.295 55.695 138.400 56.285 ;
        RECT 136.295 54.525 138.400 55.115 ;
        RECT 136.295 52.185 138.400 53.945 ;
        RECT 136.295 51.015 138.400 51.605 ;
        RECT 136.295 49.845 138.400 50.435 ;
        RECT 136.295 47.505 138.400 49.265 ;
        RECT 136.295 46.335 138.400 46.925 ;
        RECT 136.295 45.165 138.400 45.755 ;
        RECT 136.295 42.825 138.400 44.585 ;
        RECT 139.510 42.245 140.910 61.545 ;
        RECT 146.290 59.205 148.395 60.965 ;
        RECT 146.290 58.035 148.395 58.625 ;
        RECT 146.290 56.865 148.395 57.455 ;
        RECT 146.290 54.525 148.395 56.285 ;
        RECT 146.290 53.355 148.395 53.945 ;
        RECT 146.290 52.185 148.395 52.775 ;
        RECT 146.290 49.845 148.395 51.605 ;
        RECT 146.290 48.675 148.395 49.265 ;
        RECT 146.290 47.505 148.395 48.095 ;
        RECT 146.290 45.165 148.395 46.925 ;
        RECT 146.290 43.995 148.395 44.585 ;
        RECT 146.290 42.825 148.395 43.415 ;
        RECT 4.100 41.635 135.710 42.225 ;
        RECT 136.295 41.655 140.910 42.245 ;
        RECT 143.435 41.655 148.395 42.245 ;
        RECT 4.100 4.900 4.900 41.635 ;
        RECT 7.065 39.040 130.565 39.630 ;
        RECT 7.065 36.430 10.615 39.040 ;
        RECT 8.665 9.480 10.615 36.430 ;
        RECT 11.115 38.350 20.505 38.580 ;
        RECT 22.015 38.350 30.845 38.650 ;
        RECT 32.635 38.350 41.465 38.650 ;
        RECT 43.255 38.350 52.085 38.650 ;
        RECT 53.875 38.350 62.705 38.650 ;
        RECT 64.215 38.350 73.605 38.580 ;
        RECT 11.115 34.890 11.345 38.350 ;
        RECT 13.405 34.890 13.635 38.190 ;
        RECT 15.695 34.890 15.925 38.350 ;
        RECT 17.985 34.890 18.215 38.190 ;
        RECT 20.275 34.890 20.505 38.350 ;
        RECT 11.020 33.490 11.345 34.890 ;
        RECT 13.370 33.490 13.670 34.890 ;
        RECT 15.660 33.490 15.960 34.890 ;
        RECT 17.950 33.490 18.250 34.890 ;
        RECT 20.240 33.490 20.540 34.890 ;
        RECT 11.115 30.030 11.345 33.490 ;
        RECT 13.405 30.190 13.635 33.490 ;
        RECT 15.695 30.030 15.925 33.490 ;
        RECT 17.985 30.190 18.215 33.490 ;
        RECT 20.275 30.030 20.505 33.490 ;
        RECT 21.735 32.890 21.965 38.190 ;
        RECT 24.025 34.890 24.255 38.190 ;
        RECT 26.315 36.890 26.545 38.190 ;
        RECT 26.280 35.490 26.580 36.890 ;
        RECT 23.990 33.490 24.290 34.890 ;
        RECT 21.700 31.490 22.000 32.890 ;
        RECT 21.735 30.190 21.965 31.490 ;
        RECT 24.025 30.190 24.255 33.490 ;
        RECT 26.315 30.190 26.545 35.490 ;
        RECT 28.605 34.890 28.835 38.190 ;
        RECT 28.570 33.490 28.870 34.890 ;
        RECT 28.605 30.190 28.835 33.490 ;
        RECT 30.895 32.890 31.125 38.190 ;
        RECT 32.355 36.890 32.585 38.190 ;
        RECT 32.320 35.490 32.620 36.890 ;
        RECT 30.860 31.490 31.160 32.890 ;
        RECT 30.895 30.190 31.125 31.490 ;
        RECT 32.355 30.190 32.585 35.490 ;
        RECT 34.645 34.890 34.875 38.190 ;
        RECT 34.610 33.490 34.910 34.890 ;
        RECT 34.645 30.190 34.875 33.490 ;
        RECT 36.935 32.890 37.165 38.190 ;
        RECT 39.225 34.890 39.455 38.190 ;
        RECT 41.515 36.890 41.745 38.190 ;
        RECT 41.480 35.490 41.780 36.890 ;
        RECT 39.190 33.490 39.490 34.890 ;
        RECT 36.900 31.490 37.200 32.890 ;
        RECT 36.935 30.190 37.165 31.490 ;
        RECT 39.225 30.190 39.455 33.490 ;
        RECT 41.515 30.190 41.745 35.490 ;
        RECT 42.975 32.890 43.205 38.190 ;
        RECT 45.265 34.890 45.495 38.190 ;
        RECT 47.555 36.890 47.785 38.190 ;
        RECT 47.520 35.490 47.820 36.890 ;
        RECT 45.230 33.490 45.530 34.890 ;
        RECT 42.940 31.490 43.240 32.890 ;
        RECT 42.975 30.190 43.205 31.490 ;
        RECT 45.265 30.190 45.495 33.490 ;
        RECT 47.555 30.190 47.785 35.490 ;
        RECT 49.845 34.890 50.075 38.190 ;
        RECT 49.810 33.490 50.110 34.890 ;
        RECT 49.845 30.190 50.075 33.490 ;
        RECT 52.135 32.890 52.365 38.190 ;
        RECT 53.595 36.890 53.825 38.190 ;
        RECT 53.560 35.490 53.860 36.890 ;
        RECT 52.100 31.490 52.400 32.890 ;
        RECT 52.135 30.190 52.365 31.490 ;
        RECT 53.595 30.190 53.825 35.490 ;
        RECT 55.885 34.890 56.115 38.190 ;
        RECT 55.850 33.490 56.150 34.890 ;
        RECT 55.885 30.190 56.115 33.490 ;
        RECT 58.175 32.890 58.405 38.190 ;
        RECT 60.465 34.890 60.695 38.190 ;
        RECT 62.755 36.890 62.985 38.190 ;
        RECT 62.720 35.490 63.020 36.890 ;
        RECT 60.430 33.490 60.730 34.890 ;
        RECT 58.140 31.490 58.440 32.890 ;
        RECT 58.175 30.190 58.405 31.490 ;
        RECT 60.465 30.190 60.695 33.490 ;
        RECT 62.755 30.190 62.985 35.490 ;
        RECT 64.215 34.890 64.445 38.350 ;
        RECT 66.505 34.890 66.735 38.190 ;
        RECT 68.795 34.890 69.025 38.350 ;
        RECT 71.085 34.890 71.315 38.190 ;
        RECT 73.375 34.890 73.605 38.350 ;
        RECT 64.180 33.490 64.480 34.890 ;
        RECT 66.470 33.490 66.770 34.890 ;
        RECT 68.760 33.490 69.060 34.890 ;
        RECT 71.050 33.490 71.350 34.890 ;
        RECT 73.340 33.490 73.640 34.890 ;
        RECT 64.215 30.030 64.445 33.490 ;
        RECT 66.505 30.190 66.735 33.490 ;
        RECT 68.795 30.030 69.025 33.490 ;
        RECT 71.085 30.190 71.315 33.490 ;
        RECT 73.375 30.030 73.605 33.490 ;
        RECT 11.115 29.800 20.505 30.030 ;
        RECT 22.015 29.730 30.845 30.030 ;
        RECT 32.635 29.730 41.465 30.030 ;
        RECT 43.255 29.730 52.085 30.030 ;
        RECT 53.875 29.730 62.705 30.030 ;
        RECT 64.215 29.800 73.605 30.030 ;
        RECT 11.115 28.420 20.505 28.650 ;
        RECT 22.015 28.420 30.845 28.720 ;
        RECT 32.635 28.650 41.465 28.720 ;
        RECT 43.255 28.650 52.085 28.720 ;
        RECT 32.355 28.420 41.745 28.650 ;
        RECT 11.115 24.960 11.345 28.420 ;
        RECT 13.405 24.960 13.635 28.260 ;
        RECT 15.695 24.960 15.925 28.420 ;
        RECT 17.985 24.960 18.215 28.260 ;
        RECT 20.275 24.960 20.505 28.420 ;
        RECT 21.735 26.960 21.965 28.260 ;
        RECT 21.700 25.560 22.000 26.960 ;
        RECT 11.020 23.560 11.345 24.960 ;
        RECT 13.370 23.560 13.670 24.960 ;
        RECT 15.660 23.560 15.960 24.960 ;
        RECT 17.950 23.560 18.250 24.960 ;
        RECT 20.240 23.560 20.540 24.960 ;
        RECT 11.115 20.100 11.345 23.560 ;
        RECT 13.405 20.260 13.635 23.560 ;
        RECT 15.695 20.100 15.925 23.560 ;
        RECT 17.985 20.260 18.215 23.560 ;
        RECT 20.275 20.100 20.505 23.560 ;
        RECT 21.735 20.260 21.965 25.560 ;
        RECT 24.025 24.960 24.255 28.260 ;
        RECT 23.990 23.560 24.290 24.960 ;
        RECT 24.025 20.260 24.255 23.560 ;
        RECT 26.315 22.960 26.545 28.260 ;
        RECT 28.605 24.960 28.835 28.260 ;
        RECT 30.895 26.960 31.125 28.260 ;
        RECT 30.860 25.560 31.160 26.960 ;
        RECT 28.570 23.560 28.870 24.960 ;
        RECT 26.280 21.560 26.580 22.960 ;
        RECT 26.315 20.260 26.545 21.560 ;
        RECT 28.605 20.260 28.835 23.560 ;
        RECT 30.895 20.260 31.125 25.560 ;
        RECT 32.355 20.100 32.585 28.420 ;
        RECT 34.645 24.960 34.875 28.260 ;
        RECT 34.610 23.560 34.910 24.960 ;
        RECT 34.645 20.260 34.875 23.560 ;
        RECT 36.935 20.100 37.165 28.420 ;
        RECT 39.225 24.960 39.455 28.260 ;
        RECT 39.190 23.560 39.490 24.960 ;
        RECT 39.225 20.260 39.455 23.560 ;
        RECT 41.515 20.100 41.745 28.420 ;
        RECT 11.115 19.870 20.505 20.100 ;
        RECT 22.015 19.800 30.845 20.100 ;
        RECT 32.355 19.870 41.745 20.100 ;
        RECT 42.975 28.420 52.365 28.650 ;
        RECT 53.875 28.420 62.705 28.720 ;
        RECT 64.215 28.420 73.605 28.650 ;
        RECT 42.975 20.100 43.205 28.420 ;
        RECT 45.265 24.960 45.495 28.260 ;
        RECT 45.230 23.560 45.530 24.960 ;
        RECT 45.265 20.260 45.495 23.560 ;
        RECT 47.555 20.100 47.785 28.420 ;
        RECT 49.845 24.960 50.075 28.260 ;
        RECT 49.810 23.560 50.110 24.960 ;
        RECT 49.845 20.260 50.075 23.560 ;
        RECT 52.135 20.100 52.365 28.420 ;
        RECT 53.595 22.960 53.825 28.260 ;
        RECT 55.885 24.960 56.115 28.260 ;
        RECT 58.175 26.960 58.405 28.260 ;
        RECT 58.140 25.560 58.440 26.960 ;
        RECT 55.850 23.560 56.150 24.960 ;
        RECT 53.560 21.560 53.860 22.960 ;
        RECT 53.595 20.260 53.825 21.560 ;
        RECT 55.885 20.260 56.115 23.560 ;
        RECT 58.175 20.260 58.405 25.560 ;
        RECT 60.465 24.960 60.695 28.260 ;
        RECT 60.430 23.560 60.730 24.960 ;
        RECT 60.465 20.260 60.695 23.560 ;
        RECT 62.755 22.960 62.985 28.260 ;
        RECT 64.215 24.960 64.445 28.420 ;
        RECT 66.505 24.960 66.735 28.260 ;
        RECT 68.795 24.960 69.025 28.420 ;
        RECT 71.085 24.960 71.315 28.260 ;
        RECT 73.375 24.960 73.605 28.420 ;
        RECT 64.180 23.560 64.480 24.960 ;
        RECT 66.470 23.560 66.770 24.960 ;
        RECT 68.760 23.560 69.060 24.960 ;
        RECT 71.050 23.560 71.350 24.960 ;
        RECT 73.340 23.560 73.640 24.960 ;
        RECT 62.720 21.560 63.020 22.960 ;
        RECT 62.755 20.260 62.985 21.560 ;
        RECT 64.215 20.100 64.445 23.560 ;
        RECT 66.505 20.260 66.735 23.560 ;
        RECT 68.795 20.100 69.025 23.560 ;
        RECT 71.085 20.260 71.315 23.560 ;
        RECT 73.375 20.100 73.605 23.560 ;
        RECT 42.975 19.870 52.365 20.100 ;
        RECT 32.635 19.800 41.465 19.870 ;
        RECT 43.255 19.800 52.085 19.870 ;
        RECT 53.875 19.800 62.705 20.100 ;
        RECT 64.215 19.870 73.605 20.100 ;
        RECT 11.115 18.490 20.505 18.720 ;
        RECT 22.015 18.490 30.845 18.790 ;
        RECT 32.635 18.490 41.465 18.790 ;
        RECT 43.255 18.490 52.085 18.790 ;
        RECT 53.875 18.490 62.705 18.790 ;
        RECT 64.215 18.490 73.605 18.720 ;
        RECT 11.115 15.030 11.345 18.490 ;
        RECT 13.405 15.030 13.635 18.330 ;
        RECT 15.695 15.030 15.925 18.490 ;
        RECT 17.985 15.030 18.215 18.330 ;
        RECT 20.275 15.030 20.505 18.490 ;
        RECT 11.020 13.630 11.345 15.030 ;
        RECT 13.370 13.630 13.670 15.030 ;
        RECT 15.660 13.630 15.960 15.030 ;
        RECT 17.950 13.630 18.250 15.030 ;
        RECT 20.240 13.630 20.540 15.030 ;
        RECT 11.115 10.170 11.345 13.630 ;
        RECT 13.405 10.330 13.635 13.630 ;
        RECT 15.695 10.170 15.925 13.630 ;
        RECT 17.985 10.330 18.215 13.630 ;
        RECT 20.275 10.170 20.505 13.630 ;
        RECT 21.735 13.030 21.965 18.330 ;
        RECT 24.025 15.030 24.255 18.330 ;
        RECT 26.315 17.030 26.545 18.330 ;
        RECT 26.280 15.630 26.580 17.030 ;
        RECT 23.990 13.630 24.290 15.030 ;
        RECT 21.700 11.630 22.000 13.030 ;
        RECT 21.735 10.330 21.965 11.630 ;
        RECT 24.025 10.330 24.255 13.630 ;
        RECT 26.315 10.330 26.545 15.630 ;
        RECT 28.605 15.030 28.835 18.330 ;
        RECT 28.570 13.630 28.870 15.030 ;
        RECT 28.605 10.330 28.835 13.630 ;
        RECT 30.895 13.030 31.125 18.330 ;
        RECT 32.355 17.030 32.585 18.330 ;
        RECT 32.320 15.630 32.620 17.030 ;
        RECT 30.860 11.630 31.160 13.030 ;
        RECT 30.895 10.330 31.125 11.630 ;
        RECT 32.355 10.330 32.585 15.630 ;
        RECT 34.645 15.030 34.875 18.330 ;
        RECT 34.610 13.630 34.910 15.030 ;
        RECT 34.645 10.330 34.875 13.630 ;
        RECT 36.935 13.030 37.165 18.330 ;
        RECT 39.225 15.030 39.455 18.330 ;
        RECT 41.515 17.030 41.745 18.330 ;
        RECT 41.480 15.630 41.780 17.030 ;
        RECT 39.190 13.630 39.490 15.030 ;
        RECT 36.900 11.630 37.200 13.030 ;
        RECT 36.935 10.330 37.165 11.630 ;
        RECT 39.225 10.330 39.455 13.630 ;
        RECT 41.515 10.330 41.745 15.630 ;
        RECT 42.975 13.030 43.205 18.330 ;
        RECT 45.265 15.030 45.495 18.330 ;
        RECT 47.555 17.030 47.785 18.330 ;
        RECT 47.520 15.630 47.820 17.030 ;
        RECT 45.230 13.630 45.530 15.030 ;
        RECT 42.940 11.630 43.240 13.030 ;
        RECT 42.975 10.330 43.205 11.630 ;
        RECT 45.265 10.330 45.495 13.630 ;
        RECT 47.555 10.330 47.785 15.630 ;
        RECT 49.845 15.030 50.075 18.330 ;
        RECT 49.810 13.630 50.110 15.030 ;
        RECT 49.845 10.330 50.075 13.630 ;
        RECT 52.135 13.030 52.365 18.330 ;
        RECT 53.595 17.030 53.825 18.330 ;
        RECT 53.560 15.630 53.860 17.030 ;
        RECT 52.100 11.630 52.400 13.030 ;
        RECT 52.135 10.330 52.365 11.630 ;
        RECT 53.595 10.330 53.825 15.630 ;
        RECT 55.885 15.030 56.115 18.330 ;
        RECT 55.850 13.630 56.150 15.030 ;
        RECT 55.885 10.330 56.115 13.630 ;
        RECT 58.175 13.030 58.405 18.330 ;
        RECT 60.465 15.030 60.695 18.330 ;
        RECT 62.755 17.030 62.985 18.330 ;
        RECT 62.720 15.630 63.020 17.030 ;
        RECT 60.430 13.630 60.730 15.030 ;
        RECT 58.140 11.630 58.440 13.030 ;
        RECT 58.175 10.330 58.405 11.630 ;
        RECT 60.465 10.330 60.695 13.630 ;
        RECT 62.755 10.330 62.985 15.630 ;
        RECT 64.215 15.030 64.445 18.490 ;
        RECT 66.505 15.030 66.735 18.330 ;
        RECT 68.795 15.030 69.025 18.490 ;
        RECT 71.085 15.030 71.315 18.330 ;
        RECT 73.375 15.030 73.605 18.490 ;
        RECT 64.180 13.630 64.480 15.030 ;
        RECT 66.470 13.630 66.770 15.030 ;
        RECT 68.760 13.630 69.060 15.030 ;
        RECT 71.050 13.630 71.350 15.030 ;
        RECT 73.340 13.630 73.640 15.030 ;
        RECT 64.215 10.170 64.445 13.630 ;
        RECT 66.505 10.330 66.735 13.630 ;
        RECT 68.795 10.170 69.025 13.630 ;
        RECT 71.085 10.330 71.315 13.630 ;
        RECT 73.375 10.170 73.605 13.630 ;
        RECT 11.115 9.940 20.505 10.170 ;
        RECT 22.015 9.870 30.845 10.170 ;
        RECT 32.635 9.870 41.465 10.170 ;
        RECT 43.255 9.870 52.085 10.170 ;
        RECT 53.875 9.870 62.705 10.170 ;
        RECT 64.215 9.940 73.605 10.170 ;
        RECT 74.105 9.480 80.255 39.040 ;
        RECT 81.035 38.350 82.995 38.580 ;
        RECT 83.325 38.350 85.285 38.580 ;
        RECT 87.075 38.350 89.035 38.700 ;
        RECT 89.365 38.350 91.325 38.700 ;
        RECT 93.115 38.350 97.365 38.700 ;
        RECT 99.155 38.350 101.115 38.700 ;
        RECT 101.445 38.350 103.405 38.700 ;
        RECT 105.195 38.350 107.155 38.700 ;
        RECT 107.485 38.350 109.445 38.700 ;
        RECT 111.235 38.350 115.485 38.700 ;
        RECT 117.275 38.350 119.235 38.700 ;
        RECT 119.565 38.350 121.525 38.700 ;
        RECT 123.315 38.350 125.275 38.580 ;
        RECT 125.605 38.350 127.565 38.580 ;
        RECT 80.755 30.190 80.985 38.190 ;
        RECT 83.045 30.190 83.275 38.190 ;
        RECT 85.335 30.190 85.565 38.190 ;
        RECT 86.795 35.995 87.025 38.190 ;
        RECT 86.560 35.295 87.260 35.995 ;
        RECT 86.795 30.190 87.025 35.295 ;
        RECT 89.085 34.495 89.315 38.190 ;
        RECT 91.375 35.995 91.605 38.190 ;
        RECT 92.835 37.495 93.065 38.190 ;
        RECT 92.600 36.795 93.300 37.495 ;
        RECT 91.140 35.295 91.840 35.995 ;
        RECT 88.850 33.795 89.550 34.495 ;
        RECT 89.085 30.190 89.315 33.795 ;
        RECT 91.375 30.190 91.605 35.295 ;
        RECT 92.835 30.190 93.065 36.795 ;
        RECT 95.125 30.190 95.355 38.350 ;
        RECT 97.415 37.495 97.645 38.190 ;
        RECT 97.180 36.795 97.880 37.495 ;
        RECT 97.415 30.190 97.645 36.795 ;
        RECT 98.875 31.495 99.105 38.190 ;
        RECT 101.165 32.995 101.395 38.190 ;
        RECT 100.930 32.295 101.630 32.995 ;
        RECT 98.640 30.795 99.340 31.495 ;
        RECT 98.875 30.190 99.105 30.795 ;
        RECT 101.165 30.190 101.395 32.295 ;
        RECT 103.455 31.495 103.685 38.190 ;
        RECT 104.915 31.495 105.145 38.190 ;
        RECT 107.205 32.995 107.435 38.190 ;
        RECT 106.970 32.295 107.670 32.995 ;
        RECT 103.220 30.795 103.920 31.495 ;
        RECT 104.680 30.795 105.380 31.495 ;
        RECT 103.455 30.190 103.685 30.795 ;
        RECT 104.915 30.190 105.145 30.795 ;
        RECT 107.205 30.190 107.435 32.295 ;
        RECT 109.495 31.495 109.725 38.190 ;
        RECT 110.955 37.495 111.185 38.190 ;
        RECT 110.720 36.795 111.420 37.495 ;
        RECT 109.260 30.795 109.960 31.495 ;
        RECT 109.495 30.190 109.725 30.795 ;
        RECT 110.955 30.190 111.185 36.795 ;
        RECT 113.245 30.190 113.475 38.350 ;
        RECT 115.535 37.495 115.765 38.190 ;
        RECT 115.300 36.795 116.000 37.495 ;
        RECT 115.535 30.190 115.765 36.795 ;
        RECT 116.995 35.995 117.225 38.190 ;
        RECT 116.760 35.295 117.460 35.995 ;
        RECT 116.995 30.190 117.225 35.295 ;
        RECT 119.285 34.495 119.515 38.190 ;
        RECT 121.575 35.995 121.805 38.190 ;
        RECT 121.340 35.295 122.040 35.995 ;
        RECT 119.050 33.795 119.750 34.495 ;
        RECT 119.285 30.190 119.515 33.795 ;
        RECT 121.575 30.190 121.805 35.295 ;
        RECT 123.035 30.190 123.265 38.190 ;
        RECT 125.325 30.190 125.555 38.190 ;
        RECT 127.615 30.190 127.845 38.190 ;
        RECT 81.035 29.800 82.995 30.030 ;
        RECT 83.325 29.800 85.285 30.030 ;
        RECT 87.075 29.680 89.035 30.030 ;
        RECT 89.365 29.680 91.325 30.030 ;
        RECT 93.115 29.680 95.075 30.030 ;
        RECT 95.405 29.680 97.365 30.030 ;
        RECT 99.155 29.680 101.115 30.030 ;
        RECT 101.445 29.680 103.405 30.030 ;
        RECT 105.195 29.680 107.155 30.030 ;
        RECT 107.485 29.680 109.445 30.030 ;
        RECT 111.235 29.680 113.195 30.030 ;
        RECT 113.525 29.680 115.485 30.030 ;
        RECT 117.275 29.680 119.235 30.030 ;
        RECT 119.565 29.680 121.525 30.030 ;
        RECT 123.315 29.800 125.275 30.030 ;
        RECT 125.605 29.800 127.565 30.030 ;
        RECT 81.035 28.420 82.995 28.650 ;
        RECT 83.325 28.420 85.285 28.650 ;
        RECT 87.075 28.420 89.035 28.770 ;
        RECT 89.365 28.420 91.325 28.770 ;
        RECT 93.115 28.420 95.075 28.770 ;
        RECT 95.405 28.420 97.365 28.770 ;
        RECT 99.155 28.420 101.115 28.770 ;
        RECT 101.445 28.420 103.405 28.770 ;
        RECT 105.195 28.420 107.155 28.770 ;
        RECT 107.485 28.420 109.445 28.770 ;
        RECT 111.235 28.420 113.195 28.770 ;
        RECT 113.525 28.420 115.485 28.770 ;
        RECT 117.275 28.420 119.235 28.770 ;
        RECT 119.565 28.420 121.525 28.770 ;
        RECT 123.315 28.420 125.275 28.650 ;
        RECT 125.605 28.420 127.565 28.650 ;
        RECT 80.755 20.260 80.985 28.260 ;
        RECT 83.045 20.260 83.275 28.260 ;
        RECT 85.335 20.260 85.565 28.260 ;
        RECT 86.795 23.065 87.025 28.260 ;
        RECT 89.085 24.565 89.315 28.260 ;
        RECT 88.850 23.865 89.550 24.565 ;
        RECT 86.560 22.365 87.260 23.065 ;
        RECT 86.795 20.260 87.025 22.365 ;
        RECT 89.085 20.260 89.315 23.865 ;
        RECT 91.375 23.065 91.605 28.260 ;
        RECT 91.140 22.365 91.840 23.065 ;
        RECT 91.375 20.260 91.605 22.365 ;
        RECT 92.835 21.565 93.065 28.260 ;
        RECT 92.600 20.865 93.300 21.565 ;
        RECT 92.835 20.260 93.065 20.865 ;
        RECT 95.125 20.100 95.355 28.260 ;
        RECT 97.415 21.565 97.645 28.260 ;
        RECT 98.875 27.565 99.105 28.260 ;
        RECT 98.640 26.865 99.340 27.565 ;
        RECT 97.180 20.865 97.880 21.565 ;
        RECT 97.415 20.260 97.645 20.865 ;
        RECT 98.875 20.260 99.105 26.865 ;
        RECT 101.165 26.065 101.395 28.260 ;
        RECT 103.455 27.565 103.685 28.260 ;
        RECT 104.915 27.565 105.145 28.260 ;
        RECT 103.220 26.865 103.920 27.565 ;
        RECT 104.680 26.865 105.380 27.565 ;
        RECT 100.930 25.365 101.630 26.065 ;
        RECT 101.165 20.260 101.395 25.365 ;
        RECT 103.455 20.260 103.685 26.865 ;
        RECT 104.915 20.260 105.145 26.865 ;
        RECT 107.205 26.065 107.435 28.260 ;
        RECT 109.495 27.565 109.725 28.260 ;
        RECT 109.260 26.865 109.960 27.565 ;
        RECT 106.970 25.365 107.670 26.065 ;
        RECT 107.205 20.260 107.435 25.365 ;
        RECT 109.495 20.260 109.725 26.865 ;
        RECT 110.955 21.565 111.185 28.260 ;
        RECT 110.720 20.865 111.420 21.565 ;
        RECT 110.955 20.260 111.185 20.865 ;
        RECT 113.245 20.100 113.475 28.260 ;
        RECT 115.535 21.565 115.765 28.260 ;
        RECT 116.995 23.065 117.225 28.260 ;
        RECT 119.285 24.565 119.515 28.260 ;
        RECT 119.050 23.865 119.750 24.565 ;
        RECT 116.760 22.365 117.460 23.065 ;
        RECT 115.300 20.865 116.000 21.565 ;
        RECT 115.535 20.260 115.765 20.865 ;
        RECT 116.995 20.260 117.225 22.365 ;
        RECT 119.285 20.260 119.515 23.865 ;
        RECT 121.575 23.065 121.805 28.260 ;
        RECT 121.340 22.365 122.040 23.065 ;
        RECT 121.575 20.260 121.805 22.365 ;
        RECT 123.035 20.260 123.265 28.260 ;
        RECT 125.325 20.260 125.555 28.260 ;
        RECT 127.615 20.260 127.845 28.260 ;
        RECT 81.035 19.870 82.995 20.100 ;
        RECT 83.325 19.870 85.285 20.100 ;
        RECT 87.075 19.750 89.035 20.100 ;
        RECT 89.365 19.750 91.325 20.100 ;
        RECT 93.115 19.750 97.365 20.100 ;
        RECT 99.155 19.750 101.115 20.100 ;
        RECT 101.445 19.750 103.405 20.100 ;
        RECT 105.195 19.750 107.155 20.100 ;
        RECT 107.485 19.750 109.445 20.100 ;
        RECT 111.235 19.750 115.485 20.100 ;
        RECT 117.275 19.750 119.235 20.100 ;
        RECT 119.565 19.750 121.525 20.100 ;
        RECT 123.315 19.870 125.275 20.100 ;
        RECT 125.605 19.870 127.565 20.100 ;
        RECT 81.035 18.490 82.995 18.720 ;
        RECT 83.325 18.490 85.285 18.720 ;
        RECT 87.075 18.490 89.035 18.720 ;
        RECT 89.365 18.490 91.325 18.720 ;
        RECT 93.115 18.490 95.075 18.720 ;
        RECT 95.405 18.490 97.365 18.720 ;
        RECT 99.155 18.490 101.115 18.720 ;
        RECT 101.445 18.490 103.405 18.720 ;
        RECT 105.195 18.490 107.155 18.720 ;
        RECT 107.485 18.490 109.445 18.720 ;
        RECT 111.235 18.490 113.195 18.720 ;
        RECT 113.525 18.490 115.485 18.720 ;
        RECT 117.275 18.490 119.235 18.720 ;
        RECT 119.565 18.490 121.525 18.720 ;
        RECT 123.315 18.490 125.275 18.720 ;
        RECT 125.605 18.490 127.565 18.720 ;
        RECT 80.755 10.330 80.985 18.330 ;
        RECT 83.045 10.330 83.275 18.330 ;
        RECT 85.335 10.330 85.565 18.330 ;
        RECT 86.795 10.330 87.025 18.330 ;
        RECT 89.085 10.330 89.315 18.330 ;
        RECT 91.375 10.330 91.605 18.330 ;
        RECT 92.835 10.330 93.065 18.330 ;
        RECT 95.125 10.330 95.355 18.330 ;
        RECT 97.415 10.330 97.645 18.330 ;
        RECT 98.875 10.330 99.105 18.330 ;
        RECT 101.165 10.330 101.395 18.330 ;
        RECT 103.455 10.330 103.685 18.330 ;
        RECT 104.915 10.330 105.145 18.330 ;
        RECT 107.205 10.330 107.435 18.330 ;
        RECT 109.495 10.330 109.725 18.330 ;
        RECT 110.955 10.330 111.185 18.330 ;
        RECT 113.245 10.330 113.475 18.330 ;
        RECT 115.535 10.330 115.765 18.330 ;
        RECT 116.995 10.330 117.225 18.330 ;
        RECT 119.285 10.330 119.515 18.330 ;
        RECT 121.575 10.330 121.805 18.330 ;
        RECT 123.035 10.330 123.265 18.330 ;
        RECT 125.325 10.330 125.555 18.330 ;
        RECT 127.615 10.330 127.845 18.330 ;
        RECT 81.035 9.940 82.995 10.170 ;
        RECT 83.325 9.940 85.285 10.170 ;
        RECT 87.075 9.940 89.035 10.170 ;
        RECT 89.365 9.940 91.325 10.170 ;
        RECT 93.115 9.940 95.075 10.170 ;
        RECT 95.405 9.940 97.365 10.170 ;
        RECT 99.155 9.940 101.115 10.170 ;
        RECT 101.445 9.940 103.405 10.170 ;
        RECT 105.195 9.940 107.155 10.170 ;
        RECT 107.485 9.940 109.445 10.170 ;
        RECT 111.235 9.940 113.195 10.170 ;
        RECT 113.525 9.940 115.485 10.170 ;
        RECT 117.275 9.940 119.235 10.170 ;
        RECT 119.565 9.940 121.525 10.170 ;
        RECT 123.315 9.940 125.275 10.170 ;
        RECT 125.605 9.940 127.565 10.170 ;
        RECT 128.345 9.480 130.565 39.040 ;
        RECT 8.665 8.890 130.565 9.480 ;
        RECT 7.065 5.690 130.565 8.890 ;
        RECT 135.120 18.845 135.710 41.635 ;
        RECT 136.295 40.485 138.400 41.075 ;
        RECT 136.295 39.315 138.400 39.905 ;
        RECT 146.290 39.315 148.395 41.075 ;
        RECT 136.295 36.975 138.400 38.735 ;
        RECT 146.290 38.145 148.395 38.735 ;
        RECT 146.290 36.975 148.395 37.565 ;
        RECT 136.295 35.805 138.400 36.395 ;
        RECT 136.295 34.635 138.400 35.225 ;
        RECT 146.290 34.635 148.395 36.395 ;
        RECT 136.295 32.295 138.400 34.055 ;
        RECT 146.290 33.465 148.395 34.055 ;
        RECT 143.640 32.295 148.395 32.885 ;
        RECT 136.295 31.125 138.400 31.715 ;
        RECT 136.295 29.955 141.055 30.545 ;
        RECT 146.290 29.955 148.395 31.715 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 136.295 26.445 138.400 28.205 ;
        RECT 146.290 27.615 148.395 29.375 ;
        RECT 136.295 24.105 138.400 25.865 ;
        RECT 146.290 25.275 148.395 27.035 ;
        RECT 136.295 21.765 138.400 23.525 ;
        RECT 146.290 22.935 148.395 24.695 ;
        RECT 136.295 19.425 138.400 21.185 ;
        RECT 146.290 20.595 148.395 22.355 ;
        RECT 141.295 19.425 148.395 20.015 ;
        RECT 148.980 18.845 155.900 104.835 ;
        RECT 167.315 104.330 167.455 105.165 ;
        RECT 171.840 105.165 173.205 105.305 ;
        RECT 171.840 105.120 172.130 105.165 ;
        RECT 173.065 104.625 173.205 105.165 ;
        RECT 174.125 105.105 174.445 105.365 ;
        RECT 174.585 105.305 174.905 105.365 ;
        RECT 175.980 105.305 176.270 105.350 ;
        RECT 174.585 105.165 176.270 105.305 ;
        RECT 174.585 105.105 174.905 105.165 ;
        RECT 175.980 105.120 176.270 105.165 ;
        RECT 177.345 105.305 177.665 105.365 ;
        RECT 177.820 105.305 178.110 105.350 ;
        RECT 177.345 105.165 178.110 105.305 ;
        RECT 177.345 105.105 177.665 105.165 ;
        RECT 177.820 105.120 178.110 105.165 ;
        RECT 181.485 105.105 181.805 105.365 ;
        RECT 182.420 105.305 182.710 105.350 ;
        RECT 185.165 105.305 185.485 105.365 ;
        RECT 182.420 105.165 185.485 105.305 ;
        RECT 182.420 105.120 182.710 105.165 ;
        RECT 185.165 105.105 185.485 105.165 ;
        RECT 185.625 105.105 185.945 105.365 ;
        RECT 186.085 105.105 186.405 105.365 ;
        RECT 190.225 105.305 190.545 105.365 ;
        RECT 190.225 105.165 192.295 105.305 ;
        RECT 190.225 105.105 190.545 105.165 ;
        RECT 189.305 104.965 189.625 105.025 ;
        RECT 184.795 104.825 189.625 104.965 ;
        RECT 178.740 104.625 179.030 104.670 ;
        RECT 182.405 104.625 182.725 104.685 ;
        RECT 184.795 104.670 184.935 104.825 ;
        RECT 189.305 104.765 189.625 104.825 ;
        RECT 191.605 104.765 191.925 105.025 ;
        RECT 192.155 104.965 192.295 105.165 ;
        RECT 195.285 105.105 195.605 105.365 ;
        RECT 195.745 105.305 196.065 105.365 ;
        RECT 199.055 105.350 199.195 105.505 ;
        RECT 199.885 105.505 218.975 105.645 ;
        RECT 199.885 105.445 200.205 105.505 ;
        RECT 198.520 105.305 198.810 105.350 ;
        RECT 195.745 105.165 198.810 105.305 ;
        RECT 195.745 105.105 196.065 105.165 ;
        RECT 198.520 105.120 198.810 105.165 ;
        RECT 198.980 105.120 199.270 105.350 ;
        RECT 203.120 105.305 203.410 105.350 ;
        RECT 203.565 105.305 203.885 105.365 ;
        RECT 203.120 105.165 203.885 105.305 ;
        RECT 203.120 105.120 203.410 105.165 ;
        RECT 203.565 105.105 203.885 105.165 ;
        RECT 204.485 105.105 204.805 105.365 ;
        RECT 208.640 105.305 208.930 105.350 ;
        RECT 212.765 105.305 213.085 105.365 ;
        RECT 208.640 105.165 213.085 105.305 ;
        RECT 208.640 105.120 208.930 105.165 ;
        RECT 212.765 105.105 213.085 105.165 ;
        RECT 213.225 105.105 213.545 105.365 ;
        RECT 214.145 105.305 214.465 105.365 ;
        RECT 216.000 105.305 216.290 105.350 ;
        RECT 214.145 105.165 216.290 105.305 ;
        RECT 214.145 105.105 214.465 105.165 ;
        RECT 216.000 105.120 216.290 105.165 ;
        RECT 218.300 105.305 218.590 105.350 ;
        RECT 218.835 105.305 218.975 105.505 ;
        RECT 224.815 105.505 231.855 105.645 ;
        RECT 224.815 105.350 224.955 105.505 ;
        RECT 231.715 105.365 231.855 105.505 ;
        RECT 232.175 105.505 235.995 105.645 ;
        RECT 218.300 105.165 218.975 105.305 ;
        RECT 218.300 105.120 218.590 105.165 ;
        RECT 220.600 105.120 220.890 105.350 ;
        RECT 222.900 105.305 223.190 105.350 ;
        RECT 221.595 105.165 223.190 105.305 ;
        RECT 192.155 104.825 207.475 104.965 ;
        RECT 173.065 104.485 178.495 104.625 ;
        RECT 178.355 104.345 178.495 104.485 ;
        RECT 178.740 104.485 182.725 104.625 ;
        RECT 178.740 104.440 179.030 104.485 ;
        RECT 182.405 104.425 182.725 104.485 ;
        RECT 184.720 104.440 185.010 104.670 ;
        RECT 187.020 104.625 187.310 104.670 ;
        RECT 191.695 104.625 191.835 104.765 ;
        RECT 187.020 104.485 191.835 104.625 ;
        RECT 199.900 104.625 200.190 104.670 ;
        RECT 203.105 104.625 203.425 104.685 ;
        RECT 199.900 104.485 203.425 104.625 ;
        RECT 187.020 104.440 187.310 104.485 ;
        RECT 199.900 104.440 200.190 104.485 ;
        RECT 203.105 104.425 203.425 104.485 ;
        RECT 167.240 104.285 167.530 104.330 ;
        RECT 173.665 104.285 173.985 104.345 ;
        RECT 167.240 104.145 173.985 104.285 ;
        RECT 167.240 104.100 167.530 104.145 ;
        RECT 173.665 104.085 173.985 104.145 ;
        RECT 178.265 104.085 178.585 104.345 ;
        RECT 202.645 104.285 202.965 104.345 ;
        RECT 206.800 104.285 207.090 104.330 ;
        RECT 202.645 104.145 207.090 104.285 ;
        RECT 207.335 104.285 207.475 104.825 ;
        RECT 209.545 104.765 209.865 105.025 ;
        RECT 212.855 104.965 212.995 105.105 ;
        RECT 219.665 104.965 219.985 105.025 ;
        RECT 220.675 104.965 220.815 105.120 ;
        RECT 212.855 104.825 220.815 104.965 ;
        RECT 219.665 104.765 219.985 104.825 ;
        RECT 220.585 104.625 220.905 104.685 ;
        RECT 221.595 104.625 221.735 105.165 ;
        RECT 222.900 105.120 223.190 105.165 ;
        RECT 224.740 105.120 225.030 105.350 ;
        RECT 229.325 105.105 229.645 105.365 ;
        RECT 230.260 105.120 230.550 105.350 ;
        RECT 221.965 104.965 222.285 105.025 ;
        RECT 230.335 104.965 230.475 105.120 ;
        RECT 231.625 105.105 231.945 105.365 ;
        RECT 232.175 105.350 232.315 105.505 ;
        RECT 235.855 105.365 235.995 105.505 ;
        RECT 244.505 105.505 253.090 105.645 ;
        RECT 244.505 105.445 244.825 105.505 ;
        RECT 252.800 105.460 253.090 105.505 ;
        RECT 257.400 105.645 257.690 105.690 ;
        RECT 261.985 105.645 262.305 105.705 ;
        RECT 257.400 105.505 262.305 105.645 ;
        RECT 262.995 105.645 263.135 105.785 ;
        RECT 274.495 105.645 274.635 105.800 ;
        RECT 276.245 105.785 276.565 106.045 ;
        RECT 276.705 105.985 277.025 106.045 ;
        RECT 279.020 105.985 279.310 106.030 ;
        RECT 276.705 105.845 279.310 105.985 ;
        RECT 276.705 105.785 277.025 105.845 ;
        RECT 279.020 105.800 279.310 105.845 ;
        RECT 283.605 105.785 283.925 106.045 ;
        RECT 286.380 105.800 286.670 106.030 ;
        RECT 290.505 105.985 290.825 106.045 ;
        RECT 291.900 105.985 292.190 106.030 ;
        RECT 290.505 105.845 292.190 105.985 ;
        RECT 286.455 105.645 286.595 105.800 ;
        RECT 290.505 105.785 290.825 105.845 ;
        RECT 291.900 105.800 292.190 105.845 ;
        RECT 297.405 105.785 297.725 106.045 ;
        RECT 299.705 105.785 300.025 106.045 ;
        RECT 300.165 105.785 300.485 106.045 ;
        RECT 302.005 105.985 302.325 106.045 ;
        RECT 305.240 105.985 305.530 106.030 ;
        RECT 302.005 105.845 305.530 105.985 ;
        RECT 302.005 105.785 302.325 105.845 ;
        RECT 305.240 105.800 305.530 105.845 ;
        RECT 307.540 105.800 307.830 106.030 ;
        RECT 262.995 105.505 274.635 105.645 ;
        RECT 279.095 105.505 286.595 105.645 ;
        RECT 299.795 105.645 299.935 105.785 ;
        RECT 307.615 105.645 307.755 105.800 ;
        RECT 299.795 105.505 307.755 105.645 ;
        RECT 257.400 105.460 257.690 105.505 ;
        RECT 261.985 105.445 262.305 105.505 ;
        RECT 279.095 105.365 279.235 105.505 ;
        RECT 232.100 105.120 232.390 105.350 ;
        RECT 233.005 105.305 233.325 105.365 ;
        RECT 234.400 105.305 234.690 105.350 ;
        RECT 233.005 105.165 234.690 105.305 ;
        RECT 233.005 105.105 233.325 105.165 ;
        RECT 234.400 105.120 234.690 105.165 ;
        RECT 235.765 105.105 236.085 105.365 ;
        RECT 236.225 105.305 236.545 105.365 ;
        RECT 237.620 105.305 237.910 105.350 ;
        RECT 236.225 105.165 237.910 105.305 ;
        RECT 236.225 105.105 236.545 105.165 ;
        RECT 237.620 105.120 237.910 105.165 ;
        RECT 241.285 105.305 241.605 105.365 ;
        RECT 241.760 105.305 242.050 105.350 ;
        RECT 241.285 105.165 242.050 105.305 ;
        RECT 241.285 105.105 241.605 105.165 ;
        RECT 241.760 105.120 242.050 105.165 ;
        RECT 242.220 105.305 242.510 105.350 ;
        RECT 245.900 105.305 246.190 105.350 ;
        RECT 246.345 105.305 246.665 105.365 ;
        RECT 242.220 105.165 245.195 105.305 ;
        RECT 242.220 105.120 242.510 105.165 ;
        RECT 245.055 105.025 245.195 105.165 ;
        RECT 245.900 105.165 246.665 105.305 ;
        RECT 245.900 105.120 246.190 105.165 ;
        RECT 246.345 105.105 246.665 105.165 ;
        RECT 250.025 105.105 250.345 105.365 ;
        RECT 254.640 105.305 254.930 105.350 ;
        RECT 251.035 105.165 254.930 105.305 ;
        RECT 236.685 104.965 237.005 105.025 ;
        RECT 242.680 104.965 242.970 105.010 ;
        RECT 244.520 104.965 244.810 105.010 ;
        RECT 221.965 104.825 230.475 104.965 ;
        RECT 230.795 104.825 237.005 104.965 ;
        RECT 221.965 104.765 222.285 104.825 ;
        RECT 230.795 104.625 230.935 104.825 ;
        RECT 236.685 104.765 237.005 104.825 ;
        RECT 238.115 104.825 244.810 104.965 ;
        RECT 220.585 104.485 221.735 104.625 ;
        RECT 225.275 104.485 230.935 104.625 ;
        RECT 233.020 104.625 233.310 104.670 ;
        RECT 237.605 104.625 237.925 104.685 ;
        RECT 233.020 104.485 237.925 104.625 ;
        RECT 220.585 104.425 220.905 104.485 ;
        RECT 225.275 104.285 225.415 104.485 ;
        RECT 233.020 104.440 233.310 104.485 ;
        RECT 237.605 104.425 237.925 104.485 ;
        RECT 207.335 104.145 225.415 104.285 ;
        RECT 225.660 104.285 225.950 104.330 ;
        RECT 230.705 104.285 231.025 104.345 ;
        RECT 225.660 104.145 231.025 104.285 ;
        RECT 202.645 104.085 202.965 104.145 ;
        RECT 206.800 104.100 207.090 104.145 ;
        RECT 225.660 104.100 225.950 104.145 ;
        RECT 230.705 104.085 231.025 104.145 ;
        RECT 232.545 104.285 232.865 104.345 ;
        RECT 238.115 104.285 238.255 104.825 ;
        RECT 242.680 104.780 242.970 104.825 ;
        RECT 244.520 104.780 244.810 104.825 ;
        RECT 244.965 104.765 245.285 105.025 ;
        RECT 245.440 104.965 245.730 105.010 ;
        RECT 251.035 104.965 251.175 105.165 ;
        RECT 254.640 105.120 254.930 105.165 ;
        RECT 245.440 104.825 251.175 104.965 ;
        RECT 245.440 104.780 245.730 104.825 ;
        RECT 244.045 104.625 244.365 104.685 ;
        RECT 245.515 104.625 245.655 104.780 ;
        RECT 251.405 104.765 251.725 105.025 ;
        RECT 254.715 104.965 254.855 105.120 ;
        RECT 259.685 105.105 260.005 105.365 ;
        RECT 262.920 105.305 263.210 105.350 ;
        RECT 260.695 105.165 263.210 105.305 ;
        RECT 257.845 104.965 258.165 105.025 ;
        RECT 254.715 104.825 258.165 104.965 ;
        RECT 257.845 104.765 258.165 104.825 ;
        RECT 244.045 104.485 245.655 104.625 ;
        RECT 251.495 104.625 251.635 104.765 ;
        RECT 260.695 104.685 260.835 105.165 ;
        RECT 262.920 105.120 263.210 105.165 ;
        RECT 267.045 105.105 267.365 105.365 ;
        RECT 270.265 105.105 270.585 105.365 ;
        RECT 271.645 105.305 271.965 105.365 ;
        RECT 273.040 105.305 273.330 105.350 ;
        RECT 271.645 105.165 273.330 105.305 ;
        RECT 271.645 105.105 271.965 105.165 ;
        RECT 273.040 105.120 273.330 105.165 ;
        RECT 275.340 105.120 275.630 105.350 ;
        RECT 268.885 104.965 269.205 105.025 ;
        RECT 275.415 104.965 275.555 105.120 ;
        RECT 277.165 105.105 277.485 105.365 ;
        RECT 279.005 105.105 279.325 105.365 ;
        RECT 279.465 105.305 279.785 105.365 ;
        RECT 280.400 105.305 280.690 105.350 ;
        RECT 279.465 105.165 280.690 105.305 ;
        RECT 279.465 105.105 279.785 105.165 ;
        RECT 280.400 105.120 280.690 105.165 ;
        RECT 281.765 105.305 282.085 105.365 ;
        RECT 282.700 105.305 282.990 105.350 ;
        RECT 281.765 105.165 282.990 105.305 ;
        RECT 281.765 105.105 282.085 105.165 ;
        RECT 282.700 105.120 282.990 105.165 ;
        RECT 284.985 105.105 285.305 105.365 ;
        RECT 287.300 105.305 287.590 105.350 ;
        RECT 288.205 105.305 288.525 105.365 ;
        RECT 287.300 105.165 288.525 105.305 ;
        RECT 287.300 105.120 287.590 105.165 ;
        RECT 288.205 105.105 288.525 105.165 ;
        RECT 289.125 105.105 289.445 105.365 ;
        RECT 290.520 105.120 290.810 105.350 ;
        RECT 293.280 105.120 293.570 105.350 ;
        RECT 282.225 104.965 282.545 105.025 ;
        RECT 290.595 104.965 290.735 105.120 ;
        RECT 268.885 104.825 280.615 104.965 ;
        RECT 268.885 104.765 269.205 104.825 ;
        RECT 280.475 104.685 280.615 104.825 ;
        RECT 282.225 104.825 290.735 104.965 ;
        RECT 293.355 104.965 293.495 105.120 ;
        RECT 294.185 105.105 294.505 105.365 ;
        RECT 298.800 105.120 299.090 105.350 ;
        RECT 296.485 104.965 296.805 105.025 ;
        RECT 293.355 104.825 296.805 104.965 ;
        RECT 282.225 104.765 282.545 104.825 ;
        RECT 296.485 104.765 296.805 104.825 ;
        RECT 258.780 104.625 259.070 104.670 ;
        RECT 251.495 104.485 259.070 104.625 ;
        RECT 244.045 104.425 244.365 104.485 ;
        RECT 258.780 104.440 259.070 104.485 ;
        RECT 260.605 104.425 260.925 104.685 ;
        RECT 280.385 104.425 280.705 104.685 ;
        RECT 281.305 104.625 281.625 104.685 ;
        RECT 288.220 104.625 288.510 104.670 ;
        RECT 295.120 104.625 295.410 104.670 ;
        RECT 281.305 104.485 288.510 104.625 ;
        RECT 281.305 104.425 281.625 104.485 ;
        RECT 288.220 104.440 288.510 104.485 ;
        RECT 289.215 104.485 295.410 104.625 ;
        RECT 298.875 104.625 299.015 105.120 ;
        RECT 301.085 105.105 301.405 105.365 ;
        RECT 301.560 105.120 301.850 105.350 ;
        RECT 300.165 104.965 300.485 105.025 ;
        RECT 301.635 104.965 301.775 105.120 ;
        RECT 304.765 105.105 305.085 105.365 ;
        RECT 308.445 105.105 308.765 105.365 ;
        RECT 300.165 104.825 301.775 104.965 ;
        RECT 300.165 104.765 300.485 104.825 ;
        RECT 302.925 104.625 303.245 104.685 ;
        RECT 298.875 104.485 303.245 104.625 ;
        RECT 232.545 104.145 238.255 104.285 ;
        RECT 239.920 104.285 240.210 104.330 ;
        RECT 240.365 104.285 240.685 104.345 ;
        RECT 239.920 104.145 240.685 104.285 ;
        RECT 232.545 104.085 232.865 104.145 ;
        RECT 239.920 104.100 240.210 104.145 ;
        RECT 240.365 104.085 240.685 104.145 ;
        RECT 247.725 104.085 248.045 104.345 ;
        RECT 256.005 104.285 256.325 104.345 ;
        RECT 266.140 104.285 266.430 104.330 ;
        RECT 256.005 104.145 266.430 104.285 ;
        RECT 256.005 104.085 256.325 104.145 ;
        RECT 266.140 104.100 266.430 104.145 ;
        RECT 272.105 104.285 272.425 104.345 ;
        RECT 281.780 104.285 282.070 104.330 ;
        RECT 272.105 104.145 282.070 104.285 ;
        RECT 272.105 104.085 272.425 104.145 ;
        RECT 281.780 104.100 282.070 104.145 ;
        RECT 285.905 104.285 286.225 104.345 ;
        RECT 289.215 104.285 289.355 104.485 ;
        RECT 295.120 104.440 295.410 104.485 ;
        RECT 302.925 104.425 303.245 104.485 ;
        RECT 285.905 104.145 289.355 104.285 ;
        RECT 285.905 104.085 286.225 104.145 ;
        RECT 289.585 104.085 289.905 104.345 ;
        RECT 302.465 104.085 302.785 104.345 ;
        RECT 162.095 103.465 311.135 103.945 ;
        RECT 165.845 103.265 166.165 103.325 ;
        RECT 175.520 103.265 175.810 103.310 ;
        RECT 165.845 103.125 175.810 103.265 ;
        RECT 165.845 103.065 166.165 103.125 ;
        RECT 175.520 103.080 175.810 103.125 ;
        RECT 175.965 103.265 176.285 103.325 ;
        RECT 180.120 103.265 180.410 103.310 ;
        RECT 190.225 103.265 190.545 103.325 ;
        RECT 175.965 103.125 180.410 103.265 ;
        RECT 175.965 103.065 176.285 103.125 ;
        RECT 180.120 103.080 180.410 103.125 ;
        RECT 180.655 103.125 190.545 103.265 ;
        RECT 166.270 102.925 166.560 102.970 ;
        RECT 168.160 102.925 168.450 102.970 ;
        RECT 171.280 102.925 171.570 102.970 ;
        RECT 166.270 102.785 171.570 102.925 ;
        RECT 166.270 102.740 166.560 102.785 ;
        RECT 168.160 102.740 168.450 102.785 ;
        RECT 171.280 102.740 171.570 102.785 ;
        RECT 172.745 102.585 173.065 102.645 ;
        RECT 172.375 102.445 173.065 102.585 ;
        RECT 165.385 102.045 165.705 102.305 ;
        RECT 165.865 102.245 166.155 102.290 ;
        RECT 167.700 102.245 167.990 102.290 ;
        RECT 171.280 102.245 171.570 102.290 ;
        RECT 172.375 102.265 172.515 102.445 ;
        RECT 172.745 102.385 173.065 102.445 ;
        RECT 174.140 102.585 174.430 102.630 ;
        RECT 174.140 102.445 177.575 102.585 ;
        RECT 174.140 102.400 174.430 102.445 ;
        RECT 177.435 102.290 177.575 102.445 ;
        RECT 178.725 102.385 179.045 102.645 ;
        RECT 165.865 102.105 171.570 102.245 ;
        RECT 165.865 102.060 166.155 102.105 ;
        RECT 167.700 102.060 167.990 102.105 ;
        RECT 171.280 102.060 171.570 102.105 ;
        RECT 166.765 101.705 167.085 101.965 ;
        RECT 172.360 101.950 172.650 102.265 ;
        RECT 177.360 102.245 177.650 102.290 ;
        RECT 180.655 102.245 180.795 103.125 ;
        RECT 190.225 103.065 190.545 103.125 ;
        RECT 199.885 103.065 200.205 103.325 ;
        RECT 204.040 103.265 204.330 103.310 ;
        RECT 205.405 103.265 205.725 103.325 ;
        RECT 204.040 103.125 205.725 103.265 ;
        RECT 204.040 103.080 204.330 103.125 ;
        RECT 205.405 103.065 205.725 103.125 ;
        RECT 210.005 103.265 210.325 103.325 ;
        RECT 215.080 103.265 215.370 103.310 ;
        RECT 210.005 103.125 215.370 103.265 ;
        RECT 210.005 103.065 210.325 103.125 ;
        RECT 215.080 103.080 215.370 103.125 ;
        RECT 226.105 103.265 226.425 103.325 ;
        RECT 236.225 103.265 236.545 103.325 ;
        RECT 226.105 103.125 236.545 103.265 ;
        RECT 226.105 103.065 226.425 103.125 ;
        RECT 236.225 103.065 236.545 103.125 ;
        RECT 236.685 103.265 237.005 103.325 ;
        RECT 246.805 103.265 247.125 103.325 ;
        RECT 248.200 103.265 248.490 103.310 ;
        RECT 236.685 103.125 245.195 103.265 ;
        RECT 236.685 103.065 237.005 103.125 ;
        RECT 182.370 102.925 182.660 102.970 ;
        RECT 184.260 102.925 184.550 102.970 ;
        RECT 187.380 102.925 187.670 102.970 ;
        RECT 182.370 102.785 187.670 102.925 ;
        RECT 182.370 102.740 182.660 102.785 ;
        RECT 184.260 102.740 184.550 102.785 ;
        RECT 187.380 102.740 187.670 102.785 ;
        RECT 192.030 102.925 192.320 102.970 ;
        RECT 193.920 102.925 194.210 102.970 ;
        RECT 197.040 102.925 197.330 102.970 ;
        RECT 192.030 102.785 197.330 102.925 ;
        RECT 192.030 102.740 192.320 102.785 ;
        RECT 193.920 102.740 194.210 102.785 ;
        RECT 197.040 102.740 197.330 102.785 ;
        RECT 206.290 102.925 206.580 102.970 ;
        RECT 208.180 102.925 208.470 102.970 ;
        RECT 211.300 102.925 211.590 102.970 ;
        RECT 206.290 102.785 211.590 102.925 ;
        RECT 206.290 102.740 206.580 102.785 ;
        RECT 208.180 102.740 208.470 102.785 ;
        RECT 211.300 102.740 211.590 102.785 ;
        RECT 212.765 102.925 213.085 102.985 ;
        RECT 214.160 102.925 214.450 102.970 ;
        RECT 212.765 102.785 214.450 102.925 ;
        RECT 212.765 102.725 213.085 102.785 ;
        RECT 214.160 102.740 214.450 102.785 ;
        RECT 218.250 102.925 218.540 102.970 ;
        RECT 220.140 102.925 220.430 102.970 ;
        RECT 223.260 102.925 223.550 102.970 ;
        RECT 218.250 102.785 223.550 102.925 ;
        RECT 218.250 102.740 218.540 102.785 ;
        RECT 220.140 102.740 220.430 102.785 ;
        RECT 223.260 102.740 223.550 102.785 ;
        RECT 227.910 102.925 228.200 102.970 ;
        RECT 229.800 102.925 230.090 102.970 ;
        RECT 232.920 102.925 233.210 102.970 ;
        RECT 227.910 102.785 233.210 102.925 ;
        RECT 227.910 102.740 228.200 102.785 ;
        RECT 229.800 102.740 230.090 102.785 ;
        RECT 232.920 102.740 233.210 102.785 ;
        RECT 239.410 102.925 239.700 102.970 ;
        RECT 241.300 102.925 241.590 102.970 ;
        RECT 244.420 102.925 244.710 102.970 ;
        RECT 239.410 102.785 244.710 102.925 ;
        RECT 245.055 102.925 245.195 103.125 ;
        RECT 246.805 103.125 248.490 103.265 ;
        RECT 246.805 103.065 247.125 103.125 ;
        RECT 248.200 103.080 248.490 103.125 ;
        RECT 249.105 103.265 249.425 103.325 ;
        RECT 253.260 103.265 253.550 103.310 ;
        RECT 249.105 103.125 253.550 103.265 ;
        RECT 249.105 103.065 249.425 103.125 ;
        RECT 253.260 103.080 253.550 103.125 ;
        RECT 256.005 103.265 256.325 103.325 ;
        RECT 258.765 103.265 259.085 103.325 ;
        RECT 266.140 103.265 266.430 103.310 ;
        RECT 256.005 103.125 257.615 103.265 ;
        RECT 256.005 103.065 256.325 103.125 ;
        RECT 245.055 102.785 257.155 102.925 ;
        RECT 239.410 102.740 239.700 102.785 ;
        RECT 241.300 102.740 241.590 102.785 ;
        RECT 244.420 102.740 244.710 102.785 ;
        RECT 181.500 102.585 181.790 102.630 ;
        RECT 183.325 102.585 183.645 102.645 ;
        RECT 181.500 102.445 183.645 102.585 ;
        RECT 181.500 102.400 181.790 102.445 ;
        RECT 183.325 102.385 183.645 102.445 ;
        RECT 185.625 102.585 185.945 102.645 ;
        RECT 190.225 102.585 190.545 102.645 ;
        RECT 185.625 102.445 190.545 102.585 ;
        RECT 185.625 102.385 185.945 102.445 ;
        RECT 190.225 102.385 190.545 102.445 ;
        RECT 191.160 102.585 191.450 102.630 ;
        RECT 205.405 102.585 205.725 102.645 ;
        RECT 217.380 102.585 217.670 102.630 ;
        RECT 227.040 102.585 227.330 102.630 ;
        RECT 191.160 102.445 227.330 102.585 ;
        RECT 191.160 102.400 191.450 102.445 ;
        RECT 200.895 102.305 201.035 102.445 ;
        RECT 205.405 102.385 205.725 102.445 ;
        RECT 217.380 102.400 217.670 102.445 ;
        RECT 227.040 102.400 227.330 102.445 ;
        RECT 235.765 102.585 236.085 102.645 ;
        RECT 238.540 102.585 238.830 102.630 ;
        RECT 235.765 102.445 237.375 102.585 ;
        RECT 235.765 102.385 236.085 102.445 ;
        RECT 177.360 102.105 180.795 102.245 ;
        RECT 177.360 102.060 177.650 102.105 ;
        RECT 181.040 102.060 181.330 102.290 ;
        RECT 181.965 102.245 182.255 102.290 ;
        RECT 183.800 102.245 184.090 102.290 ;
        RECT 187.380 102.245 187.670 102.290 ;
        RECT 181.965 102.105 187.670 102.245 ;
        RECT 181.965 102.060 182.255 102.105 ;
        RECT 183.800 102.060 184.090 102.105 ;
        RECT 187.380 102.060 187.670 102.105 ;
        RECT 169.060 101.905 169.710 101.950 ;
        RECT 172.360 101.905 172.950 101.950 ;
        RECT 169.060 101.765 172.950 101.905 ;
        RECT 181.115 101.905 181.255 102.060 ;
        RECT 182.405 101.905 182.725 101.965 ;
        RECT 181.115 101.765 182.725 101.905 ;
        RECT 169.060 101.720 169.710 101.765 ;
        RECT 172.660 101.720 172.950 101.765 ;
        RECT 182.405 101.705 182.725 101.765 ;
        RECT 182.865 101.705 183.185 101.965 ;
        RECT 188.460 101.950 188.750 102.265 ;
        RECT 191.625 102.245 191.915 102.290 ;
        RECT 193.460 102.245 193.750 102.290 ;
        RECT 197.040 102.245 197.330 102.290 ;
        RECT 191.625 102.105 197.330 102.245 ;
        RECT 191.625 102.060 191.915 102.105 ;
        RECT 193.460 102.060 193.750 102.105 ;
        RECT 197.040 102.060 197.330 102.105 ;
        RECT 185.160 101.905 185.810 101.950 ;
        RECT 188.460 101.905 189.050 101.950 ;
        RECT 185.160 101.765 191.835 101.905 ;
        RECT 185.160 101.720 185.810 101.765 ;
        RECT 188.760 101.720 189.050 101.765 ;
        RECT 191.695 101.625 191.835 101.765 ;
        RECT 192.525 101.705 192.845 101.965 ;
        RECT 194.825 101.950 195.145 101.965 ;
        RECT 198.120 101.950 198.410 102.265 ;
        RECT 200.805 102.045 201.125 102.305 ;
        RECT 201.740 102.245 202.030 102.290 ;
        RECT 202.645 102.245 202.965 102.305 ;
        RECT 201.740 102.105 202.965 102.245 ;
        RECT 201.740 102.060 202.030 102.105 ;
        RECT 202.645 102.045 202.965 102.105 ;
        RECT 203.105 102.045 203.425 102.305 ;
        RECT 205.885 102.245 206.175 102.290 ;
        RECT 207.720 102.245 208.010 102.290 ;
        RECT 211.300 102.245 211.590 102.290 ;
        RECT 205.885 102.105 211.590 102.245 ;
        RECT 205.885 102.060 206.175 102.105 ;
        RECT 207.720 102.060 208.010 102.105 ;
        RECT 211.300 102.060 211.590 102.105 ;
        RECT 209.085 101.950 209.405 101.965 ;
        RECT 212.380 101.950 212.670 102.265 ;
        RECT 217.845 102.245 218.135 102.290 ;
        RECT 219.680 102.245 219.970 102.290 ;
        RECT 223.260 102.245 223.550 102.290 ;
        RECT 217.845 102.105 223.550 102.245 ;
        RECT 217.845 102.060 218.135 102.105 ;
        RECT 219.680 102.060 219.970 102.105 ;
        RECT 223.260 102.060 223.550 102.105 ;
        RECT 194.820 101.905 195.470 101.950 ;
        RECT 198.120 101.905 198.710 101.950 ;
        RECT 206.800 101.905 207.090 101.950 ;
        RECT 209.080 101.905 209.730 101.950 ;
        RECT 212.380 101.905 212.970 101.950 ;
        RECT 194.820 101.765 198.710 101.905 ;
        RECT 194.820 101.720 195.470 101.765 ;
        RECT 198.420 101.720 198.710 101.765 ;
        RECT 202.735 101.765 207.090 101.905 ;
        RECT 194.825 101.705 195.145 101.720 ;
        RECT 177.820 101.565 178.110 101.610 ;
        RECT 190.225 101.565 190.545 101.625 ;
        RECT 177.820 101.425 190.545 101.565 ;
        RECT 177.820 101.380 178.110 101.425 ;
        RECT 190.225 101.365 190.545 101.425 ;
        RECT 191.605 101.365 191.925 101.625 ;
        RECT 202.735 101.610 202.875 101.765 ;
        RECT 206.800 101.720 207.090 101.765 ;
        RECT 208.715 101.765 212.970 101.905 ;
        RECT 202.660 101.380 202.950 101.610 ;
        RECT 208.715 101.565 208.855 101.765 ;
        RECT 209.080 101.720 209.730 101.765 ;
        RECT 212.680 101.720 212.970 101.765 ;
        RECT 214.605 101.905 214.925 101.965 ;
        RECT 216.460 101.905 216.750 101.950 ;
        RECT 214.605 101.765 216.750 101.905 ;
        RECT 209.085 101.705 209.405 101.720 ;
        RECT 214.605 101.705 214.925 101.765 ;
        RECT 216.460 101.720 216.750 101.765 ;
        RECT 218.760 101.905 219.050 101.950 ;
        RECT 219.205 101.905 219.525 101.965 ;
        RECT 224.340 101.950 224.630 102.265 ;
        RECT 227.505 102.245 227.795 102.290 ;
        RECT 229.340 102.245 229.630 102.290 ;
        RECT 232.920 102.245 233.210 102.290 ;
        RECT 227.505 102.105 233.210 102.245 ;
        RECT 227.505 102.060 227.795 102.105 ;
        RECT 229.340 102.060 229.630 102.105 ;
        RECT 232.920 102.060 233.210 102.105 ;
        RECT 218.760 101.765 219.525 101.905 ;
        RECT 218.760 101.720 219.050 101.765 ;
        RECT 219.205 101.705 219.525 101.765 ;
        RECT 221.040 101.905 221.690 101.950 ;
        RECT 224.340 101.905 224.930 101.950 ;
        RECT 221.040 101.765 227.715 101.905 ;
        RECT 221.040 101.720 221.690 101.765 ;
        RECT 224.640 101.720 224.930 101.765 ;
        RECT 225.275 101.565 225.415 101.765 ;
        RECT 208.715 101.425 225.415 101.565 ;
        RECT 227.575 101.565 227.715 101.765 ;
        RECT 228.405 101.705 228.725 101.965 ;
        RECT 234.000 101.950 234.290 102.265 ;
        RECT 230.700 101.905 231.350 101.950 ;
        RECT 234.000 101.905 234.590 101.950 ;
        RECT 237.235 101.905 237.375 102.445 ;
        RECT 238.540 102.445 252.555 102.585 ;
        RECT 238.540 102.400 238.830 102.445 ;
        RECT 252.415 102.305 252.555 102.445 ;
        RECT 252.875 102.445 255.775 102.585 ;
        RECT 252.875 102.305 253.015 102.445 ;
        RECT 237.605 102.045 237.925 102.305 ;
        RECT 239.005 102.245 239.295 102.290 ;
        RECT 240.840 102.245 241.130 102.290 ;
        RECT 244.420 102.245 244.710 102.290 ;
        RECT 239.005 102.105 244.710 102.245 ;
        RECT 239.005 102.060 239.295 102.105 ;
        RECT 240.840 102.060 241.130 102.105 ;
        RECT 244.420 102.060 244.710 102.105 ;
        RECT 230.700 101.765 236.915 101.905 ;
        RECT 237.235 101.765 237.835 101.905 ;
        RECT 230.700 101.720 231.350 101.765 ;
        RECT 234.300 101.720 234.590 101.765 ;
        RECT 234.935 101.565 235.075 101.765 ;
        RECT 236.775 101.610 236.915 101.765 ;
        RECT 237.695 101.625 237.835 101.765 ;
        RECT 239.905 101.705 240.225 101.965 ;
        RECT 245.500 101.950 245.790 102.265 ;
        RECT 247.725 102.245 248.045 102.305 ;
        RECT 251.420 102.245 251.710 102.290 ;
        RECT 247.725 102.105 251.710 102.245 ;
        RECT 247.725 102.045 248.045 102.105 ;
        RECT 251.420 102.060 251.710 102.105 ;
        RECT 252.325 102.045 252.645 102.305 ;
        RECT 252.785 102.045 253.105 102.305 ;
        RECT 253.245 102.245 253.565 102.305 ;
        RECT 255.635 102.290 255.775 102.445 ;
        RECT 257.015 102.290 257.155 102.785 ;
        RECT 257.475 102.290 257.615 103.125 ;
        RECT 258.765 103.125 266.430 103.265 ;
        RECT 258.765 103.065 259.085 103.125 ;
        RECT 266.140 103.080 266.430 103.125 ;
        RECT 268.885 103.065 269.205 103.325 ;
        RECT 282.225 103.065 282.545 103.325 ;
        RECT 289.585 103.265 289.905 103.325 ;
        RECT 282.775 103.125 289.905 103.265 ;
        RECT 258.320 102.740 258.610 102.970 ;
        RECT 260.605 102.925 260.925 102.985 ;
        RECT 259.315 102.785 260.925 102.925 ;
        RECT 254.180 102.245 254.470 102.290 ;
        RECT 253.245 102.105 254.470 102.245 ;
        RECT 253.245 102.045 253.565 102.105 ;
        RECT 254.180 102.060 254.470 102.105 ;
        RECT 255.560 102.060 255.850 102.290 ;
        RECT 256.940 102.060 257.230 102.290 ;
        RECT 257.400 102.060 257.690 102.290 ;
        RECT 258.395 102.245 258.535 102.740 ;
        RECT 259.315 102.290 259.455 102.785 ;
        RECT 260.605 102.725 260.925 102.785 ;
        RECT 262.000 102.925 262.290 102.970 ;
        RECT 263.365 102.925 263.685 102.985 ;
        RECT 262.000 102.785 263.685 102.925 ;
        RECT 262.000 102.740 262.290 102.785 ;
        RECT 263.365 102.725 263.685 102.785 ;
        RECT 265.220 102.925 265.510 102.970 ;
        RECT 269.805 102.925 270.125 102.985 ;
        RECT 265.220 102.785 270.125 102.925 ;
        RECT 265.220 102.740 265.510 102.785 ;
        RECT 269.805 102.725 270.125 102.785 ;
        RECT 271.760 102.925 272.050 102.970 ;
        RECT 274.880 102.925 275.170 102.970 ;
        RECT 276.770 102.925 277.060 102.970 ;
        RECT 282.775 102.925 282.915 103.125 ;
        RECT 289.585 103.065 289.905 103.125 ;
        RECT 290.045 103.265 290.365 103.325 ;
        RECT 293.740 103.265 294.030 103.310 ;
        RECT 290.045 103.125 294.030 103.265 ;
        RECT 290.045 103.065 290.365 103.125 ;
        RECT 293.740 103.080 294.030 103.125 ;
        RECT 295.105 103.265 295.425 103.325 ;
        RECT 305.240 103.265 305.530 103.310 ;
        RECT 295.105 103.125 305.530 103.265 ;
        RECT 295.105 103.065 295.425 103.125 ;
        RECT 305.240 103.080 305.530 103.125 ;
        RECT 271.760 102.785 277.060 102.925 ;
        RECT 271.760 102.740 272.050 102.785 ;
        RECT 274.880 102.740 275.170 102.785 ;
        RECT 276.770 102.740 277.060 102.785 ;
        RECT 278.635 102.785 282.915 102.925 ;
        RECT 267.965 102.585 268.285 102.645 ;
        RECT 259.775 102.445 262.675 102.585 ;
        RECT 258.780 102.245 259.070 102.290 ;
        RECT 258.395 102.105 259.070 102.245 ;
        RECT 258.780 102.060 259.070 102.105 ;
        RECT 259.245 102.060 259.535 102.290 ;
        RECT 242.200 101.905 242.850 101.950 ;
        RECT 245.500 101.905 246.090 101.950 ;
        RECT 248.645 101.905 248.965 101.965 ;
        RECT 242.200 101.765 248.965 101.905 ;
        RECT 242.200 101.720 242.850 101.765 ;
        RECT 245.800 101.720 246.090 101.765 ;
        RECT 248.645 101.705 248.965 101.765 ;
        RECT 249.565 101.705 249.885 101.965 ;
        RECT 250.025 101.905 250.345 101.965 ;
        RECT 254.625 101.905 254.945 101.965 ;
        RECT 256.480 101.905 256.770 101.950 ;
        RECT 250.025 101.765 253.475 101.905 ;
        RECT 250.025 101.705 250.345 101.765 ;
        RECT 227.575 101.425 235.075 101.565 ;
        RECT 236.700 101.380 236.990 101.610 ;
        RECT 237.605 101.365 237.925 101.625 ;
        RECT 244.965 101.565 245.285 101.625 ;
        RECT 247.280 101.565 247.570 101.610 ;
        RECT 250.115 101.565 250.255 101.705 ;
        RECT 244.965 101.425 250.255 101.565 ;
        RECT 244.965 101.365 245.285 101.425 ;
        RECT 247.280 101.380 247.570 101.425 ;
        RECT 250.485 101.365 250.805 101.625 ;
        RECT 253.335 101.565 253.475 101.765 ;
        RECT 254.625 101.765 256.770 101.905 ;
        RECT 257.015 101.905 257.155 102.060 ;
        RECT 259.775 101.905 259.915 102.445 ;
        RECT 261.065 102.290 261.385 102.305 ;
        RECT 262.535 102.290 262.675 102.445 ;
        RECT 267.135 102.445 268.285 102.585 ;
        RECT 261.065 102.245 261.395 102.290 ;
        RECT 261.065 102.105 261.580 102.245 ;
        RECT 261.065 102.060 261.395 102.105 ;
        RECT 262.460 102.060 262.750 102.290 ;
        RECT 262.995 102.105 264.055 102.245 ;
        RECT 261.065 102.045 261.385 102.060 ;
        RECT 257.015 101.765 259.915 101.905 ;
        RECT 254.625 101.705 254.945 101.765 ;
        RECT 256.480 101.720 256.770 101.765 ;
        RECT 260.145 101.705 260.465 101.965 ;
        RECT 260.620 101.905 260.910 101.950 ;
        RECT 262.995 101.905 263.135 102.105 ;
        RECT 263.915 101.950 264.055 102.105 ;
        RECT 264.285 102.045 264.605 102.305 ;
        RECT 267.135 102.290 267.275 102.445 ;
        RECT 267.965 102.385 268.285 102.445 ;
        RECT 276.260 102.585 276.550 102.630 ;
        RECT 278.635 102.585 278.775 102.785 ;
        RECT 283.145 102.725 283.465 102.985 ;
        RECT 285.870 102.925 286.160 102.970 ;
        RECT 287.760 102.925 288.050 102.970 ;
        RECT 290.880 102.925 291.170 102.970 ;
        RECT 285.870 102.785 291.170 102.925 ;
        RECT 285.870 102.740 286.160 102.785 ;
        RECT 287.760 102.740 288.050 102.785 ;
        RECT 290.880 102.740 291.170 102.785 ;
        RECT 297.520 102.925 297.810 102.970 ;
        RECT 300.640 102.925 300.930 102.970 ;
        RECT 302.530 102.925 302.820 102.970 ;
        RECT 297.520 102.785 302.820 102.925 ;
        RECT 297.520 102.740 297.810 102.785 ;
        RECT 300.640 102.740 300.930 102.785 ;
        RECT 302.530 102.740 302.820 102.785 ;
        RECT 276.260 102.445 278.775 102.585 ;
        RECT 276.260 102.400 276.550 102.445 ;
        RECT 279.465 102.385 279.785 102.645 ;
        RECT 279.940 102.585 280.230 102.630 ;
        RECT 280.845 102.585 281.165 102.645 ;
        RECT 288.205 102.585 288.525 102.645 ;
        RECT 279.940 102.445 281.165 102.585 ;
        RECT 279.940 102.400 280.230 102.445 ;
        RECT 280.845 102.385 281.165 102.445 ;
        RECT 284.615 102.445 288.525 102.585 ;
        RECT 267.060 102.060 267.350 102.290 ;
        RECT 270.680 101.950 270.970 102.265 ;
        RECT 271.760 102.245 272.050 102.290 ;
        RECT 275.340 102.245 275.630 102.290 ;
        RECT 277.175 102.245 277.465 102.290 ;
        RECT 271.760 102.105 277.465 102.245 ;
        RECT 271.760 102.060 272.050 102.105 ;
        RECT 275.340 102.060 275.630 102.105 ;
        RECT 277.175 102.060 277.465 102.105 ;
        RECT 277.625 102.045 277.945 102.305 ;
        RECT 283.605 102.245 283.925 102.305 ;
        RECT 280.015 102.105 283.925 102.245 ;
        RECT 260.620 101.765 263.135 101.905 ;
        RECT 260.620 101.720 260.910 101.765 ;
        RECT 263.380 101.720 263.670 101.950 ;
        RECT 263.840 101.905 264.130 101.950 ;
        RECT 270.380 101.905 270.970 101.950 ;
        RECT 273.620 101.905 274.270 101.950 ;
        RECT 274.865 101.905 275.185 101.965 ;
        RECT 280.015 101.905 280.155 102.105 ;
        RECT 283.605 102.045 283.925 102.105 ;
        RECT 284.065 102.045 284.385 102.305 ;
        RECT 263.840 101.765 269.805 101.905 ;
        RECT 263.840 101.720 264.130 101.765 ;
        RECT 256.925 101.565 257.245 101.625 ;
        RECT 253.335 101.425 257.245 101.565 ;
        RECT 256.925 101.365 257.245 101.425 ;
        RECT 257.385 101.565 257.705 101.625 ;
        RECT 263.455 101.565 263.595 101.720 ;
        RECT 257.385 101.425 263.595 101.565 ;
        RECT 269.665 101.565 269.805 101.765 ;
        RECT 270.380 101.765 280.155 101.905 ;
        RECT 270.380 101.720 270.670 101.765 ;
        RECT 273.620 101.720 274.270 101.765 ;
        RECT 274.865 101.705 275.185 101.765 ;
        RECT 280.385 101.705 280.705 101.965 ;
        RECT 284.615 101.565 284.755 102.445 ;
        RECT 288.205 102.385 288.525 102.445 ;
        RECT 285.000 102.060 285.290 102.290 ;
        RECT 285.465 102.245 285.755 102.290 ;
        RECT 287.300 102.245 287.590 102.290 ;
        RECT 290.880 102.245 291.170 102.290 ;
        RECT 285.465 102.105 291.170 102.245 ;
        RECT 285.465 102.060 285.755 102.105 ;
        RECT 287.300 102.060 287.590 102.105 ;
        RECT 290.880 102.060 291.170 102.105 ;
        RECT 269.665 101.425 284.755 101.565 ;
        RECT 285.075 101.565 285.215 102.060 ;
        RECT 286.365 101.705 286.685 101.965 ;
        RECT 287.745 101.905 288.065 101.965 ;
        RECT 291.960 101.950 292.250 102.265 ;
        RECT 288.660 101.905 289.310 101.950 ;
        RECT 291.960 101.905 292.550 101.950 ;
        RECT 287.745 101.765 292.550 101.905 ;
        RECT 287.745 101.705 288.065 101.765 ;
        RECT 288.660 101.720 289.310 101.765 ;
        RECT 292.260 101.720 292.550 101.765 ;
        RECT 295.105 101.905 295.425 101.965 ;
        RECT 296.440 101.950 296.730 102.265 ;
        RECT 297.520 102.245 297.810 102.290 ;
        RECT 301.100 102.245 301.390 102.290 ;
        RECT 302.935 102.245 303.225 102.290 ;
        RECT 297.520 102.105 303.225 102.245 ;
        RECT 297.520 102.060 297.810 102.105 ;
        RECT 301.100 102.060 301.390 102.105 ;
        RECT 302.935 102.060 303.225 102.105 ;
        RECT 303.385 102.045 303.705 102.305 ;
        RECT 304.320 102.060 304.610 102.290 ;
        RECT 296.140 101.905 296.730 101.950 ;
        RECT 299.380 101.905 300.030 101.950 ;
        RECT 295.105 101.765 300.030 101.905 ;
        RECT 295.105 101.705 295.425 101.765 ;
        RECT 296.140 101.720 296.430 101.765 ;
        RECT 299.380 101.720 300.030 101.765 ;
        RECT 302.005 101.705 302.325 101.965 ;
        RECT 302.465 101.905 302.785 101.965 ;
        RECT 304.395 101.905 304.535 102.060 ;
        RECT 302.465 101.765 304.535 101.905 ;
        RECT 302.465 101.705 302.785 101.765 ;
        RECT 307.525 101.705 307.845 101.965 ;
        RECT 309.365 101.705 309.685 101.965 ;
        RECT 286.825 101.565 287.145 101.625 ;
        RECT 285.075 101.425 287.145 101.565 ;
        RECT 257.385 101.365 257.705 101.425 ;
        RECT 286.825 101.365 287.145 101.425 ;
        RECT 288.205 101.565 288.525 101.625 ;
        RECT 294.660 101.565 294.950 101.610 ;
        RECT 303.845 101.565 304.165 101.625 ;
        RECT 288.205 101.425 304.165 101.565 ;
        RECT 288.205 101.365 288.525 101.425 ;
        RECT 294.660 101.380 294.950 101.425 ;
        RECT 303.845 101.365 304.165 101.425 ;
        RECT 162.095 100.745 311.935 101.225 ;
        RECT 166.320 100.545 166.610 100.590 ;
        RECT 166.765 100.545 167.085 100.605 ;
        RECT 166.320 100.405 167.085 100.545 ;
        RECT 166.320 100.360 166.610 100.405 ;
        RECT 166.765 100.345 167.085 100.405 ;
        RECT 167.240 100.545 167.530 100.590 ;
        RECT 168.145 100.545 168.465 100.605 ;
        RECT 187.005 100.545 187.325 100.605 ;
        RECT 199.440 100.545 199.730 100.590 ;
        RECT 200.345 100.545 200.665 100.605 ;
        RECT 167.240 100.405 168.465 100.545 ;
        RECT 167.240 100.360 167.530 100.405 ;
        RECT 168.145 100.345 168.465 100.405 ;
        RECT 168.695 100.405 188.615 100.545 ;
        RECT 165.400 99.865 165.690 99.910 ;
        RECT 165.845 99.865 166.165 99.925 ;
        RECT 165.400 99.725 166.165 99.865 ;
        RECT 165.400 99.680 165.690 99.725 ;
        RECT 165.845 99.665 166.165 99.725 ;
        RECT 168.145 99.665 168.465 99.925 ;
        RECT 168.695 99.910 168.835 100.405 ;
        RECT 187.005 100.345 187.325 100.405 ;
        RECT 172.745 100.250 173.065 100.265 ;
        RECT 172.280 100.205 173.065 100.250 ;
        RECT 175.880 100.205 176.170 100.250 ;
        RECT 172.280 100.065 176.170 100.205 ;
        RECT 172.280 100.020 173.065 100.065 ;
        RECT 172.745 100.005 173.065 100.020 ;
        RECT 175.580 100.020 176.170 100.065 ;
        RECT 179.660 100.205 179.950 100.250 ;
        RECT 179.660 100.065 185.395 100.205 ;
        RECT 179.660 100.020 179.950 100.065 ;
        RECT 168.620 99.680 168.910 99.910 ;
        RECT 169.085 99.865 169.375 99.910 ;
        RECT 170.920 99.865 171.210 99.910 ;
        RECT 174.500 99.865 174.790 99.910 ;
        RECT 169.085 99.725 174.790 99.865 ;
        RECT 169.085 99.680 169.375 99.725 ;
        RECT 170.920 99.680 171.210 99.725 ;
        RECT 174.500 99.680 174.790 99.725 ;
        RECT 175.580 99.705 175.870 100.020 ;
        RECT 169.985 99.325 170.305 99.585 ;
        RECT 177.360 99.525 177.650 99.570 ;
        RECT 179.735 99.525 179.875 100.020 ;
        RECT 185.255 99.925 185.395 100.065 ;
        RECT 185.625 100.005 185.945 100.265 ;
        RECT 181.960 99.865 182.250 99.910 ;
        RECT 181.960 99.725 184.015 99.865 ;
        RECT 181.960 99.680 182.250 99.725 ;
        RECT 177.360 99.385 179.875 99.525 ;
        RECT 177.360 99.340 177.650 99.385 ;
        RECT 180.120 99.340 180.410 99.570 ;
        RECT 181.040 99.340 181.330 99.570 ;
        RECT 169.490 99.185 169.780 99.230 ;
        RECT 171.380 99.185 171.670 99.230 ;
        RECT 174.500 99.185 174.790 99.230 ;
        RECT 169.490 99.045 174.790 99.185 ;
        RECT 169.490 99.000 169.780 99.045 ;
        RECT 171.380 99.000 171.670 99.045 ;
        RECT 174.500 99.000 174.790 99.045 ;
        RECT 179.185 99.185 179.505 99.245 ;
        RECT 180.195 99.185 180.335 99.340 ;
        RECT 179.185 99.045 180.335 99.185 ;
        RECT 179.185 98.985 179.505 99.045 ;
        RECT 177.805 98.645 178.125 98.905 ;
        RECT 178.725 98.845 179.045 98.905 ;
        RECT 181.115 98.845 181.255 99.340 ;
        RECT 182.865 98.985 183.185 99.245 ;
        RECT 183.875 99.230 184.015 99.725 ;
        RECT 185.165 99.665 185.485 99.925 ;
        RECT 188.475 99.910 188.615 100.405 ;
        RECT 199.440 100.405 200.665 100.545 ;
        RECT 199.440 100.360 199.730 100.405 ;
        RECT 200.345 100.345 200.665 100.405 ;
        RECT 205.405 100.545 205.725 100.605 ;
        RECT 216.000 100.545 216.290 100.590 ;
        RECT 216.445 100.545 216.765 100.605 ;
        RECT 205.405 100.405 210.695 100.545 ;
        RECT 205.405 100.345 205.725 100.405 ;
        RECT 192.060 100.205 192.710 100.250 ;
        RECT 194.825 100.205 195.145 100.265 ;
        RECT 195.660 100.205 195.950 100.250 ;
        RECT 192.060 100.065 195.950 100.205 ;
        RECT 192.060 100.020 192.710 100.065 ;
        RECT 194.825 100.005 195.145 100.065 ;
        RECT 195.360 100.020 195.950 100.065 ;
        RECT 203.220 100.205 203.510 100.250 ;
        RECT 206.460 100.205 207.110 100.250 ;
        RECT 209.085 100.205 209.405 100.265 ;
        RECT 203.220 100.065 209.405 100.205 ;
        RECT 203.220 100.020 203.810 100.065 ;
        RECT 206.460 100.020 207.110 100.065 ;
        RECT 188.400 99.680 188.690 99.910 ;
        RECT 188.865 99.865 189.155 99.910 ;
        RECT 190.700 99.865 190.990 99.910 ;
        RECT 194.280 99.865 194.570 99.910 ;
        RECT 188.865 99.725 194.570 99.865 ;
        RECT 188.865 99.680 189.155 99.725 ;
        RECT 190.700 99.680 190.990 99.725 ;
        RECT 194.280 99.680 194.570 99.725 ;
        RECT 195.360 99.705 195.650 100.020 ;
        RECT 198.965 99.865 199.285 99.925 ;
        RECT 196.755 99.725 199.285 99.865 ;
        RECT 186.085 99.325 186.405 99.585 ;
        RECT 186.560 99.340 186.850 99.570 ;
        RECT 183.800 99.000 184.090 99.230 ;
        RECT 186.635 98.845 186.775 99.340 ;
        RECT 189.765 99.325 190.085 99.585 ;
        RECT 190.225 99.525 190.545 99.585 ;
        RECT 196.755 99.525 196.895 99.725 ;
        RECT 198.965 99.665 199.285 99.725 ;
        RECT 203.520 99.705 203.810 100.020 ;
        RECT 209.085 100.005 209.405 100.065 ;
        RECT 210.555 99.910 210.695 100.405 ;
        RECT 216.000 100.405 216.765 100.545 ;
        RECT 216.000 100.360 216.290 100.405 ;
        RECT 216.445 100.345 216.765 100.405 ;
        RECT 217.840 100.545 218.130 100.590 ;
        RECT 218.745 100.545 219.065 100.605 ;
        RECT 217.840 100.405 219.065 100.545 ;
        RECT 217.840 100.360 218.130 100.405 ;
        RECT 218.745 100.345 219.065 100.405 ;
        RECT 219.665 100.545 219.985 100.605 ;
        RECT 223.820 100.545 224.110 100.590 ;
        RECT 224.725 100.545 225.045 100.605 ;
        RECT 226.105 100.545 226.425 100.605 ;
        RECT 219.665 100.405 223.575 100.545 ;
        RECT 219.665 100.345 219.985 100.405 ;
        RECT 220.140 100.205 220.430 100.250 ;
        RECT 223.435 100.205 223.575 100.405 ;
        RECT 223.820 100.405 226.425 100.545 ;
        RECT 223.820 100.360 224.110 100.405 ;
        RECT 224.725 100.345 225.045 100.405 ;
        RECT 226.105 100.345 226.425 100.405 ;
        RECT 228.405 100.345 228.725 100.605 ;
        RECT 229.800 100.360 230.090 100.590 ;
        RECT 236.685 100.545 237.005 100.605 ;
        RECT 236.685 100.405 238.295 100.545 ;
        RECT 227.025 100.205 227.345 100.265 ;
        RECT 211.475 100.065 221.505 100.205 ;
        RECT 223.435 100.065 227.345 100.205 ;
        RECT 211.475 99.925 211.615 100.065 ;
        RECT 220.140 100.020 220.430 100.065 ;
        RECT 204.600 99.865 204.890 99.910 ;
        RECT 208.180 99.865 208.470 99.910 ;
        RECT 210.015 99.865 210.305 99.910 ;
        RECT 204.600 99.725 210.305 99.865 ;
        RECT 204.600 99.680 204.890 99.725 ;
        RECT 208.180 99.680 208.470 99.725 ;
        RECT 210.015 99.680 210.305 99.725 ;
        RECT 210.480 99.680 210.770 99.910 ;
        RECT 211.385 99.665 211.705 99.925 ;
        RECT 211.845 99.665 212.165 99.925 ;
        RECT 215.065 99.665 215.385 99.925 ;
        RECT 216.920 99.865 217.210 99.910 ;
        RECT 215.615 99.725 217.210 99.865 ;
        RECT 221.365 99.865 221.505 100.065 ;
        RECT 227.025 100.005 227.345 100.065 ;
        RECT 223.345 99.865 223.665 99.925 ;
        RECT 227.945 99.865 228.265 99.925 ;
        RECT 221.365 99.725 223.665 99.865 ;
        RECT 190.225 99.385 196.895 99.525 ;
        RECT 198.520 99.525 198.810 99.570 ;
        RECT 209.100 99.525 209.390 99.570 ;
        RECT 198.520 99.385 199.195 99.525 ;
        RECT 190.225 99.325 190.545 99.385 ;
        RECT 198.520 99.340 198.810 99.385 ;
        RECT 189.270 99.185 189.560 99.230 ;
        RECT 191.160 99.185 191.450 99.230 ;
        RECT 194.280 99.185 194.570 99.230 ;
        RECT 189.270 99.045 194.570 99.185 ;
        RECT 189.270 99.000 189.560 99.045 ;
        RECT 191.160 99.000 191.450 99.045 ;
        RECT 194.280 99.000 194.570 99.045 ;
        RECT 199.055 98.905 199.195 99.385 ;
        RECT 209.100 99.385 211.155 99.525 ;
        RECT 209.100 99.340 209.390 99.385 ;
        RECT 211.015 99.230 211.155 99.385 ;
        RECT 204.600 99.185 204.890 99.230 ;
        RECT 207.720 99.185 208.010 99.230 ;
        RECT 209.610 99.185 209.900 99.230 ;
        RECT 204.600 99.045 209.900 99.185 ;
        RECT 204.600 99.000 204.890 99.045 ;
        RECT 207.720 99.000 208.010 99.045 ;
        RECT 209.610 99.000 209.900 99.045 ;
        RECT 210.940 99.000 211.230 99.230 ;
        RECT 215.615 99.185 215.755 99.725 ;
        RECT 216.920 99.680 217.210 99.725 ;
        RECT 223.345 99.665 223.665 99.725 ;
        RECT 223.895 99.725 228.265 99.865 ;
        RECT 216.445 99.525 216.765 99.585 ;
        RECT 223.895 99.525 224.035 99.725 ;
        RECT 227.945 99.665 228.265 99.725 ;
        RECT 229.340 99.865 229.630 99.910 ;
        RECT 229.875 99.865 230.015 100.360 ;
        RECT 236.685 100.345 237.005 100.405 ;
        RECT 232.100 100.205 232.390 100.250 ;
        RECT 238.155 100.205 238.295 100.405 ;
        RECT 239.905 100.345 240.225 100.605 ;
        RECT 243.600 100.545 243.890 100.590 ;
        RECT 244.045 100.545 244.365 100.605 ;
        RECT 243.600 100.405 244.365 100.545 ;
        RECT 243.600 100.360 243.890 100.405 ;
        RECT 244.045 100.345 244.365 100.405 ;
        RECT 249.105 100.545 249.425 100.605 ;
        RECT 253.705 100.545 254.025 100.605 ;
        RECT 249.105 100.405 255.315 100.545 ;
        RECT 249.105 100.345 249.425 100.405 ;
        RECT 253.705 100.345 254.025 100.405 ;
        RECT 248.645 100.250 248.965 100.265 ;
        RECT 245.080 100.205 245.370 100.250 ;
        RECT 248.320 100.205 248.970 100.250 ;
        RECT 232.100 100.065 237.835 100.205 ;
        RECT 238.155 100.065 241.975 100.205 ;
        RECT 232.100 100.020 232.390 100.065 ;
        RECT 237.695 99.925 237.835 100.065 ;
        RECT 241.835 99.925 241.975 100.065 ;
        RECT 245.080 100.065 248.970 100.205 ;
        RECT 245.080 100.020 245.670 100.065 ;
        RECT 248.320 100.020 248.970 100.065 ;
        RECT 250.485 100.205 250.805 100.265 ;
        RECT 250.960 100.205 251.250 100.250 ;
        RECT 250.485 100.065 251.250 100.205 ;
        RECT 229.340 99.725 230.015 99.865 ;
        RECT 229.340 99.680 229.630 99.725 ;
        RECT 231.625 99.665 231.945 99.925 ;
        RECT 237.605 99.665 237.925 99.925 ;
        RECT 240.365 99.865 240.685 99.925 ;
        RECT 240.840 99.865 241.130 99.910 ;
        RECT 240.365 99.725 241.130 99.865 ;
        RECT 240.365 99.665 240.685 99.725 ;
        RECT 240.840 99.680 241.130 99.725 ;
        RECT 241.745 99.665 242.065 99.925 ;
        RECT 245.380 99.705 245.670 100.020 ;
        RECT 248.645 100.005 248.965 100.020 ;
        RECT 250.485 100.005 250.805 100.065 ;
        RECT 250.960 100.020 251.250 100.065 ;
        RECT 254.625 100.005 254.945 100.265 ;
        RECT 255.175 100.250 255.315 100.405 ;
        RECT 256.480 100.360 256.770 100.590 ;
        RECT 259.685 100.545 260.005 100.605 ;
        RECT 257.015 100.405 260.005 100.545 ;
        RECT 255.100 100.020 255.390 100.250 ;
        RECT 246.460 99.865 246.750 99.910 ;
        RECT 250.040 99.865 250.330 99.910 ;
        RECT 251.875 99.865 252.165 99.910 ;
        RECT 246.460 99.725 252.165 99.865 ;
        RECT 246.460 99.680 246.750 99.725 ;
        RECT 250.040 99.680 250.330 99.725 ;
        RECT 251.875 99.680 252.165 99.725 ;
        RECT 252.325 99.665 252.645 99.925 ;
        RECT 252.785 99.865 253.105 99.925 ;
        RECT 253.720 99.865 254.010 99.910 ;
        RECT 254.165 99.865 254.485 99.925 ;
        RECT 252.785 99.725 254.485 99.865 ;
        RECT 252.785 99.665 253.105 99.725 ;
        RECT 253.720 99.680 254.010 99.725 ;
        RECT 254.165 99.665 254.485 99.725 ;
        RECT 216.445 99.385 224.035 99.525 ;
        RECT 224.740 99.525 225.030 99.570 ;
        RECT 225.645 99.525 225.965 99.585 ;
        RECT 232.545 99.525 232.865 99.585 ;
        RECT 224.740 99.385 232.865 99.525 ;
        RECT 216.445 99.325 216.765 99.385 ;
        RECT 224.740 99.340 225.030 99.385 ;
        RECT 225.645 99.325 225.965 99.385 ;
        RECT 232.545 99.325 232.865 99.385 ;
        RECT 235.765 99.525 236.085 99.585 ;
        RECT 254.715 99.525 254.855 100.005 ;
        RECT 255.545 99.665 255.865 99.925 ;
        RECT 256.555 99.865 256.695 100.360 ;
        RECT 257.015 100.265 257.155 100.405 ;
        RECT 259.685 100.345 260.005 100.405 ;
        RECT 287.745 100.545 288.065 100.605 ;
        RECT 287.745 100.405 295.335 100.545 ;
        RECT 287.745 100.345 288.065 100.405 ;
        RECT 256.925 100.005 257.245 100.265 ;
        RECT 262.905 100.205 263.225 100.265 ;
        RECT 274.865 100.250 275.185 100.265 ;
        RECT 259.595 100.065 263.225 100.205 ;
        RECT 259.595 99.910 259.735 100.065 ;
        RECT 262.905 100.005 263.225 100.065 ;
        RECT 274.860 100.205 275.510 100.250 ;
        RECT 278.460 100.205 278.750 100.250 ;
        RECT 274.860 100.065 278.750 100.205 ;
        RECT 274.860 100.020 275.510 100.065 ;
        RECT 278.160 100.020 278.750 100.065 ;
        RECT 274.865 100.005 275.185 100.020 ;
        RECT 258.780 99.865 259.070 99.910 ;
        RECT 256.555 99.725 259.070 99.865 ;
        RECT 258.780 99.680 259.070 99.725 ;
        RECT 259.520 99.680 259.810 99.910 ;
        RECT 260.145 99.665 260.465 99.925 ;
        RECT 261.065 99.910 261.385 99.925 ;
        RECT 260.620 99.680 260.910 99.910 ;
        RECT 261.065 99.865 261.600 99.910 ;
        RECT 262.445 99.865 262.765 99.925 ;
        RECT 261.065 99.725 262.765 99.865 ;
        RECT 261.065 99.680 261.600 99.725 ;
        RECT 260.695 99.525 260.835 99.680 ;
        RECT 261.065 99.665 261.385 99.680 ;
        RECT 262.445 99.665 262.765 99.725 ;
        RECT 263.840 99.865 264.130 99.910 ;
        RECT 264.285 99.865 264.605 99.925 ;
        RECT 271.665 99.865 271.955 99.910 ;
        RECT 273.500 99.865 273.790 99.910 ;
        RECT 277.080 99.865 277.370 99.910 ;
        RECT 263.840 99.725 268.655 99.865 ;
        RECT 263.840 99.680 264.130 99.725 ;
        RECT 264.285 99.665 264.605 99.725 ;
        RECT 268.515 99.585 268.655 99.725 ;
        RECT 271.665 99.725 277.370 99.865 ;
        RECT 271.665 99.680 271.955 99.725 ;
        RECT 273.500 99.680 273.790 99.725 ;
        RECT 277.080 99.680 277.370 99.725 ;
        RECT 278.160 99.705 278.450 100.020 ;
        RECT 283.145 100.005 283.465 100.265 ;
        RECT 285.440 100.205 286.090 100.250 ;
        RECT 289.040 100.205 289.330 100.250 ;
        RECT 290.135 100.205 290.275 100.405 ;
        RECT 295.195 100.265 295.335 100.405 ;
        RECT 303.845 100.345 304.165 100.605 ;
        RECT 307.080 100.545 307.370 100.590 ;
        RECT 308.905 100.545 309.225 100.605 ;
        RECT 307.080 100.405 309.225 100.545 ;
        RECT 307.080 100.360 307.370 100.405 ;
        RECT 308.905 100.345 309.225 100.405 ;
        RECT 285.440 100.065 290.275 100.205 ;
        RECT 290.505 100.205 290.825 100.265 ;
        RECT 293.740 100.205 294.030 100.250 ;
        RECT 290.505 100.065 294.030 100.205 ;
        RECT 285.440 100.020 286.090 100.065 ;
        RECT 288.740 100.020 289.330 100.065 ;
        RECT 280.385 99.665 280.705 99.925 ;
        RECT 282.245 99.865 282.535 99.910 ;
        RECT 284.080 99.865 284.370 99.910 ;
        RECT 287.660 99.865 287.950 99.910 ;
        RECT 282.245 99.725 287.950 99.865 ;
        RECT 282.245 99.680 282.535 99.725 ;
        RECT 284.080 99.680 284.370 99.725 ;
        RECT 287.660 99.680 287.950 99.725 ;
        RECT 288.740 99.705 289.030 100.020 ;
        RECT 290.505 100.005 290.825 100.065 ;
        RECT 293.740 100.020 294.030 100.065 ;
        RECT 295.105 100.205 295.425 100.265 ;
        RECT 296.020 100.205 296.670 100.250 ;
        RECT 299.620 100.205 299.910 100.250 ;
        RECT 295.105 100.065 299.910 100.205 ;
        RECT 295.105 100.005 295.425 100.065 ;
        RECT 296.020 100.020 296.670 100.065 ;
        RECT 299.320 100.020 299.910 100.065 ;
        RECT 292.825 99.865 293.115 99.910 ;
        RECT 294.660 99.865 294.950 99.910 ;
        RECT 298.240 99.865 298.530 99.910 ;
        RECT 292.825 99.725 298.530 99.865 ;
        RECT 292.825 99.680 293.115 99.725 ;
        RECT 294.660 99.680 294.950 99.725 ;
        RECT 298.240 99.680 298.530 99.725 ;
        RECT 299.320 99.705 299.610 100.020 ;
        RECT 305.225 99.865 305.545 99.925 ;
        RECT 306.160 99.865 306.450 99.910 ;
        RECT 303.935 99.725 304.995 99.865 ;
        RECT 262.920 99.525 263.210 99.570 ;
        RECT 266.585 99.525 266.905 99.585 ;
        RECT 235.765 99.385 254.855 99.525 ;
        RECT 259.445 99.385 260.495 99.525 ;
        RECT 260.695 99.385 266.905 99.525 ;
        RECT 235.765 99.325 236.085 99.385 ;
        RECT 234.845 99.185 235.165 99.245 ;
        RECT 215.615 99.045 235.165 99.185 ;
        RECT 193.445 98.845 193.765 98.905 ;
        RECT 178.725 98.705 193.765 98.845 ;
        RECT 178.725 98.645 179.045 98.705 ;
        RECT 193.445 98.645 193.765 98.705 ;
        RECT 197.140 98.845 197.430 98.890 ;
        RECT 197.585 98.845 197.905 98.905 ;
        RECT 197.140 98.705 197.905 98.845 ;
        RECT 197.140 98.660 197.430 98.705 ;
        RECT 197.585 98.645 197.905 98.705 ;
        RECT 198.965 98.645 199.285 98.905 ;
        RECT 201.265 98.645 201.585 98.905 ;
        RECT 201.740 98.845 202.030 98.890 ;
        RECT 206.325 98.845 206.645 98.905 ;
        RECT 215.615 98.845 215.755 99.045 ;
        RECT 234.845 98.985 235.165 99.045 ;
        RECT 235.305 99.185 235.625 99.245 ;
        RECT 246.460 99.185 246.750 99.230 ;
        RECT 249.580 99.185 249.870 99.230 ;
        RECT 251.470 99.185 251.760 99.230 ;
        RECT 235.305 99.045 246.115 99.185 ;
        RECT 235.305 98.985 235.625 99.045 ;
        RECT 201.740 98.705 215.755 98.845 ;
        RECT 215.985 98.845 216.305 98.905 ;
        RECT 221.520 98.845 221.810 98.890 ;
        RECT 215.985 98.705 221.810 98.845 ;
        RECT 201.740 98.660 202.030 98.705 ;
        RECT 206.325 98.645 206.645 98.705 ;
        RECT 215.985 98.645 216.305 98.705 ;
        RECT 221.520 98.660 221.810 98.705 ;
        RECT 231.625 98.845 231.945 98.905 ;
        RECT 244.505 98.845 244.825 98.905 ;
        RECT 231.625 98.705 244.825 98.845 ;
        RECT 245.975 98.845 246.115 99.045 ;
        RECT 246.460 99.045 251.760 99.185 ;
        RECT 246.460 99.000 246.750 99.045 ;
        RECT 249.580 99.000 249.870 99.045 ;
        RECT 251.470 99.000 251.760 99.045 ;
        RECT 252.325 99.185 252.645 99.245 ;
        RECT 259.445 99.185 259.585 99.385 ;
        RECT 252.325 99.045 259.585 99.185 ;
        RECT 260.355 99.185 260.495 99.385 ;
        RECT 262.920 99.340 263.210 99.385 ;
        RECT 266.585 99.325 266.905 99.385 ;
        RECT 268.425 99.325 268.745 99.585 ;
        RECT 271.200 99.340 271.490 99.570 ;
        RECT 270.725 99.185 271.045 99.245 ;
        RECT 271.275 99.185 271.415 99.340 ;
        RECT 272.565 99.325 272.885 99.585 ;
        RECT 281.780 99.525 282.070 99.570 ;
        RECT 292.360 99.525 292.650 99.570 ;
        RECT 277.715 99.385 292.650 99.525 ;
        RECT 260.355 99.045 271.415 99.185 ;
        RECT 252.325 98.985 252.645 99.045 ;
        RECT 270.725 98.985 271.045 99.045 ;
        RECT 257.845 98.845 258.165 98.905 ;
        RECT 245.975 98.705 258.165 98.845 ;
        RECT 231.625 98.645 231.945 98.705 ;
        RECT 244.505 98.645 244.825 98.705 ;
        RECT 257.845 98.645 258.165 98.705 ;
        RECT 261.065 98.845 261.385 98.905 ;
        RECT 262.000 98.845 262.290 98.890 ;
        RECT 261.065 98.705 262.290 98.845 ;
        RECT 261.065 98.645 261.385 98.705 ;
        RECT 262.000 98.660 262.290 98.705 ;
        RECT 264.760 98.845 265.050 98.890 ;
        RECT 265.665 98.845 265.985 98.905 ;
        RECT 264.760 98.705 265.985 98.845 ;
        RECT 271.275 98.845 271.415 99.045 ;
        RECT 272.070 99.185 272.360 99.230 ;
        RECT 273.960 99.185 274.250 99.230 ;
        RECT 277.080 99.185 277.370 99.230 ;
        RECT 272.070 99.045 277.370 99.185 ;
        RECT 272.070 99.000 272.360 99.045 ;
        RECT 273.960 99.000 274.250 99.045 ;
        RECT 277.080 99.000 277.370 99.045 ;
        RECT 277.715 98.905 277.855 99.385 ;
        RECT 281.780 99.340 282.070 99.385 ;
        RECT 292.360 99.340 292.650 99.385 ;
        RECT 296.945 99.525 297.265 99.585 ;
        RECT 303.935 99.525 304.075 99.725 ;
        RECT 304.855 99.570 304.995 99.725 ;
        RECT 305.225 99.725 306.450 99.865 ;
        RECT 305.225 99.665 305.545 99.725 ;
        RECT 306.160 99.680 306.450 99.725 ;
        RECT 308.000 99.680 308.290 99.910 ;
        RECT 296.945 99.385 304.075 99.525 ;
        RECT 296.945 99.325 297.265 99.385 ;
        RECT 304.320 99.340 304.610 99.570 ;
        RECT 304.780 99.340 305.070 99.570 ;
        RECT 305.685 99.525 306.005 99.585 ;
        RECT 308.075 99.525 308.215 99.680 ;
        RECT 305.685 99.385 308.215 99.525 ;
        RECT 282.650 99.185 282.940 99.230 ;
        RECT 284.540 99.185 284.830 99.230 ;
        RECT 287.660 99.185 287.950 99.230 ;
        RECT 282.650 99.045 287.950 99.185 ;
        RECT 282.650 99.000 282.940 99.045 ;
        RECT 284.540 99.000 284.830 99.045 ;
        RECT 287.660 99.000 287.950 99.045 ;
        RECT 293.230 99.185 293.520 99.230 ;
        RECT 295.120 99.185 295.410 99.230 ;
        RECT 298.240 99.185 298.530 99.230 ;
        RECT 293.230 99.045 298.530 99.185 ;
        RECT 293.230 99.000 293.520 99.045 ;
        RECT 295.120 99.000 295.410 99.045 ;
        RECT 298.240 99.000 298.530 99.045 ;
        RECT 299.245 99.185 299.565 99.245 ;
        RECT 304.395 99.185 304.535 99.340 ;
        RECT 305.685 99.325 306.005 99.385 ;
        RECT 299.245 99.045 304.535 99.185 ;
        RECT 299.245 98.985 299.565 99.045 ;
        RECT 277.625 98.845 277.945 98.905 ;
        RECT 271.275 98.705 277.945 98.845 ;
        RECT 264.760 98.660 265.050 98.705 ;
        RECT 265.665 98.645 265.985 98.705 ;
        RECT 277.625 98.645 277.945 98.705 ;
        RECT 279.925 98.645 280.245 98.905 ;
        RECT 281.320 98.845 281.610 98.890 ;
        RECT 286.365 98.845 286.685 98.905 ;
        RECT 281.320 98.705 286.685 98.845 ;
        RECT 281.320 98.660 281.610 98.705 ;
        RECT 286.365 98.645 286.685 98.705 ;
        RECT 288.205 98.845 288.525 98.905 ;
        RECT 290.520 98.845 290.810 98.890 ;
        RECT 288.205 98.705 290.810 98.845 ;
        RECT 288.205 98.645 288.525 98.705 ;
        RECT 290.520 98.660 290.810 98.705 ;
        RECT 293.725 98.845 294.045 98.905 ;
        RECT 301.100 98.845 301.390 98.890 ;
        RECT 293.725 98.705 301.390 98.845 ;
        RECT 293.725 98.645 294.045 98.705 ;
        RECT 301.100 98.660 301.390 98.705 ;
        RECT 302.005 98.645 302.325 98.905 ;
        RECT 304.305 98.845 304.625 98.905 ;
        RECT 308.920 98.845 309.210 98.890 ;
        RECT 304.305 98.705 309.210 98.845 ;
        RECT 304.305 98.645 304.625 98.705 ;
        RECT 308.920 98.660 309.210 98.705 ;
        RECT 162.095 98.025 311.135 98.505 ;
        RECT 169.985 97.825 170.305 97.885 ;
        RECT 171.380 97.825 171.670 97.870 ;
        RECT 177.805 97.825 178.125 97.885 ;
        RECT 169.985 97.685 171.670 97.825 ;
        RECT 169.985 97.625 170.305 97.685 ;
        RECT 171.380 97.640 171.670 97.685 ;
        RECT 173.065 97.685 178.125 97.825 ;
        RECT 170.920 96.620 171.210 96.850 ;
        RECT 172.300 96.805 172.590 96.850 ;
        RECT 173.065 96.805 173.205 97.685 ;
        RECT 177.805 97.625 178.125 97.685 ;
        RECT 189.765 97.825 190.085 97.885 ;
        RECT 193.000 97.825 193.290 97.870 ;
        RECT 189.765 97.685 193.290 97.825 ;
        RECT 189.765 97.625 190.085 97.685 ;
        RECT 193.000 97.640 193.290 97.685 ;
        RECT 193.445 97.825 193.765 97.885 ;
        RECT 201.280 97.825 201.570 97.870 ;
        RECT 193.445 97.685 201.570 97.825 ;
        RECT 193.445 97.625 193.765 97.685 ;
        RECT 201.280 97.640 201.570 97.685 ;
        RECT 202.185 97.825 202.505 97.885 ;
        RECT 207.705 97.825 208.025 97.885 ;
        RECT 202.185 97.685 208.025 97.825 ;
        RECT 202.185 97.625 202.505 97.685 ;
        RECT 207.705 97.625 208.025 97.685 ;
        RECT 208.180 97.825 208.470 97.870 ;
        RECT 211.845 97.825 212.165 97.885 ;
        RECT 208.180 97.685 212.165 97.825 ;
        RECT 208.180 97.640 208.470 97.685 ;
        RECT 211.845 97.625 212.165 97.685 ;
        RECT 216.920 97.825 217.210 97.870 ;
        RECT 219.205 97.825 219.525 97.885 ;
        RECT 216.920 97.685 219.525 97.825 ;
        RECT 216.920 97.640 217.210 97.685 ;
        RECT 219.205 97.625 219.525 97.685 ;
        RECT 219.665 97.625 219.985 97.885 ;
        RECT 225.185 97.825 225.505 97.885 ;
        RECT 239.445 97.825 239.765 97.885 ;
        RECT 225.185 97.685 239.765 97.825 ;
        RECT 225.185 97.625 225.505 97.685 ;
        RECT 239.445 97.625 239.765 97.685 ;
        RECT 264.745 97.625 265.065 97.885 ;
        RECT 265.665 97.625 265.985 97.885 ;
        RECT 272.565 97.825 272.885 97.885 ;
        RECT 273.500 97.825 273.790 97.870 ;
        RECT 272.565 97.685 273.790 97.825 ;
        RECT 272.565 97.625 272.885 97.685 ;
        RECT 273.500 97.640 273.790 97.685 ;
        RECT 280.385 97.825 280.705 97.885 ;
        RECT 286.840 97.825 287.130 97.870 ;
        RECT 280.385 97.685 287.130 97.825 ;
        RECT 280.385 97.625 280.705 97.685 ;
        RECT 286.840 97.640 287.130 97.685 ;
        RECT 289.585 97.825 289.905 97.885 ;
        RECT 292.345 97.825 292.665 97.885 ;
        RECT 289.585 97.685 292.665 97.825 ;
        RECT 289.585 97.625 289.905 97.685 ;
        RECT 292.345 97.625 292.665 97.685 ;
        RECT 301.545 97.625 301.865 97.885 ;
        RECT 306.605 97.825 306.925 97.885 ;
        RECT 308.920 97.825 309.210 97.870 ;
        RECT 306.605 97.685 309.210 97.825 ;
        RECT 306.605 97.625 306.925 97.685 ;
        RECT 308.920 97.640 309.210 97.685 ;
        RECT 184.210 97.485 184.500 97.530 ;
        RECT 186.100 97.485 186.390 97.530 ;
        RECT 189.220 97.485 189.510 97.530 ;
        RECT 184.210 97.345 189.510 97.485 ;
        RECT 184.210 97.300 184.500 97.345 ;
        RECT 186.100 97.300 186.390 97.345 ;
        RECT 189.220 97.300 189.510 97.345 ;
        RECT 192.065 97.485 192.385 97.545 ;
        RECT 203.565 97.485 203.885 97.545 ;
        RECT 208.640 97.485 208.930 97.530 ;
        RECT 209.545 97.485 209.865 97.545 ;
        RECT 218.285 97.485 218.605 97.545 ;
        RECT 192.065 97.345 203.885 97.485 ;
        RECT 192.065 97.285 192.385 97.345 ;
        RECT 203.565 97.285 203.885 97.345 ;
        RECT 205.495 97.345 209.865 97.485 ;
        RECT 178.725 96.945 179.045 97.205 ;
        RECT 185.165 97.145 185.485 97.205 ;
        RECT 185.165 97.005 194.595 97.145 ;
        RECT 185.165 96.945 185.485 97.005 ;
        RECT 172.300 96.665 173.205 96.805 ;
        RECT 173.680 96.805 173.970 96.850 ;
        RECT 173.680 96.665 175.735 96.805 ;
        RECT 172.300 96.620 172.590 96.665 ;
        RECT 173.680 96.620 173.970 96.665 ;
        RECT 170.995 96.465 171.135 96.620 ;
        RECT 174.125 96.465 174.445 96.525 ;
        RECT 170.995 96.325 174.445 96.465 ;
        RECT 174.125 96.265 174.445 96.325 ;
        RECT 169.985 95.925 170.305 96.185 ;
        RECT 171.365 96.125 171.685 96.185 ;
        RECT 175.595 96.170 175.735 96.665 ;
        RECT 177.345 96.605 177.665 96.865 ;
        RECT 183.325 96.605 183.645 96.865 ;
        RECT 183.805 96.805 184.095 96.850 ;
        RECT 185.640 96.805 185.930 96.850 ;
        RECT 189.220 96.805 189.510 96.850 ;
        RECT 183.805 96.665 189.510 96.805 ;
        RECT 183.805 96.620 184.095 96.665 ;
        RECT 185.640 96.620 185.930 96.665 ;
        RECT 189.220 96.620 189.510 96.665 ;
        RECT 183.415 96.465 183.555 96.605 ;
        RECT 183.415 96.325 184.475 96.465 ;
        RECT 184.335 96.185 184.475 96.325 ;
        RECT 184.705 96.265 185.025 96.525 ;
        RECT 190.300 96.510 190.590 96.825 ;
        RECT 193.920 96.620 194.210 96.850 ;
        RECT 194.455 96.805 194.595 97.005 ;
        RECT 198.045 96.945 198.365 97.205 ;
        RECT 198.965 97.145 199.285 97.205 ;
        RECT 205.495 97.190 205.635 97.345 ;
        RECT 208.640 97.300 208.930 97.345 ;
        RECT 209.545 97.285 209.865 97.345 ;
        RECT 215.155 97.345 218.605 97.485 ;
        RECT 205.420 97.145 205.710 97.190 ;
        RECT 210.005 97.145 210.325 97.205 ;
        RECT 215.155 97.145 215.295 97.345 ;
        RECT 218.285 97.285 218.605 97.345 ;
        RECT 216.445 97.145 216.765 97.205 ;
        RECT 219.755 97.145 219.895 97.625 ;
        RECT 221.045 97.285 221.365 97.545 ;
        RECT 222.055 97.345 235.995 97.485 ;
        RECT 198.965 97.005 205.710 97.145 ;
        RECT 198.965 96.945 199.285 97.005 ;
        RECT 205.420 96.960 205.710 97.005 ;
        RECT 207.340 97.005 215.295 97.145 ;
        RECT 215.615 97.005 216.765 97.145 ;
        RECT 201.725 96.805 202.045 96.865 ;
        RECT 194.455 96.665 202.045 96.805 ;
        RECT 187.000 96.465 187.650 96.510 ;
        RECT 190.300 96.465 190.890 96.510 ;
        RECT 191.605 96.465 191.925 96.525 ;
        RECT 187.000 96.325 191.925 96.465 ;
        RECT 193.995 96.465 194.135 96.620 ;
        RECT 201.725 96.605 202.045 96.665 ;
        RECT 202.185 96.605 202.505 96.865 ;
        RECT 203.105 96.605 203.425 96.865 ;
        RECT 203.580 96.805 203.870 96.850 ;
        RECT 207.340 96.805 207.480 97.005 ;
        RECT 210.005 96.945 210.325 97.005 ;
        RECT 203.580 96.665 207.480 96.805 ;
        RECT 207.705 96.805 208.025 96.865 ;
        RECT 209.560 96.805 209.850 96.850 ;
        RECT 207.705 96.665 209.850 96.805 ;
        RECT 203.580 96.620 203.870 96.665 ;
        RECT 207.705 96.605 208.025 96.665 ;
        RECT 209.560 96.620 209.850 96.665 ;
        RECT 210.480 96.620 210.770 96.850 ;
        RECT 210.940 96.805 211.230 96.850 ;
        RECT 215.615 96.805 215.755 97.005 ;
        RECT 216.445 96.945 216.765 97.005 ;
        RECT 218.375 97.005 219.895 97.145 ;
        RECT 210.940 96.665 215.755 96.805 ;
        RECT 210.940 96.620 211.230 96.665 ;
        RECT 197.585 96.465 197.905 96.525 ;
        RECT 205.405 96.465 205.725 96.525 ;
        RECT 193.995 96.325 195.975 96.465 ;
        RECT 187.000 96.280 187.650 96.325 ;
        RECT 190.600 96.280 190.890 96.325 ;
        RECT 191.605 96.265 191.925 96.325 ;
        RECT 172.760 96.125 173.050 96.170 ;
        RECT 171.365 95.985 173.050 96.125 ;
        RECT 171.365 95.925 171.685 95.985 ;
        RECT 172.760 95.940 173.050 95.985 ;
        RECT 175.520 95.940 175.810 96.170 ;
        RECT 177.805 95.925 178.125 96.185 ;
        RECT 184.245 95.925 184.565 96.185 ;
        RECT 195.835 96.170 195.975 96.325 ;
        RECT 197.585 96.325 205.725 96.465 ;
        RECT 197.585 96.265 197.905 96.325 ;
        RECT 205.405 96.265 205.725 96.325 ;
        RECT 206.325 96.265 206.645 96.525 ;
        RECT 210.555 96.465 210.695 96.620 ;
        RECT 215.985 96.605 216.305 96.865 ;
        RECT 218.375 96.850 218.515 97.005 ;
        RECT 218.300 96.620 218.590 96.850 ;
        RECT 219.665 96.605 219.985 96.865 ;
        RECT 220.125 96.605 220.445 96.865 ;
        RECT 222.055 96.805 222.195 97.345 ;
        RECT 229.325 97.145 229.645 97.205 ;
        RECT 234.385 97.145 234.705 97.205 ;
        RECT 223.435 97.005 234.705 97.145 ;
        RECT 220.675 96.665 222.195 96.805 ;
        RECT 208.715 96.325 210.695 96.465 ;
        RECT 219.220 96.465 219.510 96.510 ;
        RECT 220.675 96.465 220.815 96.665 ;
        RECT 222.425 96.605 222.745 96.865 ;
        RECT 223.435 96.850 223.575 97.005 ;
        RECT 229.325 96.945 229.645 97.005 ;
        RECT 234.385 96.945 234.705 97.005 ;
        RECT 235.855 96.865 235.995 97.345 ;
        RECT 236.685 97.285 237.005 97.545 ;
        RECT 237.620 97.300 237.910 97.530 ;
        RECT 236.775 97.145 236.915 97.285 ;
        RECT 236.315 97.005 236.915 97.145 ;
        RECT 223.360 96.620 223.650 96.850 ;
        RECT 224.265 96.605 224.585 96.865 ;
        RECT 227.025 96.605 227.345 96.865 ;
        RECT 228.880 96.805 229.170 96.850 ;
        RECT 231.165 96.805 231.485 96.865 ;
        RECT 228.880 96.665 231.485 96.805 ;
        RECT 228.880 96.620 229.170 96.665 ;
        RECT 231.165 96.605 231.485 96.665 ;
        RECT 234.845 96.605 235.165 96.865 ;
        RECT 235.765 96.605 236.085 96.865 ;
        RECT 236.315 96.850 236.455 97.005 ;
        RECT 236.240 96.620 236.530 96.850 ;
        RECT 236.700 96.805 236.990 96.850 ;
        RECT 237.145 96.805 237.465 96.865 ;
        RECT 236.700 96.665 237.465 96.805 ;
        RECT 237.695 96.805 237.835 97.300 ;
        RECT 238.080 96.805 238.370 96.850 ;
        RECT 237.695 96.665 238.370 96.805 ;
        RECT 236.700 96.620 236.990 96.665 ;
        RECT 237.145 96.605 237.465 96.665 ;
        RECT 238.080 96.620 238.370 96.665 ;
        RECT 238.525 96.805 238.845 96.865 ;
        RECT 239.535 96.850 239.675 97.625 ;
        RECT 257.385 97.285 257.705 97.545 ;
        RECT 260.605 97.485 260.925 97.545 ;
        RECT 258.395 97.345 260.925 97.485 ;
        RECT 254.165 97.145 254.485 97.205 ;
        RECT 240.580 97.005 254.485 97.145 ;
        RECT 238.525 96.665 239.040 96.805 ;
        RECT 238.525 96.605 238.845 96.665 ;
        RECT 239.460 96.620 239.750 96.850 ;
        RECT 239.905 96.605 240.225 96.865 ;
        RECT 240.580 96.850 240.720 97.005 ;
        RECT 254.165 96.945 254.485 97.005 ;
        RECT 255.175 97.005 257.615 97.145 ;
        RECT 240.500 96.805 240.790 96.850 ;
        RECT 247.265 96.805 247.585 96.865 ;
        RECT 240.460 96.620 240.790 96.805 ;
        RECT 241.045 96.665 247.585 96.805 ;
        RECT 222.900 96.465 223.190 96.510 ;
        RECT 219.220 96.325 220.815 96.465 ;
        RECT 221.135 96.325 223.190 96.465 ;
        RECT 208.715 96.185 208.855 96.325 ;
        RECT 219.220 96.280 219.510 96.325 ;
        RECT 195.760 95.940 196.050 96.170 ;
        RECT 200.345 96.125 200.665 96.185 ;
        RECT 205.880 96.125 206.170 96.170 ;
        RECT 208.165 96.125 208.485 96.185 ;
        RECT 200.345 95.985 208.485 96.125 ;
        RECT 200.345 95.925 200.665 95.985 ;
        RECT 205.880 95.940 206.170 95.985 ;
        RECT 208.165 95.925 208.485 95.985 ;
        RECT 208.625 95.925 208.945 96.185 ;
        RECT 215.985 96.125 216.305 96.185 ;
        RECT 219.295 96.125 219.435 96.280 ;
        RECT 215.985 95.985 219.435 96.125 ;
        RECT 219.665 96.125 219.985 96.185 ;
        RECT 221.135 96.125 221.275 96.325 ;
        RECT 222.900 96.280 223.190 96.325 ;
        RECT 227.945 96.265 228.265 96.525 ;
        RECT 228.405 96.465 228.725 96.525 ;
        RECT 234.385 96.465 234.705 96.525 ;
        RECT 240.460 96.465 240.600 96.620 ;
        RECT 241.045 96.465 241.185 96.665 ;
        RECT 247.265 96.605 247.585 96.665 ;
        RECT 253.705 96.805 254.025 96.865 ;
        RECT 254.640 96.805 254.930 96.850 ;
        RECT 253.705 96.665 254.930 96.805 ;
        RECT 253.705 96.605 254.025 96.665 ;
        RECT 254.640 96.620 254.930 96.665 ;
        RECT 228.405 96.325 232.315 96.465 ;
        RECT 228.405 96.265 228.725 96.325 ;
        RECT 219.665 95.985 221.275 96.125 ;
        RECT 215.985 95.925 216.305 95.985 ;
        RECT 219.665 95.925 219.985 95.985 ;
        RECT 221.505 95.925 221.825 96.185 ;
        RECT 222.425 96.125 222.745 96.185 ;
        RECT 225.185 96.125 225.505 96.185 ;
        RECT 222.425 95.985 225.505 96.125 ;
        RECT 222.425 95.925 222.745 95.985 ;
        RECT 225.185 95.925 225.505 95.985 ;
        RECT 229.785 95.925 230.105 96.185 ;
        RECT 232.175 96.125 232.315 96.325 ;
        RECT 234.385 96.325 240.600 96.465 ;
        RECT 240.915 96.325 241.185 96.465 ;
        RECT 242.205 96.465 242.525 96.525 ;
        RECT 255.175 96.465 255.315 97.005 ;
        RECT 255.545 96.605 255.865 96.865 ;
        RECT 256.465 96.605 256.785 96.865 ;
        RECT 242.205 96.325 255.315 96.465 ;
        RECT 234.385 96.265 234.705 96.325 ;
        RECT 240.915 96.125 241.055 96.325 ;
        RECT 242.205 96.265 242.525 96.325 ;
        RECT 256.005 96.265 256.325 96.525 ;
        RECT 257.475 96.465 257.615 97.005 ;
        RECT 257.845 96.685 258.165 96.945 ;
        RECT 258.395 96.850 258.535 97.345 ;
        RECT 260.605 97.285 260.925 97.345 ;
        RECT 264.300 97.485 264.590 97.530 ;
        RECT 264.300 97.345 265.435 97.485 ;
        RECT 264.300 97.300 264.590 97.345 ;
        RECT 265.295 97.190 265.435 97.345 ;
        RECT 259.315 97.005 263.595 97.145 ;
        RECT 257.860 96.620 258.150 96.685 ;
        RECT 258.325 96.620 258.615 96.850 ;
        RECT 259.315 96.510 259.455 97.005 ;
        RECT 259.685 96.605 260.005 96.865 ;
        RECT 260.145 96.850 260.465 96.865 ;
        RECT 260.145 96.805 260.475 96.850 ;
        RECT 260.145 96.665 260.660 96.805 ;
        RECT 260.145 96.620 260.475 96.665 ;
        RECT 260.145 96.605 260.465 96.620 ;
        RECT 261.525 96.605 261.845 96.865 ;
        RECT 263.455 96.850 263.595 97.005 ;
        RECT 265.220 96.960 265.510 97.190 ;
        RECT 263.380 96.620 263.670 96.850 ;
        RECT 263.825 96.805 264.145 96.865 ;
        RECT 264.760 96.805 265.050 96.850 ;
        RECT 263.825 96.665 265.050 96.805 ;
        RECT 265.755 96.805 265.895 97.625 ;
        RECT 267.045 97.485 267.365 97.545 ;
        RECT 267.045 97.345 285.675 97.485 ;
        RECT 267.045 97.285 267.365 97.345 ;
        RECT 266.585 97.145 266.905 97.205 ;
        RECT 279.465 97.145 279.785 97.205 ;
        RECT 281.320 97.145 281.610 97.190 ;
        RECT 282.225 97.145 282.545 97.205 ;
        RECT 283.605 97.145 283.925 97.205 ;
        RECT 266.585 97.005 279.235 97.145 ;
        RECT 266.585 96.945 266.905 97.005 ;
        RECT 266.140 96.805 266.430 96.850 ;
        RECT 265.755 96.665 266.430 96.805 ;
        RECT 263.825 96.605 264.145 96.665 ;
        RECT 264.760 96.620 265.050 96.665 ;
        RECT 266.140 96.620 266.430 96.665 ;
        RECT 268.885 96.605 269.205 96.865 ;
        RECT 274.420 96.805 274.710 96.850 ;
        RECT 274.420 96.665 278.775 96.805 ;
        RECT 274.420 96.620 274.710 96.665 ;
        RECT 259.240 96.465 259.530 96.510 ;
        RECT 257.475 96.325 259.530 96.465 ;
        RECT 259.240 96.280 259.530 96.325 ;
        RECT 260.605 96.465 260.925 96.525 ;
        RECT 262.905 96.510 263.225 96.525 ;
        RECT 262.460 96.465 262.750 96.510 ;
        RECT 260.605 96.325 262.750 96.465 ;
        RECT 260.605 96.265 260.925 96.325 ;
        RECT 262.460 96.280 262.750 96.325 ;
        RECT 262.900 96.465 263.225 96.510 ;
        RECT 268.975 96.465 269.115 96.605 ;
        RECT 262.900 96.325 269.115 96.465 ;
        RECT 262.900 96.280 263.225 96.325 ;
        RECT 262.905 96.265 263.225 96.280 ;
        RECT 232.175 95.985 241.055 96.125 ;
        RECT 241.285 95.925 241.605 96.185 ;
        RECT 261.065 95.925 261.385 96.185 ;
        RECT 265.205 96.125 265.525 96.185 ;
        RECT 278.635 96.170 278.775 96.665 ;
        RECT 279.095 96.465 279.235 97.005 ;
        RECT 279.465 97.005 283.925 97.145 ;
        RECT 279.465 96.945 279.785 97.005 ;
        RECT 281.320 96.960 281.610 97.005 ;
        RECT 282.225 96.945 282.545 97.005 ;
        RECT 283.605 96.945 283.925 97.005 ;
        RECT 284.065 97.145 284.385 97.205 ;
        RECT 285.000 97.145 285.290 97.190 ;
        RECT 284.065 97.005 285.290 97.145 ;
        RECT 284.065 96.945 284.385 97.005 ;
        RECT 285.000 96.960 285.290 97.005 ;
        RECT 279.925 96.805 280.245 96.865 ;
        RECT 280.400 96.805 280.690 96.850 ;
        RECT 279.925 96.665 280.690 96.805 ;
        RECT 279.925 96.605 280.245 96.665 ;
        RECT 280.400 96.620 280.690 96.665 ;
        RECT 280.845 96.605 281.165 96.865 ;
        RECT 281.855 96.665 283.835 96.805 ;
        RECT 281.855 96.465 281.995 96.665 ;
        RECT 283.695 96.525 283.835 96.665 ;
        RECT 284.540 96.685 284.830 96.850 ;
        RECT 285.535 96.805 285.675 97.345 ;
        RECT 300.180 97.300 300.470 97.530 ;
        RECT 285.905 97.145 286.225 97.205 ;
        RECT 289.600 97.145 289.890 97.190 ;
        RECT 285.905 97.005 289.890 97.145 ;
        RECT 285.905 96.945 286.225 97.005 ;
        RECT 289.600 96.960 289.890 97.005 ;
        RECT 292.805 97.145 293.125 97.205 ;
        RECT 294.660 97.145 294.950 97.190 ;
        RECT 296.945 97.145 297.265 97.205 ;
        RECT 292.805 97.005 297.265 97.145 ;
        RECT 292.805 96.945 293.125 97.005 ;
        RECT 294.660 96.960 294.950 97.005 ;
        RECT 296.945 96.945 297.265 97.005 ;
        RECT 297.865 96.945 298.185 97.205 ;
        RECT 300.255 97.145 300.395 97.300 ;
        RECT 300.255 97.005 303.155 97.145 ;
        RECT 288.205 96.805 288.525 96.865 ;
        RECT 285.535 96.685 288.525 96.805 ;
        RECT 284.540 96.665 288.525 96.685 ;
        RECT 284.540 96.620 285.675 96.665 ;
        RECT 284.615 96.545 285.675 96.620 ;
        RECT 288.205 96.605 288.525 96.665 ;
        RECT 288.680 96.805 288.970 96.850 ;
        RECT 290.045 96.805 290.365 96.865 ;
        RECT 288.680 96.665 290.365 96.805 ;
        RECT 288.680 96.620 288.970 96.665 ;
        RECT 290.045 96.605 290.365 96.665 ;
        RECT 293.725 96.605 294.045 96.865 ;
        RECT 300.640 96.805 300.930 96.850 ;
        RECT 302.005 96.805 302.325 96.865 ;
        RECT 303.015 96.850 303.155 97.005 ;
        RECT 300.640 96.665 302.325 96.805 ;
        RECT 300.640 96.620 300.930 96.665 ;
        RECT 302.005 96.605 302.325 96.665 ;
        RECT 302.940 96.620 303.230 96.850 ;
        RECT 307.985 96.605 308.305 96.865 ;
        RECT 279.095 96.325 281.995 96.465 ;
        RECT 282.315 96.325 283.375 96.465 ;
        RECT 267.060 96.125 267.350 96.170 ;
        RECT 265.205 95.985 267.350 96.125 ;
        RECT 265.205 95.925 265.525 95.985 ;
        RECT 267.060 95.940 267.350 95.985 ;
        RECT 278.560 95.940 278.850 96.170 ;
        RECT 279.465 96.125 279.785 96.185 ;
        RECT 282.315 96.125 282.455 96.325 ;
        RECT 279.465 95.985 282.455 96.125 ;
        RECT 279.465 95.925 279.785 95.985 ;
        RECT 282.685 95.925 283.005 96.185 ;
        RECT 283.235 96.125 283.375 96.325 ;
        RECT 283.605 96.265 283.925 96.525 ;
        RECT 289.125 96.465 289.445 96.525 ;
        RECT 290.965 96.465 291.285 96.525 ;
        RECT 294.200 96.465 294.490 96.510 ;
        RECT 289.125 96.325 294.490 96.465 ;
        RECT 289.125 96.265 289.445 96.325 ;
        RECT 290.965 96.265 291.285 96.325 ;
        RECT 294.200 96.280 294.490 96.325 ;
        RECT 284.065 96.125 284.385 96.185 ;
        RECT 283.235 95.985 284.385 96.125 ;
        RECT 284.065 95.925 284.385 95.985 ;
        RECT 291.885 95.925 292.205 96.185 ;
        RECT 292.345 96.125 292.665 96.185 ;
        RECT 298.340 96.125 298.630 96.170 ;
        RECT 292.345 95.985 298.630 96.125 ;
        RECT 292.345 95.925 292.665 95.985 ;
        RECT 298.340 95.940 298.630 95.985 ;
        RECT 302.005 95.925 302.325 96.185 ;
        RECT 162.095 95.305 311.935 95.785 ;
        RECT 177.345 94.905 177.665 95.165 ;
        RECT 184.705 95.105 185.025 95.165 ;
        RECT 186.100 95.105 186.390 95.150 ;
        RECT 184.705 94.965 186.390 95.105 ;
        RECT 184.705 94.905 185.025 94.965 ;
        RECT 186.100 94.920 186.390 94.965 ;
        RECT 188.400 94.920 188.690 95.150 ;
        RECT 190.240 95.105 190.530 95.150 ;
        RECT 192.065 95.105 192.385 95.165 ;
        RECT 190.240 94.965 192.385 95.105 ;
        RECT 190.240 94.920 190.530 94.965 ;
        RECT 170.000 94.765 170.290 94.810 ;
        RECT 171.365 94.765 171.685 94.825 ;
        RECT 170.000 94.625 171.685 94.765 ;
        RECT 170.000 94.580 170.290 94.625 ;
        RECT 171.365 94.565 171.685 94.625 ;
        RECT 172.280 94.765 172.930 94.810 ;
        RECT 173.205 94.765 173.525 94.825 ;
        RECT 175.880 94.765 176.170 94.810 ;
        RECT 172.280 94.625 176.170 94.765 ;
        RECT 172.280 94.580 172.930 94.625 ;
        RECT 173.205 94.565 173.525 94.625 ;
        RECT 175.580 94.580 176.170 94.625 ;
        RECT 163.545 94.225 163.865 94.485 ;
        RECT 165.400 94.425 165.690 94.470 ;
        RECT 165.845 94.425 166.165 94.485 ;
        RECT 165.400 94.285 166.165 94.425 ;
        RECT 165.400 94.240 165.690 94.285 ;
        RECT 165.845 94.225 166.165 94.285 ;
        RECT 169.085 94.425 169.375 94.470 ;
        RECT 170.920 94.425 171.210 94.470 ;
        RECT 174.500 94.425 174.790 94.470 ;
        RECT 169.085 94.285 174.790 94.425 ;
        RECT 169.085 94.240 169.375 94.285 ;
        RECT 170.920 94.240 171.210 94.285 ;
        RECT 174.500 94.240 174.790 94.285 ;
        RECT 175.580 94.265 175.870 94.580 ;
        RECT 177.805 94.425 178.125 94.485 ;
        RECT 187.020 94.425 187.310 94.470 ;
        RECT 188.475 94.425 188.615 94.920 ;
        RECT 192.065 94.905 192.385 94.965 ;
        RECT 201.265 94.905 201.585 95.165 ;
        RECT 215.065 95.105 215.385 95.165 ;
        RECT 219.205 95.105 219.525 95.165 ;
        RECT 215.065 94.965 219.525 95.105 ;
        RECT 215.065 94.905 215.385 94.965 ;
        RECT 219.205 94.905 219.525 94.965 ;
        RECT 219.665 94.905 219.985 95.165 ;
        RECT 220.140 94.920 220.430 95.150 ;
        RECT 221.045 95.105 221.365 95.165 ;
        RECT 221.045 94.965 221.735 95.105 ;
        RECT 190.700 94.765 190.990 94.810 ;
        RECT 200.345 94.765 200.665 94.825 ;
        RECT 177.805 94.285 186.775 94.425 ;
        RECT 177.805 94.225 178.125 94.285 ;
        RECT 168.620 94.085 168.910 94.130 ;
        RECT 184.245 94.085 184.565 94.145 ;
        RECT 168.620 93.945 184.565 94.085 ;
        RECT 186.635 94.085 186.775 94.285 ;
        RECT 187.020 94.285 188.615 94.425 ;
        RECT 188.935 94.625 200.665 94.765 ;
        RECT 187.020 94.240 187.310 94.285 ;
        RECT 188.935 94.085 189.075 94.625 ;
        RECT 190.700 94.580 190.990 94.625 ;
        RECT 200.345 94.565 200.665 94.625 ;
        RECT 192.525 94.425 192.845 94.485 ;
        RECT 193.460 94.425 193.750 94.470 ;
        RECT 194.825 94.425 195.145 94.485 ;
        RECT 192.525 94.285 193.215 94.425 ;
        RECT 192.525 94.225 192.845 94.285 ;
        RECT 186.635 93.945 189.075 94.085 ;
        RECT 191.620 94.085 191.910 94.130 ;
        RECT 192.065 94.085 192.385 94.145 ;
        RECT 191.620 93.945 192.385 94.085 ;
        RECT 168.620 93.900 168.910 93.945 ;
        RECT 165.385 93.745 165.705 93.805 ;
        RECT 168.695 93.745 168.835 93.900 ;
        RECT 184.245 93.885 184.565 93.945 ;
        RECT 191.620 93.900 191.910 93.945 ;
        RECT 192.065 93.885 192.385 93.945 ;
        RECT 165.385 93.605 168.835 93.745 ;
        RECT 169.490 93.745 169.780 93.790 ;
        RECT 171.380 93.745 171.670 93.790 ;
        RECT 174.500 93.745 174.790 93.790 ;
        RECT 169.490 93.605 174.790 93.745 ;
        RECT 193.075 93.745 193.215 94.285 ;
        RECT 193.460 94.285 195.145 94.425 ;
        RECT 201.355 94.425 201.495 94.905 ;
        RECT 201.725 94.765 202.045 94.825 ;
        RECT 219.755 94.765 219.895 94.905 ;
        RECT 201.725 94.625 219.895 94.765 ;
        RECT 220.215 94.765 220.355 94.920 ;
        RECT 221.045 94.905 221.365 94.965 ;
        RECT 220.215 94.625 221.300 94.765 ;
        RECT 201.725 94.565 202.045 94.625 ;
        RECT 202.200 94.425 202.490 94.470 ;
        RECT 201.355 94.285 202.490 94.425 ;
        RECT 193.460 94.240 193.750 94.285 ;
        RECT 194.825 94.225 195.145 94.285 ;
        RECT 202.200 94.240 202.490 94.285 ;
        RECT 203.105 94.425 203.425 94.485 ;
        RECT 208.625 94.425 208.945 94.485 ;
        RECT 203.105 94.285 208.945 94.425 ;
        RECT 203.105 94.225 203.425 94.285 ;
        RECT 208.625 94.225 208.945 94.285 ;
        RECT 216.445 94.425 216.765 94.485 ;
        RECT 217.455 94.470 217.595 94.625 ;
        RECT 216.920 94.425 217.210 94.470 ;
        RECT 216.445 94.285 217.210 94.425 ;
        RECT 216.445 94.225 216.765 94.285 ;
        RECT 216.920 94.240 217.210 94.285 ;
        RECT 217.385 94.240 217.675 94.470 ;
        RECT 218.285 94.225 218.605 94.485 ;
        RECT 218.745 94.225 219.065 94.485 ;
        RECT 219.665 94.470 219.985 94.485 ;
        RECT 219.450 94.240 219.985 94.470 ;
        RECT 219.665 94.225 219.985 94.240 ;
        RECT 220.125 94.425 220.445 94.485 ;
        RECT 220.600 94.425 220.890 94.470 ;
        RECT 220.125 94.285 220.890 94.425 ;
        RECT 220.125 94.225 220.445 94.285 ;
        RECT 220.600 94.240 220.890 94.285 ;
        RECT 221.160 94.085 221.300 94.625 ;
        RECT 221.595 94.470 221.735 94.965 ;
        RECT 222.425 94.905 222.745 95.165 ;
        RECT 227.945 95.105 228.265 95.165 ;
        RECT 238.525 95.105 238.845 95.165 ;
        RECT 242.665 95.105 242.985 95.165 ;
        RECT 222.975 94.965 224.495 95.105 ;
        RECT 222.975 94.765 223.115 94.965 ;
        RECT 223.805 94.810 224.125 94.825 ;
        RECT 222.055 94.625 223.115 94.765 ;
        RECT 221.520 94.240 221.810 94.470 ;
        RECT 222.055 94.085 222.195 94.625 ;
        RECT 223.690 94.580 224.125 94.810 ;
        RECT 224.355 94.765 224.495 94.965 ;
        RECT 227.945 94.965 237.375 95.105 ;
        RECT 227.945 94.905 228.265 94.965 ;
        RECT 226.580 94.765 226.870 94.810 ;
        RECT 229.785 94.765 230.105 94.825 ;
        RECT 224.355 94.625 226.870 94.765 ;
        RECT 226.580 94.580 226.870 94.625 ;
        RECT 227.575 94.625 230.105 94.765 ;
        RECT 223.805 94.565 224.125 94.580 ;
        RECT 224.280 94.425 224.570 94.470 ;
        RECT 222.560 94.285 224.570 94.425 ;
        RECT 222.560 94.145 222.700 94.285 ;
        RECT 224.280 94.240 224.570 94.285 ;
        RECT 224.725 94.225 225.045 94.485 ;
        RECT 227.575 94.470 227.715 94.625 ;
        RECT 229.785 94.565 230.105 94.625 ;
        RECT 234.845 94.765 235.165 94.825 ;
        RECT 237.235 94.810 237.375 94.965 ;
        RECT 238.525 94.965 242.985 95.105 ;
        RECT 238.525 94.905 238.845 94.965 ;
        RECT 242.665 94.905 242.985 94.965 ;
        RECT 243.140 94.920 243.430 95.150 ;
        RECT 243.585 95.105 243.905 95.165 ;
        RECT 261.080 95.105 261.370 95.150 ;
        RECT 264.745 95.105 265.065 95.165 ;
        RECT 243.585 94.965 246.575 95.105 ;
        RECT 237.160 94.765 237.450 94.810 ;
        RECT 234.845 94.625 236.460 94.765 ;
        RECT 234.845 94.565 235.165 94.625 ;
        RECT 225.200 94.425 225.490 94.470 ;
        RECT 225.200 94.345 225.875 94.425 ;
        RECT 226.425 94.345 227.285 94.375 ;
        RECT 225.200 94.285 227.285 94.345 ;
        RECT 225.200 94.240 225.490 94.285 ;
        RECT 225.735 94.235 227.285 94.285 ;
        RECT 227.500 94.240 227.790 94.470 ;
        RECT 227.960 94.425 228.250 94.470 ;
        RECT 232.545 94.425 232.865 94.485 ;
        RECT 235.765 94.425 236.085 94.485 ;
        RECT 236.320 94.470 236.460 94.625 ;
        RECT 237.160 94.625 239.675 94.765 ;
        RECT 237.160 94.580 237.450 94.625 ;
        RECT 239.535 94.485 239.675 94.625 ;
        RECT 241.745 94.565 242.065 94.825 ;
        RECT 227.960 94.285 236.085 94.425 ;
        RECT 227.960 94.240 228.250 94.285 ;
        RECT 225.735 94.205 226.565 94.235 ;
        RECT 221.160 93.945 222.195 94.085 ;
        RECT 222.425 93.885 222.745 94.145 ;
        RECT 222.885 93.885 223.205 94.145 ;
        RECT 201.280 93.745 201.570 93.790 ;
        RECT 193.075 93.605 201.570 93.745 ;
        RECT 165.385 93.545 165.705 93.605 ;
        RECT 169.490 93.560 169.780 93.605 ;
        RECT 171.380 93.560 171.670 93.605 ;
        RECT 174.500 93.560 174.790 93.605 ;
        RECT 201.280 93.560 201.570 93.605 ;
        RECT 208.165 93.745 208.485 93.805 ;
        RECT 209.085 93.745 209.405 93.805 ;
        RECT 208.165 93.605 209.405 93.745 ;
        RECT 208.165 93.545 208.485 93.605 ;
        RECT 209.085 93.545 209.405 93.605 ;
        RECT 213.685 93.745 214.005 93.805 ;
        RECT 222.515 93.745 222.655 93.885 ;
        RECT 213.685 93.605 222.655 93.745 ;
        RECT 227.145 93.745 227.285 94.235 ;
        RECT 232.545 94.225 232.865 94.285 ;
        RECT 235.765 94.225 236.085 94.285 ;
        RECT 236.245 94.240 236.535 94.470 ;
        RECT 237.605 94.225 237.925 94.485 ;
        RECT 238.065 94.470 238.385 94.485 ;
        RECT 238.065 94.425 238.395 94.470 ;
        RECT 238.065 94.285 238.580 94.425 ;
        RECT 238.065 94.240 238.395 94.285 ;
        RECT 238.065 94.225 238.385 94.240 ;
        RECT 239.445 94.225 239.765 94.485 ;
        RECT 239.905 94.225 240.225 94.485 ;
        RECT 242.205 94.470 242.525 94.485 ;
        RECT 240.385 94.240 240.675 94.470 ;
        RECT 241.300 94.425 241.590 94.470 ;
        RECT 240.915 94.285 241.590 94.425 ;
        RECT 235.305 94.085 235.625 94.145 ;
        RECT 240.460 94.085 240.600 94.240 ;
        RECT 235.305 93.945 240.600 94.085 ;
        RECT 235.305 93.885 235.625 93.945 ;
        RECT 240.915 93.805 241.055 94.285 ;
        RECT 241.300 94.240 241.590 94.285 ;
        RECT 242.205 94.425 242.535 94.470 ;
        RECT 243.215 94.425 243.355 94.920 ;
        RECT 243.585 94.905 243.905 94.965 ;
        RECT 244.965 94.565 245.285 94.825 ;
        RECT 243.585 94.425 243.905 94.485 ;
        RECT 242.205 94.285 242.720 94.425 ;
        RECT 243.215 94.285 243.905 94.425 ;
        RECT 242.205 94.240 242.535 94.285 ;
        RECT 242.205 94.225 242.525 94.240 ;
        RECT 243.585 94.225 243.905 94.285 ;
        RECT 244.045 94.425 244.365 94.485 ;
        RECT 246.435 94.470 246.575 94.965 ;
        RECT 261.080 94.965 265.065 95.105 ;
        RECT 261.080 94.920 261.370 94.965 ;
        RECT 264.745 94.905 265.065 94.965 ;
        RECT 282.685 94.905 283.005 95.165 ;
        RECT 283.145 94.905 283.465 95.165 ;
        RECT 283.605 95.105 283.925 95.165 ;
        RECT 289.585 95.105 289.905 95.165 ;
        RECT 283.605 94.965 289.905 95.105 ;
        RECT 283.605 94.905 283.925 94.965 ;
        RECT 289.585 94.905 289.905 94.965 ;
        RECT 290.505 94.905 290.825 95.165 ;
        RECT 291.885 94.905 292.205 95.165 ;
        RECT 302.005 95.105 302.325 95.165 ;
        RECT 298.875 94.965 302.325 95.105 ;
        RECT 262.460 94.765 262.750 94.810 ;
        RECT 256.555 94.625 262.750 94.765 ;
        RECT 244.520 94.425 244.810 94.470 ;
        RECT 244.045 94.285 244.810 94.425 ;
        RECT 244.045 94.225 244.365 94.285 ;
        RECT 244.520 94.240 244.810 94.285 ;
        RECT 245.440 94.240 245.730 94.470 ;
        RECT 246.360 94.240 246.650 94.470 ;
        RECT 244.965 94.085 245.285 94.145 ;
        RECT 245.515 94.085 245.655 94.240 ;
        RECT 256.555 94.145 256.695 94.625 ;
        RECT 262.460 94.580 262.750 94.625 ;
        RECT 278.175 94.625 281.075 94.765 ;
        RECT 278.175 94.485 278.315 94.625 ;
        RECT 257.845 94.225 258.165 94.485 ;
        RECT 258.765 94.470 259.085 94.485 ;
        RECT 258.600 94.240 259.085 94.470 ;
        RECT 258.765 94.225 259.085 94.240 ;
        RECT 259.225 94.225 259.545 94.485 ;
        RECT 260.145 94.470 260.465 94.485 ;
        RECT 259.700 94.240 259.990 94.470 ;
        RECT 260.145 94.240 260.570 94.470 ;
        RECT 255.545 94.085 255.865 94.145 ;
        RECT 242.755 93.945 243.355 94.085 ;
        RECT 238.065 93.745 238.385 93.805 ;
        RECT 227.145 93.605 238.385 93.745 ;
        RECT 213.685 93.545 214.005 93.605 ;
        RECT 238.065 93.545 238.385 93.605 ;
        RECT 240.825 93.545 241.145 93.805 ;
        RECT 241.745 93.745 242.065 93.805 ;
        RECT 242.755 93.745 242.895 93.945 ;
        RECT 241.745 93.605 242.895 93.745 ;
        RECT 243.215 93.745 243.355 93.945 ;
        RECT 244.965 93.945 255.865 94.085 ;
        RECT 244.965 93.885 245.285 93.945 ;
        RECT 255.545 93.885 255.865 93.945 ;
        RECT 256.465 93.885 256.785 94.145 ;
        RECT 259.775 94.085 259.915 94.240 ;
        RECT 260.145 94.225 260.465 94.240 ;
        RECT 261.525 94.225 261.845 94.485 ;
        RECT 262.905 94.225 263.225 94.485 ;
        RECT 263.380 94.240 263.670 94.470 ;
        RECT 268.885 94.425 269.205 94.485 ;
        RECT 277.640 94.425 277.930 94.470 ;
        RECT 268.885 94.285 277.930 94.425 ;
        RECT 258.395 93.945 259.915 94.085 ;
        RECT 262.445 94.085 262.765 94.145 ;
        RECT 263.455 94.085 263.595 94.240 ;
        RECT 268.885 94.225 269.205 94.285 ;
        RECT 277.640 94.240 277.930 94.285 ;
        RECT 278.085 94.225 278.405 94.485 ;
        RECT 279.005 94.425 279.325 94.485 ;
        RECT 279.005 94.285 280.155 94.425 ;
        RECT 279.005 94.225 279.325 94.285 ;
        RECT 271.185 94.085 271.505 94.145 ;
        RECT 262.445 93.945 271.505 94.085 ;
        RECT 280.015 94.085 280.155 94.285 ;
        RECT 280.385 94.225 280.705 94.485 ;
        RECT 280.935 94.470 281.075 94.625 ;
        RECT 280.860 94.240 281.150 94.470 ;
        RECT 281.780 94.425 282.070 94.470 ;
        RECT 281.395 94.285 282.070 94.425 ;
        RECT 282.775 94.425 282.915 94.905 ;
        RECT 284.080 94.425 284.370 94.470 ;
        RECT 282.775 94.285 284.370 94.425 ;
        RECT 281.395 94.085 281.535 94.285 ;
        RECT 281.780 94.240 282.070 94.285 ;
        RECT 284.080 94.240 284.370 94.285 ;
        RECT 289.600 94.425 289.890 94.470 ;
        RECT 291.975 94.425 292.115 94.905 ;
        RECT 292.920 94.765 293.210 94.810 ;
        RECT 295.105 94.765 295.425 94.825 ;
        RECT 298.875 94.810 299.015 94.965 ;
        RECT 302.005 94.905 302.325 94.965 ;
        RECT 303.845 94.905 304.165 95.165 ;
        RECT 296.160 94.765 296.810 94.810 ;
        RECT 292.920 94.625 296.810 94.765 ;
        RECT 292.920 94.580 293.510 94.625 ;
        RECT 289.600 94.285 292.115 94.425 ;
        RECT 289.600 94.240 289.890 94.285 ;
        RECT 293.220 94.265 293.510 94.580 ;
        RECT 295.105 94.565 295.425 94.625 ;
        RECT 296.160 94.580 296.810 94.625 ;
        RECT 298.800 94.580 299.090 94.810 ;
        RECT 303.385 94.765 303.705 94.825 ;
        RECT 300.715 94.625 303.705 94.765 ;
        RECT 303.935 94.765 304.075 94.905 ;
        RECT 304.300 94.765 304.950 94.810 ;
        RECT 307.900 94.765 308.190 94.810 ;
        RECT 303.935 94.625 308.190 94.765 ;
        RECT 300.715 94.485 300.855 94.625 ;
        RECT 303.385 94.565 303.705 94.625 ;
        RECT 304.300 94.580 304.950 94.625 ;
        RECT 307.600 94.580 308.190 94.625 ;
        RECT 294.300 94.425 294.590 94.470 ;
        RECT 297.880 94.425 298.170 94.470 ;
        RECT 299.715 94.425 300.005 94.470 ;
        RECT 294.300 94.285 300.005 94.425 ;
        RECT 294.300 94.240 294.590 94.285 ;
        RECT 297.880 94.240 298.170 94.285 ;
        RECT 299.715 94.240 300.005 94.285 ;
        RECT 300.180 94.425 300.470 94.470 ;
        RECT 300.625 94.425 300.945 94.485 ;
        RECT 300.180 94.285 300.945 94.425 ;
        RECT 300.180 94.240 300.470 94.285 ;
        RECT 300.625 94.225 300.945 94.285 ;
        RECT 301.105 94.425 301.395 94.470 ;
        RECT 302.940 94.425 303.230 94.470 ;
        RECT 306.520 94.425 306.810 94.470 ;
        RECT 301.105 94.285 306.810 94.425 ;
        RECT 301.105 94.240 301.395 94.285 ;
        RECT 302.940 94.240 303.230 94.285 ;
        RECT 306.520 94.240 306.810 94.285 ;
        RECT 307.600 94.265 307.890 94.580 ;
        RECT 280.015 93.945 281.535 94.085 ;
        RECT 282.225 94.085 282.545 94.145 ;
        RECT 282.700 94.085 282.990 94.130 ;
        RECT 292.805 94.085 293.125 94.145 ;
        RECT 282.225 93.945 282.990 94.085 ;
        RECT 243.600 93.745 243.890 93.790 ;
        RECT 256.555 93.745 256.695 93.885 ;
        RECT 258.395 93.805 258.535 93.945 ;
        RECT 262.445 93.885 262.765 93.945 ;
        RECT 271.185 93.885 271.505 93.945 ;
        RECT 282.225 93.885 282.545 93.945 ;
        RECT 282.700 93.900 282.990 93.945 ;
        RECT 283.465 93.945 293.125 94.085 ;
        RECT 243.215 93.605 243.890 93.745 ;
        RECT 241.745 93.545 242.065 93.605 ;
        RECT 243.600 93.560 243.890 93.605 ;
        RECT 244.135 93.605 256.695 93.745 ;
        RECT 192.525 93.205 192.845 93.465 ;
        RECT 197.125 93.405 197.445 93.465 ;
        RECT 215.525 93.405 215.845 93.465 ;
        RECT 218.745 93.405 219.065 93.465 ;
        RECT 197.125 93.265 219.065 93.405 ;
        RECT 197.125 93.205 197.445 93.265 ;
        RECT 215.525 93.205 215.845 93.265 ;
        RECT 218.745 93.205 219.065 93.265 ;
        RECT 221.045 93.205 221.365 93.465 ;
        RECT 226.120 93.405 226.410 93.450 ;
        RECT 226.580 93.405 226.870 93.450 ;
        RECT 226.120 93.265 226.870 93.405 ;
        RECT 226.120 93.220 226.410 93.265 ;
        RECT 226.580 93.220 226.870 93.265 ;
        RECT 228.865 93.205 229.185 93.465 ;
        RECT 238.985 93.205 239.305 93.465 ;
        RECT 240.915 93.405 241.055 93.545 ;
        RECT 244.135 93.405 244.275 93.605 ;
        RECT 258.305 93.545 258.625 93.805 ;
        RECT 259.225 93.745 259.545 93.805 ;
        RECT 260.605 93.745 260.925 93.805 ;
        RECT 278.545 93.745 278.865 93.805 ;
        RECT 259.225 93.605 260.925 93.745 ;
        RECT 259.225 93.545 259.545 93.605 ;
        RECT 260.605 93.545 260.925 93.605 ;
        RECT 262.995 93.605 278.865 93.745 ;
        RECT 240.915 93.265 244.275 93.405 ;
        RECT 247.265 93.405 247.585 93.465 ;
        RECT 262.995 93.405 263.135 93.605 ;
        RECT 278.545 93.545 278.865 93.605 ;
        RECT 279.940 93.745 280.230 93.790 ;
        RECT 281.765 93.745 282.085 93.805 ;
        RECT 283.465 93.745 283.605 93.945 ;
        RECT 292.805 93.885 293.125 93.945 ;
        RECT 302.005 93.885 302.325 94.145 ;
        RECT 294.300 93.745 294.590 93.790 ;
        RECT 297.420 93.745 297.710 93.790 ;
        RECT 299.310 93.745 299.600 93.790 ;
        RECT 279.940 93.605 283.605 93.745 ;
        RECT 291.055 93.605 293.955 93.745 ;
        RECT 279.940 93.560 280.230 93.605 ;
        RECT 281.765 93.545 282.085 93.605 ;
        RECT 247.265 93.265 263.135 93.405 ;
        RECT 247.265 93.205 247.585 93.265 ;
        RECT 264.285 93.205 264.605 93.465 ;
        RECT 278.635 93.405 278.775 93.545 ;
        RECT 291.055 93.405 291.195 93.605 ;
        RECT 293.815 93.465 293.955 93.605 ;
        RECT 294.300 93.605 299.600 93.745 ;
        RECT 294.300 93.560 294.590 93.605 ;
        RECT 297.420 93.560 297.710 93.605 ;
        RECT 299.310 93.560 299.600 93.605 ;
        RECT 301.510 93.745 301.800 93.790 ;
        RECT 303.400 93.745 303.690 93.790 ;
        RECT 306.520 93.745 306.810 93.790 ;
        RECT 301.510 93.605 306.810 93.745 ;
        RECT 301.510 93.560 301.800 93.605 ;
        RECT 303.400 93.560 303.690 93.605 ;
        RECT 306.520 93.560 306.810 93.605 ;
        RECT 278.635 93.265 291.195 93.405 ;
        RECT 291.440 93.405 291.730 93.450 ;
        RECT 292.345 93.405 292.665 93.465 ;
        RECT 291.440 93.265 292.665 93.405 ;
        RECT 291.440 93.220 291.730 93.265 ;
        RECT 292.345 93.205 292.665 93.265 ;
        RECT 293.725 93.205 294.045 93.465 ;
        RECT 296.945 93.405 297.265 93.465 ;
        RECT 302.925 93.405 303.245 93.465 ;
        RECT 309.380 93.405 309.670 93.450 ;
        RECT 296.945 93.265 309.670 93.405 ;
        RECT 296.945 93.205 297.265 93.265 ;
        RECT 302.925 93.205 303.245 93.265 ;
        RECT 309.380 93.220 309.670 93.265 ;
        RECT 162.095 92.585 311.135 93.065 ;
        RECT 165.845 92.385 166.165 92.445 ;
        RECT 174.125 92.385 174.445 92.445 ;
        RECT 175.520 92.385 175.810 92.430 ;
        RECT 209.085 92.385 209.405 92.445 ;
        RECT 165.845 92.245 172.055 92.385 ;
        RECT 165.845 92.185 166.165 92.245 ;
        RECT 166.270 92.045 166.560 92.090 ;
        RECT 168.160 92.045 168.450 92.090 ;
        RECT 171.280 92.045 171.570 92.090 ;
        RECT 166.270 91.905 171.570 92.045 ;
        RECT 171.915 92.045 172.055 92.245 ;
        RECT 174.125 92.245 175.810 92.385 ;
        RECT 174.125 92.185 174.445 92.245 ;
        RECT 175.520 92.200 175.810 92.245 ;
        RECT 183.875 92.245 209.405 92.385 ;
        RECT 183.875 92.045 184.015 92.245 ;
        RECT 209.085 92.185 209.405 92.245 ;
        RECT 216.445 92.385 216.765 92.445 ;
        RECT 217.380 92.385 217.670 92.430 ;
        RECT 216.445 92.245 217.670 92.385 ;
        RECT 216.445 92.185 216.765 92.245 ;
        RECT 217.380 92.200 217.670 92.245 ;
        RECT 220.585 92.385 220.905 92.445 ;
        RECT 226.565 92.385 226.885 92.445 ;
        RECT 220.585 92.245 226.885 92.385 ;
        RECT 220.585 92.185 220.905 92.245 ;
        RECT 226.565 92.185 226.885 92.245 ;
        RECT 227.945 92.185 228.265 92.445 ;
        RECT 239.905 92.385 240.225 92.445 ;
        RECT 241.300 92.385 241.590 92.430 ;
        RECT 239.905 92.245 241.590 92.385 ;
        RECT 239.905 92.185 240.225 92.245 ;
        RECT 241.300 92.200 241.590 92.245 ;
        RECT 241.745 92.185 242.065 92.445 ;
        RECT 244.505 92.385 244.825 92.445 ;
        RECT 279.465 92.385 279.785 92.445 ;
        RECT 244.505 92.245 279.785 92.385 ;
        RECT 244.505 92.185 244.825 92.245 ;
        RECT 279.465 92.185 279.785 92.245 ;
        RECT 193.445 92.045 193.765 92.105 ;
        RECT 171.915 91.905 184.015 92.045 ;
        RECT 184.795 91.905 193.765 92.045 ;
        RECT 166.270 91.860 166.560 91.905 ;
        RECT 168.160 91.860 168.450 91.905 ;
        RECT 171.280 91.860 171.570 91.905 ;
        RECT 165.385 91.505 165.705 91.765 ;
        RECT 166.780 91.705 167.070 91.750 ;
        RECT 169.985 91.705 170.305 91.765 ;
        RECT 166.780 91.565 170.305 91.705 ;
        RECT 166.780 91.520 167.070 91.565 ;
        RECT 169.985 91.505 170.305 91.565 ;
        RECT 177.805 91.505 178.125 91.765 ;
        RECT 178.725 91.705 179.045 91.765 ;
        RECT 184.795 91.750 184.935 91.905 ;
        RECT 193.445 91.845 193.765 91.905 ;
        RECT 193.920 92.045 194.210 92.090 ;
        RECT 194.825 92.045 195.145 92.105 ;
        RECT 204.485 92.045 204.805 92.105 ;
        RECT 229.785 92.045 230.105 92.105 ;
        RECT 193.920 91.905 195.145 92.045 ;
        RECT 193.920 91.860 194.210 91.905 ;
        RECT 194.825 91.845 195.145 91.905 ;
        RECT 196.755 91.905 197.815 92.045 ;
        RECT 184.720 91.705 185.010 91.750 ;
        RECT 178.725 91.565 185.010 91.705 ;
        RECT 178.725 91.505 179.045 91.565 ;
        RECT 184.720 91.520 185.010 91.565 ;
        RECT 185.180 91.705 185.470 91.750 ;
        RECT 186.085 91.705 186.405 91.765 ;
        RECT 185.180 91.565 186.405 91.705 ;
        RECT 185.180 91.520 185.470 91.565 ;
        RECT 186.085 91.505 186.405 91.565 ;
        RECT 190.225 91.705 190.545 91.765 ;
        RECT 191.160 91.705 191.450 91.750 ;
        RECT 190.225 91.565 191.450 91.705 ;
        RECT 190.225 91.505 190.545 91.565 ;
        RECT 191.160 91.520 191.450 91.565 ;
        RECT 192.065 91.705 192.385 91.765 ;
        RECT 196.755 91.750 196.895 91.905 ;
        RECT 196.680 91.705 196.970 91.750 ;
        RECT 192.065 91.565 196.970 91.705 ;
        RECT 197.675 91.705 197.815 91.905 ;
        RECT 204.485 91.905 230.105 92.045 ;
        RECT 204.485 91.845 204.805 91.905 ;
        RECT 229.785 91.845 230.105 91.905 ;
        RECT 238.985 91.845 239.305 92.105 ;
        RECT 240.365 92.045 240.685 92.105 ;
        RECT 262.445 92.045 262.765 92.105 ;
        RECT 239.995 91.905 260.835 92.045 ;
        RECT 205.880 91.705 206.170 91.750 ;
        RECT 206.800 91.705 207.090 91.750 ;
        RECT 197.675 91.565 207.090 91.705 ;
        RECT 192.065 91.505 192.385 91.565 ;
        RECT 196.680 91.520 196.970 91.565 ;
        RECT 205.880 91.520 206.170 91.565 ;
        RECT 206.800 91.520 207.090 91.565 ;
        RECT 208.625 91.505 208.945 91.765 ;
        RECT 209.100 91.705 209.390 91.750 ;
        RECT 209.545 91.705 209.865 91.765 ;
        RECT 219.665 91.705 219.985 91.765 ;
        RECT 209.100 91.565 219.985 91.705 ;
        RECT 209.100 91.520 209.390 91.565 ;
        RECT 209.545 91.505 209.865 91.565 ;
        RECT 219.665 91.505 219.985 91.565 ;
        RECT 222.055 91.565 232.315 91.705 ;
        RECT 165.865 91.365 166.155 91.410 ;
        RECT 167.700 91.365 167.990 91.410 ;
        RECT 171.280 91.365 171.570 91.410 ;
        RECT 165.865 91.225 171.570 91.365 ;
        RECT 165.865 91.180 166.155 91.225 ;
        RECT 167.700 91.180 167.990 91.225 ;
        RECT 171.280 91.180 171.570 91.225 ;
        RECT 172.360 91.365 172.650 91.385 ;
        RECT 173.205 91.365 173.525 91.425 ;
        RECT 182.865 91.365 183.185 91.425 ;
        RECT 194.365 91.365 194.685 91.425 ;
        RECT 199.900 91.365 200.190 91.410 ;
        RECT 201.265 91.365 201.585 91.425 ;
        RECT 172.360 91.225 183.185 91.365 ;
        RECT 172.360 91.070 172.650 91.225 ;
        RECT 173.205 91.165 173.525 91.225 ;
        RECT 182.865 91.165 183.185 91.225 ;
        RECT 187.095 91.225 190.455 91.365 ;
        RECT 169.060 91.025 169.710 91.070 ;
        RECT 172.360 91.025 172.950 91.070 ;
        RECT 169.060 90.885 172.950 91.025 ;
        RECT 169.060 90.840 169.710 90.885 ;
        RECT 172.660 90.840 172.950 90.885 ;
        RECT 177.345 90.825 177.665 91.085 ;
        RECT 179.185 91.025 179.505 91.085 ;
        RECT 187.095 91.025 187.235 91.225 ;
        RECT 189.305 91.025 189.625 91.085 ;
        RECT 179.185 90.885 187.235 91.025 ;
        RECT 187.555 90.885 189.625 91.025 ;
        RECT 179.185 90.825 179.505 90.885 ;
        RECT 173.665 90.685 173.985 90.745 ;
        RECT 174.140 90.685 174.430 90.730 ;
        RECT 177.435 90.685 177.575 90.825 ;
        RECT 173.665 90.545 177.575 90.685 ;
        RECT 185.640 90.685 185.930 90.730 ;
        RECT 186.545 90.685 186.865 90.745 ;
        RECT 187.555 90.730 187.695 90.885 ;
        RECT 189.305 90.825 189.625 90.885 ;
        RECT 185.640 90.545 186.865 90.685 ;
        RECT 173.665 90.485 173.985 90.545 ;
        RECT 174.140 90.500 174.430 90.545 ;
        RECT 185.640 90.500 185.930 90.545 ;
        RECT 186.545 90.485 186.865 90.545 ;
        RECT 187.480 90.500 187.770 90.730 ;
        RECT 188.845 90.485 189.165 90.745 ;
        RECT 190.315 90.685 190.455 91.225 ;
        RECT 194.365 91.225 201.585 91.365 ;
        RECT 194.365 91.165 194.685 91.225 ;
        RECT 199.900 91.180 200.190 91.225 ;
        RECT 201.265 91.165 201.585 91.225 ;
        RECT 204.485 91.165 204.805 91.425 ;
        RECT 207.705 91.165 208.025 91.425 ;
        RECT 213.240 91.365 213.530 91.410 ;
        RECT 216.460 91.365 216.750 91.410 ;
        RECT 220.585 91.365 220.905 91.425 ;
        RECT 222.055 91.365 222.195 91.565 ;
        RECT 213.240 91.225 220.905 91.365 ;
        RECT 213.240 91.180 213.530 91.225 ;
        RECT 216.460 91.180 216.750 91.225 ;
        RECT 220.585 91.165 220.905 91.225 ;
        RECT 221.160 91.225 222.195 91.365 ;
        RECT 222.440 91.365 222.730 91.410 ;
        RECT 227.025 91.365 227.345 91.425 ;
        RECT 229.800 91.365 230.090 91.410 ;
        RECT 222.440 91.225 230.090 91.365 ;
        RECT 190.700 91.025 190.990 91.070 ;
        RECT 192.985 91.025 193.305 91.085 ;
        RECT 196.220 91.025 196.510 91.070 ;
        RECT 190.700 90.885 193.305 91.025 ;
        RECT 190.700 90.840 190.990 90.885 ;
        RECT 192.985 90.825 193.305 90.885 ;
        RECT 195.375 90.885 196.510 91.025 ;
        RECT 194.825 90.685 195.145 90.745 ;
        RECT 195.375 90.685 195.515 90.885 ;
        RECT 196.220 90.840 196.510 90.885 ;
        RECT 198.045 90.825 198.365 91.085 ;
        RECT 198.505 91.025 198.825 91.085 ;
        RECT 204.945 91.025 205.265 91.085 ;
        RECT 198.505 90.885 205.265 91.025 ;
        RECT 198.505 90.825 198.825 90.885 ;
        RECT 204.945 90.825 205.265 90.885 ;
        RECT 213.685 91.025 214.005 91.085 ;
        RECT 214.620 91.025 214.910 91.070 ;
        RECT 215.540 91.025 215.830 91.070 ;
        RECT 213.685 90.885 214.910 91.025 ;
        RECT 213.685 90.825 214.005 90.885 ;
        RECT 214.620 90.840 214.910 90.885 ;
        RECT 215.155 90.885 215.830 91.025 ;
        RECT 215.155 90.745 215.295 90.885 ;
        RECT 215.540 90.840 215.830 90.885 ;
        RECT 216.000 91.025 216.290 91.070 ;
        RECT 216.905 91.025 217.225 91.085 ;
        RECT 221.160 91.025 221.300 91.225 ;
        RECT 222.440 91.180 222.730 91.225 ;
        RECT 227.025 91.165 227.345 91.225 ;
        RECT 229.800 91.180 230.090 91.225 ;
        RECT 232.175 91.085 232.315 91.565 ;
        RECT 234.385 91.165 234.705 91.425 ;
        RECT 234.845 91.365 235.165 91.425 ;
        RECT 238.080 91.365 238.370 91.410 ;
        RECT 234.845 91.225 238.370 91.365 ;
        RECT 239.075 91.365 239.215 91.845 ;
        RECT 239.995 91.750 240.135 91.905 ;
        RECT 240.365 91.845 240.685 91.905 ;
        RECT 239.920 91.520 240.210 91.750 ;
        RECT 242.220 91.705 242.510 91.750 ;
        RECT 243.125 91.705 243.445 91.765 ;
        RECT 242.220 91.565 243.445 91.705 ;
        RECT 242.220 91.520 242.510 91.565 ;
        RECT 243.125 91.505 243.445 91.565 ;
        RECT 251.955 91.565 260.375 91.705 ;
        RECT 251.955 91.425 252.095 91.565 ;
        RECT 241.785 91.365 242.075 91.410 ;
        RECT 239.075 91.225 242.075 91.365 ;
        RECT 234.845 91.165 235.165 91.225 ;
        RECT 238.080 91.180 238.370 91.225 ;
        RECT 241.785 91.180 242.075 91.225 ;
        RECT 242.665 91.365 242.985 91.425 ;
        RECT 246.345 91.365 246.665 91.425 ;
        RECT 242.665 91.225 246.665 91.365 ;
        RECT 242.665 91.165 242.985 91.225 ;
        RECT 246.345 91.165 246.665 91.225 ;
        RECT 251.865 91.165 252.185 91.425 ;
        RECT 259.225 91.365 259.545 91.425 ;
        RECT 260.235 91.410 260.375 91.565 ;
        RECT 259.700 91.365 259.990 91.410 ;
        RECT 259.225 91.225 259.990 91.365 ;
        RECT 259.225 91.165 259.545 91.225 ;
        RECT 259.700 91.180 259.990 91.225 ;
        RECT 260.160 91.180 260.450 91.410 ;
        RECT 216.000 90.885 221.300 91.025 ;
        RECT 216.000 90.840 216.290 90.885 ;
        RECT 216.905 90.825 217.225 90.885 ;
        RECT 221.505 90.825 221.825 91.085 ;
        RECT 227.960 91.025 228.250 91.070 ;
        RECT 223.895 90.885 228.250 91.025 ;
        RECT 223.895 90.745 224.035 90.885 ;
        RECT 227.960 90.840 228.250 90.885 ;
        RECT 232.085 90.825 232.405 91.085 ;
        RECT 190.315 90.545 195.515 90.685 ;
        RECT 195.760 90.685 196.050 90.730 ;
        RECT 197.125 90.685 197.445 90.745 ;
        RECT 195.760 90.545 197.445 90.685 ;
        RECT 194.825 90.485 195.145 90.545 ;
        RECT 195.760 90.500 196.050 90.545 ;
        RECT 197.125 90.485 197.445 90.545 ;
        RECT 202.645 90.485 202.965 90.745 ;
        RECT 215.065 90.485 215.385 90.745 ;
        RECT 219.665 90.485 219.985 90.745 ;
        RECT 221.060 90.685 221.350 90.730 ;
        RECT 223.805 90.685 224.125 90.745 ;
        RECT 221.060 90.545 224.125 90.685 ;
        RECT 221.060 90.500 221.350 90.545 ;
        RECT 223.805 90.485 224.125 90.545 ;
        RECT 224.265 90.485 224.585 90.745 ;
        RECT 226.565 90.685 226.885 90.745 ;
        RECT 227.040 90.685 227.330 90.730 ;
        RECT 234.475 90.685 234.615 91.165 ;
        RECT 238.525 91.025 238.845 91.085 ;
        RECT 240.505 91.025 240.795 91.070 ;
        RECT 238.525 90.885 240.795 91.025 ;
        RECT 260.695 91.025 260.835 91.905 ;
        RECT 262.445 91.905 288.895 92.045 ;
        RECT 262.445 91.845 262.765 91.905 ;
        RECT 277.255 91.565 279.235 91.705 ;
        RECT 261.065 91.165 261.385 91.425 ;
        RECT 261.540 91.365 261.830 91.410 ;
        RECT 264.285 91.365 264.605 91.425 ;
        RECT 261.540 91.225 264.605 91.365 ;
        RECT 261.540 91.180 261.830 91.225 ;
        RECT 264.285 91.165 264.605 91.225 ;
        RECT 277.255 91.025 277.395 91.565 ;
        RECT 277.640 91.365 277.930 91.410 ;
        RECT 279.095 91.365 279.235 91.565 ;
        RECT 281.765 91.505 282.085 91.765 ;
        RECT 277.640 91.225 278.775 91.365 ;
        RECT 279.095 91.225 280.615 91.365 ;
        RECT 277.640 91.180 277.930 91.225 ;
        RECT 260.695 90.885 277.395 91.025 ;
        RECT 238.525 90.825 238.845 90.885 ;
        RECT 240.505 90.840 240.795 90.885 ;
        RECT 226.565 90.545 234.615 90.685 ;
        RECT 226.565 90.485 226.885 90.545 ;
        RECT 227.040 90.500 227.330 90.545 ;
        RECT 239.445 90.485 239.765 90.745 ;
        RECT 243.600 90.685 243.890 90.730 ;
        RECT 248.185 90.685 248.505 90.745 ;
        RECT 243.600 90.545 248.505 90.685 ;
        RECT 243.600 90.500 243.890 90.545 ;
        RECT 248.185 90.485 248.505 90.545 ;
        RECT 258.780 90.685 259.070 90.730 ;
        RECT 269.345 90.685 269.665 90.745 ;
        RECT 258.780 90.545 269.665 90.685 ;
        RECT 258.780 90.500 259.070 90.545 ;
        RECT 269.345 90.485 269.665 90.545 ;
        RECT 276.705 90.485 277.025 90.745 ;
        RECT 278.635 90.730 278.775 91.225 ;
        RECT 279.465 90.825 279.785 91.085 ;
        RECT 280.475 91.070 280.615 91.225 ;
        RECT 282.685 91.165 283.005 91.425 ;
        RECT 280.400 91.025 280.690 91.070 ;
        RECT 284.985 91.025 285.305 91.085 ;
        RECT 280.400 90.885 285.305 91.025 ;
        RECT 288.755 91.025 288.895 91.905 ;
        RECT 299.720 91.860 300.010 92.090 ;
        RECT 301.100 92.045 301.390 92.090 ;
        RECT 301.545 92.045 301.865 92.105 ;
        RECT 301.100 91.905 301.865 92.045 ;
        RECT 301.100 91.860 301.390 91.905 ;
        RECT 289.125 91.705 289.445 91.765 ;
        RECT 292.820 91.705 293.110 91.750 ;
        RECT 295.565 91.705 295.885 91.765 ;
        RECT 296.500 91.705 296.790 91.750 ;
        RECT 289.125 91.565 296.790 91.705 ;
        RECT 289.125 91.505 289.445 91.565 ;
        RECT 292.820 91.520 293.110 91.565 ;
        RECT 295.565 91.505 295.885 91.565 ;
        RECT 296.500 91.520 296.790 91.565 ;
        RECT 297.420 91.705 297.710 91.750 ;
        RECT 297.865 91.705 298.185 91.765 ;
        RECT 297.420 91.565 298.185 91.705 ;
        RECT 297.420 91.520 297.710 91.565 ;
        RECT 297.865 91.505 298.185 91.565 ;
        RECT 290.965 91.365 291.285 91.425 ;
        RECT 292.360 91.365 292.650 91.410 ;
        RECT 290.965 91.225 292.650 91.365 ;
        RECT 299.795 91.365 299.935 91.860 ;
        RECT 301.545 91.845 301.865 91.905 ;
        RECT 300.180 91.365 300.470 91.410 ;
        RECT 299.795 91.225 300.470 91.365 ;
        RECT 290.965 91.165 291.285 91.225 ;
        RECT 292.360 91.180 292.650 91.225 ;
        RECT 300.180 91.180 300.470 91.225 ;
        RECT 302.465 91.165 302.785 91.425 ;
        RECT 291.885 91.025 292.205 91.085 ;
        RECT 302.555 91.025 302.695 91.165 ;
        RECT 288.755 90.885 291.195 91.025 ;
        RECT 280.400 90.840 280.690 90.885 ;
        RECT 284.985 90.825 285.305 90.885 ;
        RECT 278.560 90.500 278.850 90.730 ;
        RECT 279.555 90.685 279.695 90.825 ;
        RECT 280.860 90.685 281.150 90.730 ;
        RECT 283.145 90.685 283.465 90.745 ;
        RECT 279.555 90.545 283.465 90.685 ;
        RECT 280.860 90.500 281.150 90.545 ;
        RECT 283.145 90.485 283.465 90.545 ;
        RECT 283.620 90.685 283.910 90.730 ;
        RECT 284.525 90.685 284.845 90.745 ;
        RECT 283.620 90.545 284.845 90.685 ;
        RECT 283.620 90.500 283.910 90.545 ;
        RECT 284.525 90.485 284.845 90.545 ;
        RECT 290.045 90.485 290.365 90.745 ;
        RECT 291.055 90.685 291.195 90.885 ;
        RECT 291.885 90.885 302.695 91.025 ;
        RECT 291.885 90.825 292.205 90.885 ;
        RECT 297.880 90.685 298.170 90.730 ;
        RECT 308.445 90.685 308.765 90.745 ;
        RECT 291.055 90.545 308.765 90.685 ;
        RECT 297.880 90.500 298.170 90.545 ;
        RECT 308.445 90.485 308.765 90.545 ;
        RECT 162.095 89.865 311.935 90.345 ;
        RECT 181.945 89.665 182.265 89.725 ;
        RECT 184.720 89.665 185.010 89.710 ;
        RECT 181.945 89.525 185.010 89.665 ;
        RECT 181.945 89.465 182.265 89.525 ;
        RECT 184.720 89.480 185.010 89.525 ;
        RECT 188.845 89.465 189.165 89.725 ;
        RECT 189.305 89.465 189.625 89.725 ;
        RECT 191.605 89.665 191.925 89.725 ;
        RECT 198.045 89.665 198.365 89.725 ;
        RECT 191.605 89.525 198.365 89.665 ;
        RECT 191.605 89.465 191.925 89.525 ;
        RECT 198.045 89.465 198.365 89.525 ;
        RECT 202.645 89.465 202.965 89.725 ;
        RECT 204.485 89.665 204.805 89.725 ;
        RECT 210.020 89.665 210.310 89.710 ;
        RECT 204.485 89.525 210.310 89.665 ;
        RECT 204.485 89.465 204.805 89.525 ;
        RECT 210.020 89.480 210.310 89.525 ;
        RECT 211.860 89.665 212.150 89.710 ;
        RECT 213.685 89.665 214.005 89.725 ;
        RECT 211.860 89.525 214.005 89.665 ;
        RECT 211.860 89.480 212.150 89.525 ;
        RECT 213.685 89.465 214.005 89.525 ;
        RECT 215.525 89.665 215.845 89.725 ;
        RECT 219.220 89.665 219.510 89.710 ;
        RECT 215.525 89.525 219.510 89.665 ;
        RECT 215.525 89.465 215.845 89.525 ;
        RECT 219.220 89.480 219.510 89.525 ;
        RECT 219.665 89.465 219.985 89.725 ;
        RECT 220.125 89.665 220.445 89.725 ;
        RECT 222.440 89.665 222.730 89.710 ;
        RECT 220.125 89.525 222.730 89.665 ;
        RECT 220.125 89.465 220.445 89.525 ;
        RECT 222.440 89.480 222.730 89.525 ;
        RECT 223.345 89.665 223.665 89.725 ;
        RECT 223.820 89.665 224.110 89.710 ;
        RECT 242.665 89.665 242.985 89.725 ;
        RECT 258.765 89.665 259.085 89.725 ;
        RECT 262.445 89.665 262.765 89.725 ;
        RECT 223.345 89.525 224.110 89.665 ;
        RECT 223.345 89.465 223.665 89.525 ;
        RECT 223.820 89.480 224.110 89.525 ;
        RECT 238.155 89.525 257.615 89.665 ;
        RECT 169.980 89.325 170.630 89.370 ;
        RECT 173.580 89.325 173.870 89.370 ;
        RECT 169.980 89.185 173.870 89.325 ;
        RECT 169.980 89.140 170.630 89.185 ;
        RECT 173.280 89.140 173.870 89.185 ;
        RECT 179.640 89.325 180.290 89.370 ;
        RECT 183.240 89.325 183.530 89.370 ;
        RECT 179.640 89.185 183.530 89.325 ;
        RECT 179.640 89.140 180.290 89.185 ;
        RECT 182.940 89.140 183.530 89.185 ;
        RECT 173.280 89.045 173.570 89.140 ;
        RECT 164.925 88.785 165.245 89.045 ;
        RECT 165.385 88.985 165.705 89.045 ;
        RECT 166.320 88.985 166.610 89.030 ;
        RECT 165.385 88.845 166.610 88.985 ;
        RECT 165.385 88.785 165.705 88.845 ;
        RECT 166.320 88.800 166.610 88.845 ;
        RECT 166.785 88.985 167.075 89.030 ;
        RECT 168.620 88.985 168.910 89.030 ;
        RECT 172.200 88.985 172.490 89.030 ;
        RECT 166.785 88.845 172.490 88.985 ;
        RECT 166.785 88.800 167.075 88.845 ;
        RECT 168.620 88.800 168.910 88.845 ;
        RECT 172.200 88.800 172.490 88.845 ;
        RECT 173.205 88.825 173.570 89.045 ;
        RECT 176.445 88.985 176.735 89.030 ;
        RECT 178.280 88.985 178.570 89.030 ;
        RECT 181.860 88.985 182.150 89.030 ;
        RECT 176.445 88.845 182.150 88.985 ;
        RECT 173.205 88.785 173.525 88.825 ;
        RECT 176.445 88.800 176.735 88.845 ;
        RECT 178.280 88.800 178.570 88.845 ;
        RECT 181.860 88.800 182.150 88.845 ;
        RECT 182.940 88.825 183.230 89.140 ;
        RECT 187.480 88.985 187.770 89.030 ;
        RECT 188.935 88.985 189.075 89.465 ;
        RECT 189.395 89.030 189.535 89.465 ;
        RECT 191.160 89.325 191.450 89.370 ;
        RECT 192.525 89.325 192.845 89.385 ;
        RECT 191.160 89.185 192.845 89.325 ;
        RECT 191.160 89.140 191.450 89.185 ;
        RECT 192.525 89.125 192.845 89.185 ;
        RECT 193.440 89.325 194.090 89.370 ;
        RECT 197.040 89.325 197.330 89.370 ;
        RECT 198.135 89.325 198.275 89.465 ;
        RECT 202.735 89.325 202.875 89.465 ;
        RECT 193.440 89.185 198.275 89.325 ;
        RECT 199.975 89.185 202.875 89.325 ;
        RECT 204.940 89.325 205.590 89.370 ;
        RECT 208.540 89.325 208.830 89.370 ;
        RECT 204.940 89.185 208.830 89.325 ;
        RECT 219.755 89.325 219.895 89.465 ;
        RECT 221.045 89.325 221.365 89.385 ;
        RECT 226.580 89.325 226.870 89.370 ;
        RECT 219.755 89.185 220.815 89.325 ;
        RECT 193.440 89.140 194.090 89.185 ;
        RECT 196.740 89.140 197.330 89.185 ;
        RECT 187.480 88.845 189.075 88.985 ;
        RECT 167.700 88.645 167.990 88.690 ;
        RECT 165.935 88.505 167.990 88.645 ;
        RECT 165.935 88.350 166.075 88.505 ;
        RECT 167.700 88.460 167.990 88.505 ;
        RECT 168.145 88.645 168.465 88.705 ;
        RECT 172.745 88.645 173.065 88.705 ;
        RECT 168.145 88.505 173.205 88.645 ;
        RECT 168.145 88.445 168.465 88.505 ;
        RECT 172.745 88.445 173.205 88.505 ;
        RECT 175.980 88.460 176.270 88.690 ;
        RECT 165.860 88.120 166.150 88.350 ;
        RECT 167.190 88.305 167.480 88.350 ;
        RECT 169.080 88.305 169.370 88.350 ;
        RECT 172.200 88.305 172.490 88.350 ;
        RECT 167.190 88.165 172.490 88.305 ;
        RECT 173.065 88.305 173.205 88.445 ;
        RECT 175.045 88.305 175.365 88.365 ;
        RECT 173.065 88.165 175.365 88.305 ;
        RECT 167.190 88.120 167.480 88.165 ;
        RECT 169.080 88.120 169.370 88.165 ;
        RECT 172.200 88.120 172.490 88.165 ;
        RECT 175.045 88.105 175.365 88.165 ;
        RECT 176.055 87.965 176.195 88.460 ;
        RECT 177.345 88.445 177.665 88.705 ;
        RECT 182.955 88.365 183.095 88.825 ;
        RECT 187.480 88.800 187.770 88.845 ;
        RECT 189.320 88.800 189.610 89.030 ;
        RECT 190.245 88.985 190.535 89.030 ;
        RECT 192.080 88.985 192.370 89.030 ;
        RECT 195.660 88.985 195.950 89.030 ;
        RECT 190.245 88.845 195.950 88.985 ;
        RECT 190.245 88.800 190.535 88.845 ;
        RECT 192.080 88.800 192.370 88.845 ;
        RECT 195.660 88.800 195.950 88.845 ;
        RECT 196.740 88.825 197.030 89.140 ;
        RECT 199.975 89.030 200.115 89.185 ;
        RECT 204.940 89.140 205.590 89.185 ;
        RECT 208.240 89.140 208.830 89.185 ;
        RECT 208.240 89.045 208.530 89.140 ;
        RECT 199.900 88.800 200.190 89.030 ;
        RECT 201.745 88.985 202.035 89.030 ;
        RECT 203.580 88.985 203.870 89.030 ;
        RECT 207.160 88.985 207.450 89.030 ;
        RECT 201.745 88.845 207.450 88.985 ;
        RECT 201.745 88.800 202.035 88.845 ;
        RECT 203.580 88.800 203.870 88.845 ;
        RECT 207.160 88.800 207.450 88.845 ;
        RECT 208.165 88.825 208.530 89.045 ;
        RECT 209.085 88.985 209.405 89.045 ;
        RECT 210.940 88.985 211.230 89.030 ;
        RECT 211.385 88.985 211.705 89.045 ;
        RECT 220.675 89.030 220.815 89.185 ;
        RECT 221.045 89.185 226.870 89.325 ;
        RECT 221.045 89.125 221.365 89.185 ;
        RECT 226.580 89.140 226.870 89.185 ;
        RECT 209.085 88.845 211.705 88.985 ;
        RECT 208.165 88.785 208.485 88.825 ;
        RECT 209.085 88.785 209.405 88.845 ;
        RECT 210.940 88.800 211.230 88.845 ;
        RECT 211.385 88.785 211.705 88.845 ;
        RECT 218.760 88.800 219.050 89.030 ;
        RECT 220.600 88.800 220.890 89.030 ;
        RECT 223.345 88.985 223.665 89.045 ;
        RECT 226.105 88.985 226.425 89.045 ;
        RECT 223.345 88.845 226.425 88.985 ;
        RECT 226.655 88.985 226.795 89.140 ;
        RECT 227.945 88.985 228.265 89.045 ;
        RECT 236.240 88.985 236.530 89.030 ;
        RECT 226.655 88.845 228.265 88.985 ;
        RECT 188.845 88.645 189.165 88.705 ;
        RECT 189.780 88.645 190.070 88.690 ;
        RECT 191.605 88.645 191.925 88.705 ;
        RECT 188.845 88.505 190.070 88.645 ;
        RECT 188.845 88.445 189.165 88.505 ;
        RECT 189.780 88.460 190.070 88.505 ;
        RECT 190.315 88.505 191.925 88.645 ;
        RECT 176.850 88.305 177.140 88.350 ;
        RECT 178.740 88.305 179.030 88.350 ;
        RECT 181.860 88.305 182.150 88.350 ;
        RECT 176.850 88.165 182.150 88.305 ;
        RECT 176.850 88.120 177.140 88.165 ;
        RECT 178.740 88.120 179.030 88.165 ;
        RECT 181.860 88.120 182.150 88.165 ;
        RECT 182.865 88.305 183.185 88.365 ;
        RECT 190.315 88.305 190.455 88.505 ;
        RECT 191.605 88.445 191.925 88.505 ;
        RECT 197.125 88.645 197.445 88.705 ;
        RECT 198.520 88.645 198.810 88.690 ;
        RECT 197.125 88.505 198.810 88.645 ;
        RECT 197.125 88.445 197.445 88.505 ;
        RECT 198.520 88.460 198.810 88.505 ;
        RECT 200.805 88.645 201.125 88.705 ;
        RECT 201.280 88.645 201.570 88.690 ;
        RECT 202.660 88.645 202.950 88.690 ;
        RECT 200.805 88.505 201.570 88.645 ;
        RECT 200.805 88.445 201.125 88.505 ;
        RECT 201.280 88.460 201.570 88.505 ;
        RECT 201.815 88.505 202.950 88.645 ;
        RECT 182.865 88.165 190.455 88.305 ;
        RECT 190.650 88.305 190.940 88.350 ;
        RECT 192.540 88.305 192.830 88.350 ;
        RECT 195.660 88.305 195.950 88.350 ;
        RECT 201.815 88.305 201.955 88.505 ;
        RECT 202.660 88.460 202.950 88.505 ;
        RECT 206.325 88.645 206.645 88.705 ;
        RECT 216.905 88.645 217.225 88.705 ;
        RECT 206.325 88.505 217.225 88.645 ;
        RECT 218.835 88.645 218.975 88.800 ;
        RECT 223.345 88.785 223.665 88.845 ;
        RECT 226.105 88.785 226.425 88.845 ;
        RECT 227.945 88.785 228.265 88.845 ;
        RECT 234.015 88.845 236.530 88.985 ;
        RECT 234.015 88.705 234.155 88.845 ;
        RECT 236.240 88.800 236.530 88.845 ;
        RECT 236.685 88.785 237.005 89.045 ;
        RECT 237.145 88.985 237.465 89.045 ;
        RECT 238.155 89.030 238.295 89.525 ;
        RECT 242.665 89.465 242.985 89.525 ;
        RECT 239.000 89.325 239.290 89.370 ;
        RECT 242.205 89.325 242.525 89.385 ;
        RECT 256.940 89.325 257.230 89.370 ;
        RECT 239.000 89.185 241.515 89.325 ;
        RECT 239.000 89.140 239.290 89.185 ;
        RECT 237.620 88.985 237.910 89.030 ;
        RECT 237.145 88.845 237.910 88.985 ;
        RECT 237.145 88.785 237.465 88.845 ;
        RECT 237.620 88.800 237.910 88.845 ;
        RECT 238.080 88.800 238.370 89.030 ;
        RECT 239.920 88.985 240.210 89.030 ;
        RECT 240.365 88.985 240.685 89.045 ;
        RECT 241.375 89.030 241.515 89.185 ;
        RECT 242.205 89.185 242.895 89.325 ;
        RECT 242.205 89.125 242.525 89.185 ;
        RECT 242.755 89.030 242.895 89.185 ;
        RECT 254.255 89.185 257.230 89.325 ;
        RECT 239.920 88.845 240.685 88.985 ;
        RECT 239.920 88.800 240.210 88.845 ;
        RECT 240.365 88.785 240.685 88.845 ;
        RECT 240.840 88.800 241.130 89.030 ;
        RECT 241.300 88.800 241.590 89.030 ;
        RECT 241.760 88.985 242.050 89.030 ;
        RECT 242.680 88.985 242.970 89.030 ;
        RECT 243.125 88.985 243.445 89.045 ;
        RECT 241.760 88.845 242.435 88.985 ;
        RECT 241.760 88.800 242.050 88.845 ;
        RECT 221.045 88.645 221.365 88.705 ;
        RECT 218.835 88.505 221.365 88.645 ;
        RECT 206.325 88.445 206.645 88.505 ;
        RECT 216.905 88.445 217.225 88.505 ;
        RECT 221.045 88.445 221.365 88.505 ;
        RECT 224.280 88.645 224.570 88.690 ;
        RECT 230.245 88.645 230.565 88.705 ;
        RECT 224.280 88.505 230.565 88.645 ;
        RECT 224.280 88.460 224.570 88.505 ;
        RECT 230.245 88.445 230.565 88.505 ;
        RECT 233.925 88.445 234.245 88.705 ;
        RECT 240.915 88.645 241.055 88.800 ;
        RECT 240.915 88.505 241.975 88.645 ;
        RECT 241.835 88.365 241.975 88.505 ;
        RECT 242.295 88.365 242.435 88.845 ;
        RECT 242.680 88.845 243.445 88.985 ;
        RECT 242.680 88.800 242.970 88.845 ;
        RECT 243.125 88.785 243.445 88.845 ;
        RECT 253.245 88.985 253.565 89.045 ;
        RECT 254.255 89.030 254.395 89.185 ;
        RECT 256.940 89.140 257.230 89.185 ;
        RECT 257.475 89.045 257.615 89.525 ;
        RECT 258.765 89.525 262.765 89.665 ;
        RECT 258.765 89.465 259.085 89.525 ;
        RECT 258.305 89.125 258.625 89.385 ;
        RECT 253.720 88.985 254.010 89.030 ;
        RECT 253.245 88.845 254.010 88.985 ;
        RECT 253.245 88.785 253.565 88.845 ;
        RECT 253.720 88.800 254.010 88.845 ;
        RECT 254.180 88.800 254.470 89.030 ;
        RECT 255.085 88.785 255.405 89.045 ;
        RECT 255.560 88.985 255.850 89.030 ;
        RECT 257.385 88.985 257.705 89.045 ;
        RECT 255.560 88.845 257.705 88.985 ;
        RECT 255.560 88.800 255.850 88.845 ;
        RECT 257.385 88.785 257.705 88.845 ;
        RECT 257.845 88.785 258.165 89.045 ;
        RECT 260.235 89.030 260.375 89.525 ;
        RECT 262.445 89.465 262.765 89.525 ;
        RECT 262.905 89.465 263.225 89.725 ;
        RECT 274.865 89.665 275.185 89.725 ;
        RECT 282.685 89.665 283.005 89.725 ;
        RECT 284.080 89.665 284.370 89.710 ;
        RECT 274.865 89.525 278.315 89.665 ;
        RECT 274.865 89.465 275.185 89.525 ;
        RECT 260.605 89.325 260.925 89.385 ;
        RECT 262.000 89.325 262.290 89.370 ;
        RECT 260.605 89.185 262.290 89.325 ;
        RECT 262.995 89.325 263.135 89.465 ;
        RECT 262.995 89.185 269.805 89.325 ;
        RECT 260.605 89.125 260.925 89.185 ;
        RECT 262.000 89.140 262.290 89.185 ;
        RECT 258.785 88.985 259.075 89.030 ;
        RECT 259.370 88.985 259.660 89.030 ;
        RECT 258.675 88.800 259.075 88.985 ;
        RECT 259.320 88.800 259.660 88.985 ;
        RECT 260.160 88.800 260.450 89.030 ;
        RECT 261.540 88.985 261.830 89.030 ;
        RECT 260.695 88.845 261.830 88.985 ;
        RECT 255.175 88.645 255.315 88.785 ;
        RECT 256.465 88.645 256.785 88.705 ;
        RECT 258.675 88.645 258.815 88.800 ;
        RECT 243.215 88.505 255.315 88.645 ;
        RECT 256.095 88.505 258.815 88.645 ;
        RECT 190.650 88.165 195.950 88.305 ;
        RECT 182.865 88.105 183.185 88.165 ;
        RECT 190.650 88.120 190.940 88.165 ;
        RECT 192.540 88.120 192.830 88.165 ;
        RECT 195.660 88.120 195.950 88.165 ;
        RECT 200.895 88.165 201.955 88.305 ;
        RECT 202.150 88.305 202.440 88.350 ;
        RECT 204.040 88.305 204.330 88.350 ;
        RECT 207.160 88.305 207.450 88.350 ;
        RECT 202.150 88.165 207.450 88.305 ;
        RECT 184.245 87.965 184.565 88.025 ;
        RECT 176.055 87.825 184.565 87.965 ;
        RECT 184.245 87.765 184.565 87.825 ;
        RECT 185.625 87.965 185.945 88.025 ;
        RECT 186.560 87.965 186.850 88.010 ;
        RECT 185.625 87.825 186.850 87.965 ;
        RECT 185.625 87.765 185.945 87.825 ;
        RECT 186.560 87.780 186.850 87.825 ;
        RECT 188.385 87.765 188.705 88.025 ;
        RECT 200.895 88.010 201.035 88.165 ;
        RECT 202.150 88.120 202.440 88.165 ;
        RECT 204.040 88.120 204.330 88.165 ;
        RECT 207.160 88.120 207.450 88.165 ;
        RECT 220.140 88.305 220.430 88.350 ;
        RECT 222.900 88.305 223.190 88.350 ;
        RECT 220.140 88.165 223.190 88.305 ;
        RECT 220.140 88.120 220.430 88.165 ;
        RECT 222.900 88.120 223.190 88.165 ;
        RECT 224.725 88.305 225.045 88.365 ;
        RECT 226.580 88.305 226.870 88.350 ;
        RECT 227.025 88.305 227.345 88.365 ;
        RECT 224.725 88.165 226.335 88.305 ;
        RECT 224.725 88.105 225.045 88.165 ;
        RECT 226.195 88.025 226.335 88.165 ;
        RECT 226.580 88.165 227.345 88.305 ;
        RECT 226.580 88.120 226.870 88.165 ;
        RECT 227.025 88.105 227.345 88.165 ;
        RECT 229.785 88.105 230.105 88.365 ;
        RECT 232.085 88.305 232.405 88.365 ;
        RECT 237.145 88.305 237.465 88.365 ;
        RECT 239.445 88.305 239.765 88.365 ;
        RECT 232.085 88.165 239.765 88.305 ;
        RECT 232.085 88.105 232.405 88.165 ;
        RECT 237.145 88.105 237.465 88.165 ;
        RECT 239.445 88.105 239.765 88.165 ;
        RECT 241.745 88.105 242.065 88.365 ;
        RECT 242.205 88.105 242.525 88.365 ;
        RECT 200.820 87.780 201.110 88.010 ;
        RECT 221.060 87.965 221.350 88.010 ;
        RECT 223.345 87.965 223.665 88.025 ;
        RECT 221.060 87.825 223.665 87.965 ;
        RECT 221.060 87.780 221.350 87.825 ;
        RECT 223.345 87.765 223.665 87.825 ;
        RECT 226.105 87.765 226.425 88.025 ;
        RECT 229.875 87.965 230.015 88.105 ;
        RECT 243.215 87.965 243.355 88.505 ;
        RECT 244.505 88.305 244.825 88.365 ;
        RECT 256.095 88.305 256.235 88.505 ;
        RECT 256.465 88.445 256.785 88.505 ;
        RECT 258.305 88.305 258.625 88.365 ;
        RECT 244.505 88.165 256.235 88.305 ;
        RECT 256.555 88.165 258.625 88.305 ;
        RECT 259.320 88.305 259.460 88.800 ;
        RECT 260.695 88.705 260.835 88.845 ;
        RECT 261.540 88.800 261.830 88.845 ;
        RECT 262.445 88.785 262.765 89.045 ;
        RECT 263.915 89.030 264.055 89.185 ;
        RECT 263.050 88.800 263.340 89.030 ;
        RECT 263.840 88.800 264.130 89.030 ;
        RECT 265.680 88.800 265.970 89.030 ;
        RECT 266.125 88.985 266.445 89.045 ;
        RECT 266.600 88.985 266.890 89.030 ;
        RECT 266.125 88.845 266.890 88.985 ;
        RECT 260.605 88.445 260.925 88.705 ;
        RECT 263.125 88.645 263.265 88.800 ;
        RECT 261.155 88.505 263.265 88.645 ;
        RECT 261.155 88.305 261.295 88.505 ;
        RECT 259.320 88.165 261.295 88.305 ;
        RECT 244.505 88.105 244.825 88.165 ;
        RECT 229.875 87.825 243.355 87.965 ;
        RECT 243.600 87.965 243.890 88.010 ;
        RECT 244.965 87.965 245.285 88.025 ;
        RECT 256.555 88.010 256.695 88.165 ;
        RECT 258.305 88.105 258.625 88.165 ;
        RECT 261.155 88.025 261.295 88.165 ;
        RECT 265.755 88.025 265.895 88.800 ;
        RECT 266.125 88.785 266.445 88.845 ;
        RECT 266.600 88.800 266.890 88.845 ;
        RECT 243.600 87.825 245.285 87.965 ;
        RECT 243.600 87.780 243.890 87.825 ;
        RECT 244.965 87.765 245.285 87.825 ;
        RECT 256.480 87.780 256.770 88.010 ;
        RECT 256.925 87.965 257.245 88.025 ;
        RECT 260.620 87.965 260.910 88.010 ;
        RECT 256.925 87.825 260.910 87.965 ;
        RECT 256.925 87.765 257.245 87.825 ;
        RECT 260.620 87.780 260.910 87.825 ;
        RECT 261.065 87.765 261.385 88.025 ;
        RECT 265.665 87.765 265.985 88.025 ;
        RECT 267.520 87.965 267.810 88.010 ;
        RECT 268.425 87.965 268.745 88.025 ;
        RECT 267.520 87.825 268.745 87.965 ;
        RECT 269.665 87.965 269.805 89.185 ;
        RECT 270.725 89.125 271.045 89.385 ;
        RECT 274.420 89.325 274.710 89.370 ;
        RECT 277.625 89.325 277.945 89.385 ;
        RECT 274.420 89.185 277.945 89.325 ;
        RECT 278.175 89.325 278.315 89.525 ;
        RECT 282.685 89.525 284.370 89.665 ;
        RECT 282.685 89.465 283.005 89.525 ;
        RECT 284.080 89.480 284.370 89.525 ;
        RECT 286.825 89.665 287.145 89.725 ;
        RECT 286.825 89.525 300.855 89.665 ;
        RECT 286.825 89.465 287.145 89.525 ;
        RECT 278.540 89.325 279.190 89.370 ;
        RECT 282.140 89.325 282.430 89.370 ;
        RECT 278.175 89.185 282.430 89.325 ;
        RECT 274.420 89.140 274.710 89.185 ;
        RECT 277.625 89.125 277.945 89.185 ;
        RECT 278.540 89.140 279.190 89.185 ;
        RECT 281.840 89.140 282.430 89.185 ;
        RECT 283.145 89.325 283.465 89.385 ;
        RECT 286.380 89.325 286.670 89.370 ;
        RECT 283.145 89.185 286.670 89.325 ;
        RECT 275.345 88.985 275.635 89.030 ;
        RECT 277.180 88.985 277.470 89.030 ;
        RECT 280.760 88.985 281.050 89.030 ;
        RECT 275.345 88.845 281.050 88.985 ;
        RECT 275.345 88.800 275.635 88.845 ;
        RECT 277.180 88.800 277.470 88.845 ;
        RECT 280.760 88.800 281.050 88.845 ;
        RECT 281.840 88.825 282.130 89.140 ;
        RECT 283.145 89.125 283.465 89.185 ;
        RECT 286.380 89.140 286.670 89.185 ;
        RECT 290.045 89.125 290.365 89.385 ;
        RECT 285.905 88.985 286.225 89.045 ;
        RECT 288.205 88.985 288.525 89.045 ;
        RECT 285.905 88.845 288.525 88.985 ;
        RECT 285.905 88.785 286.225 88.845 ;
        RECT 288.205 88.785 288.525 88.845 ;
        RECT 289.600 88.985 289.890 89.030 ;
        RECT 290.135 88.985 290.275 89.125 ;
        RECT 291.515 89.030 291.655 89.525 ;
        RECT 295.105 89.370 295.425 89.385 ;
        RECT 295.100 89.325 295.750 89.370 ;
        RECT 298.700 89.325 298.990 89.370 ;
        RECT 295.100 89.185 298.990 89.325 ;
        RECT 295.100 89.140 295.750 89.185 ;
        RECT 298.400 89.140 298.990 89.185 ;
        RECT 295.105 89.125 295.425 89.140 ;
        RECT 289.600 88.845 290.275 88.985 ;
        RECT 289.600 88.800 289.890 88.845 ;
        RECT 291.440 88.800 291.730 89.030 ;
        RECT 291.905 88.985 292.195 89.030 ;
        RECT 293.740 88.985 294.030 89.030 ;
        RECT 297.320 88.985 297.610 89.030 ;
        RECT 291.905 88.845 297.610 88.985 ;
        RECT 291.905 88.800 292.195 88.845 ;
        RECT 293.740 88.800 294.030 88.845 ;
        RECT 297.320 88.800 297.610 88.845 ;
        RECT 298.400 88.825 298.690 89.140 ;
        RECT 300.715 89.045 300.855 89.525 ;
        RECT 303.845 89.465 304.165 89.725 ;
        RECT 308.445 89.665 308.765 89.725 ;
        RECT 309.380 89.665 309.670 89.710 ;
        RECT 308.445 89.525 309.670 89.665 ;
        RECT 308.445 89.465 308.765 89.525 ;
        RECT 309.380 89.480 309.670 89.525 ;
        RECT 301.545 89.325 301.865 89.385 ;
        RECT 302.020 89.325 302.310 89.370 ;
        RECT 301.545 89.185 302.310 89.325 ;
        RECT 303.935 89.325 304.075 89.465 ;
        RECT 304.300 89.325 304.950 89.370 ;
        RECT 307.900 89.325 308.190 89.370 ;
        RECT 303.935 89.185 308.190 89.325 ;
        RECT 301.545 89.125 301.865 89.185 ;
        RECT 302.020 89.140 302.310 89.185 ;
        RECT 304.300 89.140 304.950 89.185 ;
        RECT 307.600 89.140 308.190 89.185 ;
        RECT 300.625 88.785 300.945 89.045 ;
        RECT 301.105 88.985 301.395 89.030 ;
        RECT 302.940 88.985 303.230 89.030 ;
        RECT 306.520 88.985 306.810 89.030 ;
        RECT 301.105 88.845 306.810 88.985 ;
        RECT 301.105 88.800 301.395 88.845 ;
        RECT 302.940 88.800 303.230 88.845 ;
        RECT 306.520 88.800 306.810 88.845 ;
        RECT 307.600 88.825 307.890 89.140 ;
        RECT 274.865 88.445 275.185 88.705 ;
        RECT 276.260 88.645 276.550 88.690 ;
        RECT 276.705 88.645 277.025 88.705 ;
        RECT 286.365 88.645 286.685 88.705 ;
        RECT 276.260 88.505 277.025 88.645 ;
        RECT 276.260 88.460 276.550 88.505 ;
        RECT 276.705 88.445 277.025 88.505 ;
        RECT 282.315 88.505 286.685 88.645 ;
        RECT 275.750 88.305 276.040 88.350 ;
        RECT 277.640 88.305 277.930 88.350 ;
        RECT 280.760 88.305 281.050 88.350 ;
        RECT 275.750 88.165 281.050 88.305 ;
        RECT 275.750 88.120 276.040 88.165 ;
        RECT 277.640 88.120 277.930 88.165 ;
        RECT 280.760 88.120 281.050 88.165 ;
        RECT 282.315 87.965 282.455 88.505 ;
        RECT 286.365 88.445 286.685 88.505 ;
        RECT 286.840 88.645 287.130 88.690 ;
        RECT 289.125 88.645 289.445 88.705 ;
        RECT 292.820 88.645 293.110 88.690 ;
        RECT 286.840 88.505 289.445 88.645 ;
        RECT 286.840 88.460 287.130 88.505 ;
        RECT 282.685 88.305 283.005 88.365 ;
        RECT 286.915 88.305 287.055 88.460 ;
        RECT 289.125 88.445 289.445 88.505 ;
        RECT 290.595 88.505 293.110 88.645 ;
        RECT 290.595 88.350 290.735 88.505 ;
        RECT 292.820 88.460 293.110 88.505 ;
        RECT 300.180 88.645 300.470 88.690 ;
        RECT 302.465 88.645 302.785 88.705 ;
        RECT 300.180 88.505 302.785 88.645 ;
        RECT 300.180 88.460 300.470 88.505 ;
        RECT 302.465 88.445 302.785 88.505 ;
        RECT 282.685 88.165 287.055 88.305 ;
        RECT 282.685 88.105 283.005 88.165 ;
        RECT 290.520 88.120 290.810 88.350 ;
        RECT 292.310 88.305 292.600 88.350 ;
        RECT 294.200 88.305 294.490 88.350 ;
        RECT 297.320 88.305 297.610 88.350 ;
        RECT 292.310 88.165 297.610 88.305 ;
        RECT 292.310 88.120 292.600 88.165 ;
        RECT 294.200 88.120 294.490 88.165 ;
        RECT 297.320 88.120 297.610 88.165 ;
        RECT 301.510 88.305 301.800 88.350 ;
        RECT 303.400 88.305 303.690 88.350 ;
        RECT 306.520 88.305 306.810 88.350 ;
        RECT 301.510 88.165 306.810 88.305 ;
        RECT 301.510 88.120 301.800 88.165 ;
        RECT 303.400 88.120 303.690 88.165 ;
        RECT 306.520 88.120 306.810 88.165 ;
        RECT 269.665 87.825 282.455 87.965 ;
        RECT 283.620 87.965 283.910 88.010 ;
        RECT 284.985 87.965 285.305 88.025 ;
        RECT 283.620 87.825 285.305 87.965 ;
        RECT 267.520 87.780 267.810 87.825 ;
        RECT 268.425 87.765 268.745 87.825 ;
        RECT 283.620 87.780 283.910 87.825 ;
        RECT 284.985 87.765 285.305 87.825 ;
        RECT 293.725 87.965 294.045 88.025 ;
        RECT 300.165 87.965 300.485 88.025 ;
        RECT 293.725 87.825 300.485 87.965 ;
        RECT 293.725 87.765 294.045 87.825 ;
        RECT 300.165 87.765 300.485 87.825 ;
        RECT 162.095 87.145 311.135 87.625 ;
        RECT 164.925 86.945 165.245 87.005 ;
        RECT 170.920 86.945 171.210 86.990 ;
        RECT 164.925 86.805 171.210 86.945 ;
        RECT 164.925 86.745 165.245 86.805 ;
        RECT 170.920 86.760 171.210 86.805 ;
        RECT 175.965 86.945 176.285 87.005 ;
        RECT 182.405 86.945 182.725 87.005 ;
        RECT 175.965 86.805 182.725 86.945 ;
        RECT 175.965 86.745 176.285 86.805 ;
        RECT 182.405 86.745 182.725 86.805 ;
        RECT 188.845 86.945 189.165 87.005 ;
        RECT 200.805 86.945 201.125 87.005 ;
        RECT 207.705 86.945 208.025 87.005 ;
        RECT 188.845 86.805 201.125 86.945 ;
        RECT 188.845 86.745 189.165 86.805 ;
        RECT 200.805 86.745 201.125 86.805 ;
        RECT 202.275 86.805 208.025 86.945 ;
        RECT 170.460 86.605 170.750 86.650 ;
        RECT 177.345 86.605 177.665 86.665 ;
        RECT 170.460 86.465 177.665 86.605 ;
        RECT 170.460 86.420 170.750 86.465 ;
        RECT 177.345 86.405 177.665 86.465 ;
        RECT 185.130 86.605 185.420 86.650 ;
        RECT 187.020 86.605 187.310 86.650 ;
        RECT 190.140 86.605 190.430 86.650 ;
        RECT 185.130 86.465 190.430 86.605 ;
        RECT 185.130 86.420 185.420 86.465 ;
        RECT 187.020 86.420 187.310 86.465 ;
        RECT 190.140 86.420 190.430 86.465 ;
        RECT 193.905 86.605 194.225 86.665 ;
        RECT 201.280 86.605 201.570 86.650 ;
        RECT 193.905 86.465 201.570 86.605 ;
        RECT 193.905 86.405 194.225 86.465 ;
        RECT 201.280 86.420 201.570 86.465 ;
        RECT 174.140 86.265 174.430 86.310 ;
        RECT 178.725 86.265 179.045 86.325 ;
        RECT 174.140 86.125 179.045 86.265 ;
        RECT 174.140 86.080 174.430 86.125 ;
        RECT 178.725 86.065 179.045 86.125 ;
        RECT 184.245 86.265 184.565 86.325 ;
        RECT 186.085 86.265 186.405 86.325 ;
        RECT 184.245 86.125 186.405 86.265 ;
        RECT 184.245 86.065 184.565 86.125 ;
        RECT 186.085 86.065 186.405 86.125 ;
        RECT 169.540 85.740 169.830 85.970 ;
        RECT 169.615 85.245 169.755 85.740 ;
        RECT 172.745 85.725 173.065 85.985 ;
        RECT 173.220 85.925 173.510 85.970 ;
        RECT 177.360 85.925 177.650 85.970 ;
        RECT 181.945 85.925 182.265 85.985 ;
        RECT 173.220 85.785 177.115 85.925 ;
        RECT 173.220 85.740 173.510 85.785 ;
        RECT 176.975 85.585 177.115 85.785 ;
        RECT 177.360 85.785 182.265 85.925 ;
        RECT 177.360 85.740 177.650 85.785 ;
        RECT 181.945 85.725 182.265 85.785 ;
        RECT 184.725 85.925 185.015 85.970 ;
        RECT 186.560 85.925 186.850 85.970 ;
        RECT 190.140 85.925 190.430 85.970 ;
        RECT 184.725 85.785 190.430 85.925 ;
        RECT 184.725 85.740 185.015 85.785 ;
        RECT 186.560 85.740 186.850 85.785 ;
        RECT 190.140 85.740 190.430 85.785 ;
        RECT 191.220 85.925 191.510 85.945 ;
        RECT 194.365 85.925 194.685 85.985 ;
        RECT 202.275 85.970 202.415 86.805 ;
        RECT 207.705 86.745 208.025 86.805 ;
        RECT 208.625 86.745 208.945 87.005 ;
        RECT 222.900 86.945 223.195 87.000 ;
        RECT 225.660 86.945 225.955 87.000 ;
        RECT 222.900 86.805 225.955 86.945 ;
        RECT 222.900 86.730 223.195 86.805 ;
        RECT 225.660 86.730 225.955 86.805 ;
        RECT 226.120 86.945 226.410 86.990 ;
        RECT 226.565 86.945 226.885 87.005 ;
        RECT 236.685 86.945 237.005 87.005 ;
        RECT 238.540 86.945 238.830 86.990 ;
        RECT 244.505 86.945 244.825 87.005 ;
        RECT 226.120 86.805 234.155 86.945 ;
        RECT 226.120 86.760 226.410 86.805 ;
        RECT 226.565 86.745 226.885 86.805 ;
        RECT 234.015 86.665 234.155 86.805 ;
        RECT 236.685 86.805 238.830 86.945 ;
        RECT 236.685 86.745 237.005 86.805 ;
        RECT 238.540 86.760 238.830 86.805 ;
        RECT 240.455 86.805 244.825 86.945 ;
        RECT 212.320 86.605 212.610 86.650 ;
        RECT 222.425 86.605 222.745 86.665 ;
        RECT 203.655 86.465 222.745 86.605 ;
        RECT 203.655 86.310 203.795 86.465 ;
        RECT 212.320 86.420 212.610 86.465 ;
        RECT 222.425 86.405 222.745 86.465 ;
        RECT 229.785 86.605 230.105 86.665 ;
        RECT 233.005 86.605 233.325 86.665 ;
        RECT 229.785 86.465 233.325 86.605 ;
        RECT 229.785 86.405 230.105 86.465 ;
        RECT 233.005 86.405 233.325 86.465 ;
        RECT 233.925 86.405 234.245 86.665 ;
        RECT 239.445 86.605 239.765 86.665 ;
        RECT 239.445 86.465 240.135 86.605 ;
        RECT 239.445 86.405 239.765 86.465 ;
        RECT 203.580 86.080 203.870 86.310 ;
        RECT 205.880 86.265 206.170 86.310 ;
        RECT 225.200 86.265 225.490 86.310 ;
        RECT 227.485 86.265 227.805 86.325 ;
        RECT 237.605 86.265 237.925 86.325 ;
        RECT 205.880 86.125 210.235 86.265 ;
        RECT 205.880 86.080 206.170 86.125 ;
        RECT 191.220 85.785 194.685 85.925 ;
        RECT 182.035 85.585 182.175 85.725 ;
        RECT 184.245 85.585 184.565 85.645 ;
        RECT 173.065 85.445 175.735 85.585 ;
        RECT 176.975 85.445 181.715 85.585 ;
        RECT 182.035 85.445 184.565 85.585 ;
        RECT 173.065 85.245 173.205 85.445 ;
        RECT 175.595 85.290 175.735 85.445 ;
        RECT 169.615 85.105 173.205 85.245 ;
        RECT 175.520 85.060 175.810 85.290 ;
        RECT 177.820 85.245 178.110 85.290 ;
        RECT 179.185 85.245 179.505 85.305 ;
        RECT 177.820 85.105 179.505 85.245 ;
        RECT 181.575 85.245 181.715 85.445 ;
        RECT 184.245 85.385 184.565 85.445 ;
        RECT 185.625 85.385 185.945 85.645 ;
        RECT 191.220 85.630 191.510 85.785 ;
        RECT 194.365 85.725 194.685 85.785 ;
        RECT 202.200 85.740 202.490 85.970 ;
        RECT 203.105 85.725 203.425 85.985 ;
        RECT 206.325 85.725 206.645 85.985 ;
        RECT 206.785 85.725 207.105 85.985 ;
        RECT 207.720 85.925 208.010 85.970 ;
        RECT 208.625 85.925 208.945 85.985 ;
        RECT 209.560 85.925 209.850 85.970 ;
        RECT 207.720 85.785 208.945 85.925 ;
        RECT 207.720 85.740 208.010 85.785 ;
        RECT 208.625 85.725 208.945 85.785 ;
        RECT 209.175 85.785 209.850 85.925 ;
        RECT 187.920 85.585 188.570 85.630 ;
        RECT 191.220 85.585 191.810 85.630 ;
        RECT 187.920 85.445 191.810 85.585 ;
        RECT 187.920 85.400 188.570 85.445 ;
        RECT 191.520 85.400 191.810 85.445 ;
        RECT 204.485 85.585 204.805 85.645 ;
        RECT 204.960 85.585 205.250 85.630 ;
        RECT 204.485 85.445 206.555 85.585 ;
        RECT 204.485 85.385 204.805 85.445 ;
        RECT 204.960 85.400 205.250 85.445 ;
        RECT 190.225 85.245 190.545 85.305 ;
        RECT 181.575 85.105 190.545 85.245 ;
        RECT 177.820 85.060 178.110 85.105 ;
        RECT 179.185 85.045 179.505 85.105 ;
        RECT 190.225 85.045 190.545 85.105 ;
        RECT 192.985 85.045 193.305 85.305 ;
        RECT 206.415 85.290 206.555 85.445 ;
        RECT 209.175 85.305 209.315 85.785 ;
        RECT 209.560 85.740 209.850 85.785 ;
        RECT 210.095 85.585 210.235 86.125 ;
        RECT 225.200 86.125 227.805 86.265 ;
        RECT 225.200 86.080 225.490 86.125 ;
        RECT 227.485 86.065 227.805 86.125 ;
        RECT 235.855 86.125 237.925 86.265 ;
        RECT 210.480 85.925 210.770 85.970 ;
        RECT 220.125 85.925 220.445 85.985 ;
        RECT 210.480 85.785 220.445 85.925 ;
        RECT 210.480 85.740 210.770 85.785 ;
        RECT 220.125 85.725 220.445 85.785 ;
        RECT 221.980 85.915 222.270 85.970 ;
        RECT 223.345 85.925 223.665 85.985 ;
        RECT 222.515 85.915 223.665 85.925 ;
        RECT 221.980 85.785 223.665 85.915 ;
        RECT 221.980 85.775 222.655 85.785 ;
        RECT 221.980 85.740 222.270 85.775 ;
        RECT 223.345 85.725 223.665 85.785 ;
        RECT 224.740 85.925 225.030 85.970 ;
        RECT 228.405 85.925 228.725 85.985 ;
        RECT 234.400 85.925 234.690 85.970 ;
        RECT 235.305 85.925 235.625 85.985 ;
        RECT 235.855 85.970 235.995 86.125 ;
        RECT 237.605 86.065 237.925 86.125 ;
        RECT 224.740 85.785 228.725 85.925 ;
        RECT 224.740 85.740 225.030 85.785 ;
        RECT 228.405 85.725 228.725 85.785 ;
        RECT 228.955 85.785 235.625 85.925 ;
        RECT 211.400 85.585 211.690 85.630 ;
        RECT 224.265 85.585 224.585 85.645 ;
        RECT 210.095 85.445 224.585 85.585 ;
        RECT 211.400 85.400 211.690 85.445 ;
        RECT 224.265 85.385 224.585 85.445 ;
        RECT 206.340 85.060 206.630 85.290 ;
        RECT 209.085 85.045 209.405 85.305 ;
        RECT 215.065 85.245 215.385 85.305 ;
        RECT 228.955 85.245 229.095 85.785 ;
        RECT 234.400 85.740 234.690 85.785 ;
        RECT 235.305 85.725 235.625 85.785 ;
        RECT 235.780 85.740 236.070 85.970 ;
        RECT 239.465 85.645 239.755 85.860 ;
        RECT 230.705 85.585 231.025 85.645 ;
        RECT 230.705 85.445 239.215 85.585 ;
        RECT 230.705 85.385 231.025 85.445 ;
        RECT 215.065 85.105 229.095 85.245 ;
        RECT 233.465 85.245 233.785 85.305 ;
        RECT 238.065 85.245 238.385 85.305 ;
        RECT 233.465 85.105 238.385 85.245 ;
        RECT 239.075 85.245 239.215 85.445 ;
        RECT 239.445 85.385 239.765 85.645 ;
        RECT 239.995 85.630 240.135 86.465 ;
        RECT 240.455 85.645 240.595 86.805 ;
        RECT 244.505 86.745 244.825 86.805 ;
        RECT 256.465 86.945 256.785 87.005 ;
        RECT 262.445 86.945 262.765 87.005 ;
        RECT 256.465 86.805 262.765 86.945 ;
        RECT 256.465 86.745 256.785 86.805 ;
        RECT 262.445 86.745 262.765 86.805 ;
        RECT 278.085 86.945 278.405 87.005 ;
        RECT 279.020 86.945 279.310 86.990 ;
        RECT 278.085 86.805 279.310 86.945 ;
        RECT 278.085 86.745 278.405 86.805 ;
        RECT 279.020 86.760 279.310 86.805 ;
        RECT 280.860 86.945 281.150 86.990 ;
        RECT 282.685 86.945 283.005 87.005 ;
        RECT 284.985 86.945 285.305 87.005 ;
        RECT 286.825 86.945 287.145 87.005 ;
        RECT 280.860 86.805 283.005 86.945 ;
        RECT 280.860 86.760 281.150 86.805 ;
        RECT 282.685 86.745 283.005 86.805 ;
        RECT 283.235 86.805 287.145 86.945 ;
        RECT 240.825 86.605 241.145 86.665 ;
        RECT 250.025 86.605 250.345 86.665 ;
        RECT 262.905 86.605 263.225 86.665 ;
        RECT 240.825 86.465 263.225 86.605 ;
        RECT 240.825 86.405 241.145 86.465 ;
        RECT 250.025 86.405 250.345 86.465 ;
        RECT 241.760 86.265 242.050 86.310 ;
        RECT 245.425 86.265 245.745 86.325 ;
        RECT 241.760 86.125 245.745 86.265 ;
        RECT 241.760 86.080 242.050 86.125 ;
        RECT 245.425 86.065 245.745 86.125 ;
        RECT 242.665 85.925 242.985 85.985 ;
        RECT 243.140 85.925 243.430 85.970 ;
        RECT 253.705 85.925 254.025 85.985 ;
        RECT 256.925 85.970 257.245 85.985 ;
        RECT 255.970 85.925 256.260 85.970 ;
        RECT 242.665 85.785 243.430 85.925 ;
        RECT 242.665 85.725 242.985 85.785 ;
        RECT 243.140 85.740 243.430 85.785 ;
        RECT 243.675 85.785 254.025 85.925 ;
        RECT 239.920 85.400 240.210 85.630 ;
        RECT 240.365 85.385 240.685 85.645 ;
        RECT 240.970 85.400 241.260 85.630 ;
        RECT 242.220 85.585 242.510 85.630 ;
        RECT 243.675 85.585 243.815 85.785 ;
        RECT 253.705 85.725 254.025 85.785 ;
        RECT 255.175 85.785 256.260 85.925 ;
        RECT 242.220 85.445 243.815 85.585 ;
        RECT 244.505 85.585 244.825 85.645 ;
        RECT 253.245 85.585 253.565 85.645 ;
        RECT 255.175 85.585 255.315 85.785 ;
        RECT 255.970 85.740 256.260 85.785 ;
        RECT 256.685 85.740 257.245 85.970 ;
        RECT 257.400 85.740 257.690 85.970 ;
        RECT 256.925 85.725 257.245 85.740 ;
        RECT 244.505 85.445 253.015 85.585 ;
        RECT 242.220 85.400 242.510 85.445 ;
        RECT 241.045 85.245 241.185 85.400 ;
        RECT 244.505 85.385 244.825 85.445 ;
        RECT 252.875 85.305 253.015 85.445 ;
        RECT 253.245 85.445 255.315 85.585 ;
        RECT 253.245 85.385 253.565 85.445 ;
        RECT 242.665 85.245 242.985 85.305 ;
        RECT 239.075 85.105 242.985 85.245 ;
        RECT 215.065 85.045 215.385 85.105 ;
        RECT 233.465 85.045 233.785 85.105 ;
        RECT 238.065 85.045 238.385 85.105 ;
        RECT 242.665 85.045 242.985 85.105 ;
        RECT 244.060 85.245 244.350 85.290 ;
        RECT 245.425 85.245 245.745 85.305 ;
        RECT 244.060 85.105 245.745 85.245 ;
        RECT 244.060 85.060 244.350 85.105 ;
        RECT 245.425 85.045 245.745 85.105 ;
        RECT 252.785 85.045 253.105 85.305 ;
        RECT 255.175 85.245 255.315 85.445 ;
        RECT 256.465 85.245 256.785 85.305 ;
        RECT 255.175 85.105 256.785 85.245 ;
        RECT 256.465 85.045 256.785 85.105 ;
        RECT 256.925 85.245 257.245 85.305 ;
        RECT 257.475 85.245 257.615 85.740 ;
        RECT 257.845 85.725 258.165 85.985 ;
        RECT 258.395 85.925 258.535 86.465 ;
        RECT 262.905 86.405 263.225 86.465 ;
        RECT 263.380 86.605 263.670 86.650 ;
        RECT 263.825 86.605 264.145 86.665 ;
        RECT 266.585 86.605 266.905 86.665 ;
        RECT 263.380 86.465 264.145 86.605 ;
        RECT 263.380 86.420 263.670 86.465 ;
        RECT 263.825 86.405 264.145 86.465 ;
        RECT 265.755 86.465 266.905 86.605 ;
        RECT 258.765 86.265 259.085 86.325 ;
        RECT 265.755 86.310 265.895 86.465 ;
        RECT 266.585 86.405 266.905 86.465 ;
        RECT 283.235 86.310 283.375 86.805 ;
        RECT 284.985 86.745 285.305 86.805 ;
        RECT 286.825 86.745 287.145 86.805 ;
        RECT 288.205 86.945 288.525 87.005 ;
        RECT 291.900 86.945 292.190 86.990 ;
        RECT 293.725 86.945 294.045 87.005 ;
        RECT 299.245 86.945 299.565 87.005 ;
        RECT 288.205 86.805 294.045 86.945 ;
        RECT 288.205 86.745 288.525 86.805 ;
        RECT 291.900 86.760 292.190 86.805 ;
        RECT 293.725 86.745 294.045 86.805 ;
        RECT 296.575 86.805 299.565 86.945 ;
        RECT 284.030 86.605 284.320 86.650 ;
        RECT 285.920 86.605 286.210 86.650 ;
        RECT 289.040 86.605 289.330 86.650 ;
        RECT 284.030 86.465 289.330 86.605 ;
        RECT 284.030 86.420 284.320 86.465 ;
        RECT 285.920 86.420 286.210 86.465 ;
        RECT 289.040 86.420 289.330 86.465 ;
        RECT 294.200 86.605 294.490 86.650 ;
        RECT 294.645 86.605 294.965 86.665 ;
        RECT 294.200 86.465 294.965 86.605 ;
        RECT 294.200 86.420 294.490 86.465 ;
        RECT 294.645 86.405 294.965 86.465 ;
        RECT 261.080 86.265 261.370 86.310 ;
        RECT 258.765 86.125 261.370 86.265 ;
        RECT 258.765 86.065 259.085 86.125 ;
        RECT 261.080 86.080 261.370 86.125 ;
        RECT 261.540 86.265 261.830 86.310 ;
        RECT 265.680 86.265 265.970 86.310 ;
        RECT 261.540 86.125 265.970 86.265 ;
        RECT 261.540 86.080 261.830 86.125 ;
        RECT 265.680 86.080 265.970 86.125 ;
        RECT 279.555 86.125 281.075 86.265 ;
        RECT 259.700 85.925 259.990 85.970 ;
        RECT 258.395 85.785 259.990 85.925 ;
        RECT 259.700 85.740 259.990 85.785 ;
        RECT 260.145 85.925 260.465 85.985 ;
        RECT 260.620 85.925 260.910 85.970 ;
        RECT 260.145 85.785 260.910 85.925 ;
        RECT 260.145 85.725 260.465 85.785 ;
        RECT 260.620 85.740 260.910 85.785 ;
        RECT 262.445 85.725 262.765 85.985 ;
        RECT 262.905 85.925 263.225 85.985 ;
        RECT 263.840 85.925 264.130 85.970 ;
        RECT 262.905 85.785 264.130 85.925 ;
        RECT 262.905 85.725 263.225 85.785 ;
        RECT 263.840 85.740 264.130 85.785 ;
        RECT 264.285 85.925 264.605 85.985 ;
        RECT 264.760 85.925 265.050 85.970 ;
        RECT 264.285 85.785 265.050 85.925 ;
        RECT 264.285 85.725 264.605 85.785 ;
        RECT 264.760 85.740 265.050 85.785 ;
        RECT 265.220 85.740 265.510 85.970 ;
        RECT 266.125 85.925 266.445 85.985 ;
        RECT 266.600 85.925 266.890 85.970 ;
        RECT 266.125 85.785 266.890 85.925 ;
        RECT 258.780 85.585 259.070 85.630 ;
        RECT 265.295 85.585 265.435 85.740 ;
        RECT 266.125 85.725 266.445 85.785 ;
        RECT 266.600 85.740 266.890 85.785 ;
        RECT 267.980 85.740 268.270 85.970 ;
        RECT 268.425 85.925 268.745 85.985 ;
        RECT 268.900 85.925 269.190 85.970 ;
        RECT 268.425 85.785 269.190 85.925 ;
        RECT 268.055 85.585 268.195 85.740 ;
        RECT 268.425 85.725 268.745 85.785 ;
        RECT 268.900 85.740 269.190 85.785 ;
        RECT 269.345 85.725 269.665 85.985 ;
        RECT 269.805 85.725 270.125 85.985 ;
        RECT 271.185 85.925 271.505 85.985 ;
        RECT 278.085 85.925 278.405 85.985 ;
        RECT 278.560 85.925 278.850 85.970 ;
        RECT 271.185 85.785 278.850 85.925 ;
        RECT 271.185 85.725 271.505 85.785 ;
        RECT 278.085 85.725 278.405 85.785 ;
        RECT 278.560 85.740 278.850 85.785 ;
        RECT 279.555 85.585 279.695 86.125 ;
        RECT 279.940 85.740 280.230 85.970 ;
        RECT 258.780 85.445 265.435 85.585 ;
        RECT 266.215 85.445 268.195 85.585 ;
        RECT 272.195 85.445 279.695 85.585 ;
        RECT 258.780 85.400 259.070 85.445 ;
        RECT 266.215 85.305 266.355 85.445 ;
        RECT 272.195 85.305 272.335 85.445 ;
        RECT 261.525 85.245 261.845 85.305 ;
        RECT 256.925 85.105 261.845 85.245 ;
        RECT 256.925 85.045 257.245 85.105 ;
        RECT 261.525 85.045 261.845 85.105 ;
        RECT 266.125 85.045 266.445 85.305 ;
        RECT 267.505 85.045 267.825 85.305 ;
        RECT 267.965 85.245 268.285 85.305 ;
        RECT 271.200 85.245 271.490 85.290 ;
        RECT 267.965 85.105 271.490 85.245 ;
        RECT 267.965 85.045 268.285 85.105 ;
        RECT 271.200 85.060 271.490 85.105 ;
        RECT 272.105 85.045 272.425 85.305 ;
        RECT 276.705 85.245 277.025 85.305 ;
        RECT 279.005 85.245 279.325 85.305 ;
        RECT 280.015 85.245 280.155 85.740 ;
        RECT 276.705 85.105 280.155 85.245 ;
        RECT 280.935 85.245 281.075 86.125 ;
        RECT 283.160 86.080 283.450 86.310 ;
        RECT 284.525 86.065 284.845 86.325 ;
        RECT 286.365 86.265 286.685 86.325 ;
        RECT 286.365 86.125 295.335 86.265 ;
        RECT 286.365 86.065 286.685 86.125 ;
        RECT 283.625 85.925 283.915 85.970 ;
        RECT 285.460 85.925 285.750 85.970 ;
        RECT 289.040 85.925 289.330 85.970 ;
        RECT 283.625 85.785 289.330 85.925 ;
        RECT 283.625 85.740 283.915 85.785 ;
        RECT 285.460 85.740 285.750 85.785 ;
        RECT 289.040 85.740 289.330 85.785 ;
        RECT 290.120 85.630 290.410 85.945 ;
        RECT 293.265 85.725 293.585 85.985 ;
        RECT 295.195 85.925 295.335 86.125 ;
        RECT 295.565 86.065 295.885 86.325 ;
        RECT 296.575 86.310 296.715 86.805 ;
        RECT 299.245 86.745 299.565 86.805 ;
        RECT 300.180 86.945 300.470 86.990 ;
        RECT 302.005 86.945 302.325 87.005 ;
        RECT 300.180 86.805 302.325 86.945 ;
        RECT 300.180 86.760 300.470 86.805 ;
        RECT 302.005 86.745 302.325 86.805 ;
        RECT 298.800 86.420 299.090 86.650 ;
        RECT 296.500 86.080 296.790 86.310 ;
        RECT 296.945 85.925 297.265 85.985 ;
        RECT 295.195 85.785 297.265 85.925 ;
        RECT 298.875 85.925 299.015 86.420 ;
        RECT 310.745 86.265 311.065 86.325 ;
        RECT 309.455 86.125 311.065 86.265 ;
        RECT 309.455 85.970 309.595 86.125 ;
        RECT 310.745 86.065 311.065 86.125 ;
        RECT 299.260 85.925 299.550 85.970 ;
        RECT 298.875 85.785 299.550 85.925 ;
        RECT 296.945 85.725 297.265 85.785 ;
        RECT 299.260 85.740 299.550 85.785 ;
        RECT 309.380 85.740 309.670 85.970 ;
        RECT 286.820 85.585 287.470 85.630 ;
        RECT 290.120 85.585 290.710 85.630 ;
        RECT 292.345 85.585 292.665 85.645 ;
        RECT 295.105 85.585 295.425 85.645 ;
        RECT 286.820 85.445 295.425 85.585 ;
        RECT 286.820 85.400 287.470 85.445 ;
        RECT 290.420 85.400 290.710 85.445 ;
        RECT 292.345 85.385 292.665 85.445 ;
        RECT 295.105 85.385 295.425 85.445 ;
        RECT 296.025 85.585 296.345 85.645 ;
        RECT 303.845 85.585 304.165 85.645 ;
        RECT 296.025 85.445 304.165 85.585 ;
        RECT 296.025 85.385 296.345 85.445 ;
        RECT 303.845 85.385 304.165 85.445 ;
        RECT 297.405 85.245 297.725 85.305 ;
        RECT 305.685 85.245 306.005 85.305 ;
        RECT 280.935 85.105 306.005 85.245 ;
        RECT 276.705 85.045 277.025 85.105 ;
        RECT 279.005 85.045 279.325 85.105 ;
        RECT 297.405 85.045 297.725 85.105 ;
        RECT 305.685 85.045 306.005 85.105 ;
        RECT 306.145 85.245 306.465 85.305 ;
        RECT 308.460 85.245 308.750 85.290 ;
        RECT 306.145 85.105 308.750 85.245 ;
        RECT 306.145 85.045 306.465 85.105 ;
        RECT 308.460 85.060 308.750 85.105 ;
        RECT 162.095 84.425 311.935 84.905 ;
        RECT 178.265 84.225 178.585 84.285 ;
        RECT 178.740 84.225 179.030 84.270 ;
        RECT 186.545 84.225 186.865 84.285 ;
        RECT 178.265 84.085 186.865 84.225 ;
        RECT 178.265 84.025 178.585 84.085 ;
        RECT 178.740 84.040 179.030 84.085 ;
        RECT 186.545 84.025 186.865 84.085 ;
        RECT 194.825 84.225 195.145 84.285 ;
        RECT 207.720 84.225 208.010 84.270 ;
        RECT 194.825 84.085 208.010 84.225 ;
        RECT 194.825 84.025 195.145 84.085 ;
        RECT 207.720 84.040 208.010 84.085 ;
        RECT 180.220 83.885 180.510 83.930 ;
        RECT 182.865 83.885 183.185 83.945 ;
        RECT 183.460 83.885 184.110 83.930 ;
        RECT 180.220 83.745 184.110 83.885 ;
        RECT 180.220 83.700 180.810 83.745 ;
        RECT 180.520 83.385 180.810 83.700 ;
        RECT 182.865 83.685 183.185 83.745 ;
        RECT 183.460 83.700 184.110 83.745 ;
        RECT 186.100 83.885 186.390 83.930 ;
        RECT 188.385 83.885 188.705 83.945 ;
        RECT 186.100 83.745 188.705 83.885 ;
        RECT 186.100 83.700 186.390 83.745 ;
        RECT 188.385 83.685 188.705 83.745 ;
        RECT 200.805 83.885 201.125 83.945 ;
        RECT 205.420 83.885 205.710 83.930 ;
        RECT 200.805 83.745 205.710 83.885 ;
        RECT 207.795 83.885 207.935 84.040 ;
        RECT 210.925 84.025 211.245 84.285 ;
        RECT 211.845 84.025 212.165 84.285 ;
        RECT 222.425 84.225 222.745 84.285 ;
        RECT 232.545 84.225 232.865 84.285 ;
        RECT 222.425 84.085 232.865 84.225 ;
        RECT 222.425 84.025 222.745 84.085 ;
        RECT 232.545 84.025 232.865 84.085 ;
        RECT 234.845 84.225 235.165 84.285 ;
        RECT 239.445 84.225 239.765 84.285 ;
        RECT 245.440 84.225 245.730 84.270 ;
        RECT 248.645 84.225 248.965 84.285 ;
        RECT 234.845 84.085 244.760 84.225 ;
        RECT 234.845 84.025 235.165 84.085 ;
        RECT 239.445 84.025 239.765 84.085 ;
        RECT 211.935 83.885 212.075 84.025 ;
        RECT 227.025 83.885 227.345 83.945 ;
        RECT 207.795 83.745 212.075 83.885 ;
        RECT 223.435 83.745 227.345 83.885 ;
        RECT 200.805 83.685 201.125 83.745 ;
        RECT 205.420 83.700 205.710 83.745 ;
        RECT 223.435 83.605 223.575 83.745 ;
        RECT 227.025 83.685 227.345 83.745 ;
        RECT 227.960 83.700 228.250 83.930 ;
        RECT 232.635 83.885 232.775 84.025 ;
        RECT 238.985 83.885 239.305 83.945 ;
        RECT 232.635 83.745 239.305 83.885 ;
        RECT 181.600 83.545 181.890 83.590 ;
        RECT 185.180 83.545 185.470 83.590 ;
        RECT 187.015 83.545 187.305 83.590 ;
        RECT 181.600 83.405 187.305 83.545 ;
        RECT 181.600 83.360 181.890 83.405 ;
        RECT 185.180 83.360 185.470 83.405 ;
        RECT 187.015 83.360 187.305 83.405 ;
        RECT 187.480 83.545 187.770 83.590 ;
        RECT 188.845 83.545 189.165 83.605 ;
        RECT 187.480 83.405 189.165 83.545 ;
        RECT 187.480 83.360 187.770 83.405 ;
        RECT 188.845 83.345 189.165 83.405 ;
        RECT 190.240 83.360 190.530 83.590 ;
        RECT 193.445 83.545 193.765 83.605 ;
        RECT 196.220 83.545 196.510 83.590 ;
        RECT 201.740 83.545 202.030 83.590 ;
        RECT 193.445 83.405 202.030 83.545 ;
        RECT 181.600 82.865 181.890 82.910 ;
        RECT 184.720 82.865 185.010 82.910 ;
        RECT 186.610 82.865 186.900 82.910 ;
        RECT 181.600 82.725 186.900 82.865 ;
        RECT 190.315 82.865 190.455 83.360 ;
        RECT 193.445 83.345 193.765 83.405 ;
        RECT 196.220 83.360 196.510 83.405 ;
        RECT 201.740 83.360 202.030 83.405 ;
        RECT 208.640 83.545 208.930 83.590 ;
        RECT 209.085 83.545 209.405 83.605 ;
        RECT 211.860 83.545 212.150 83.590 ;
        RECT 208.640 83.405 213.455 83.545 ;
        RECT 208.640 83.360 208.930 83.405 ;
        RECT 209.085 83.345 209.405 83.405 ;
        RECT 211.860 83.360 212.150 83.405 ;
        RECT 213.315 83.265 213.455 83.405 ;
        RECT 220.140 83.360 220.430 83.590 ;
        RECT 222.440 83.545 222.730 83.590 ;
        RECT 223.345 83.545 223.665 83.605 ;
        RECT 222.440 83.405 223.665 83.545 ;
        RECT 222.440 83.360 222.730 83.405 ;
        RECT 192.540 83.205 192.830 83.250 ;
        RECT 193.905 83.205 194.225 83.265 ;
        RECT 192.540 83.065 194.225 83.205 ;
        RECT 192.540 83.020 192.830 83.065 ;
        RECT 193.905 83.005 194.225 83.065 ;
        RECT 209.560 83.020 209.850 83.250 ;
        RECT 194.365 82.865 194.685 82.925 ;
        RECT 190.315 82.725 194.685 82.865 ;
        RECT 209.635 82.865 209.775 83.020 ;
        RECT 212.765 83.005 213.085 83.265 ;
        RECT 213.225 83.005 213.545 83.265 ;
        RECT 220.215 83.205 220.355 83.360 ;
        RECT 223.345 83.345 223.665 83.405 ;
        RECT 223.805 83.545 224.125 83.605 ;
        RECT 228.035 83.545 228.175 83.700 ;
        RECT 238.985 83.685 239.305 83.745 ;
        RECT 243.600 83.700 243.890 83.930 ;
        RECT 223.805 83.405 228.175 83.545 ;
        RECT 223.805 83.345 224.125 83.405 ;
        RECT 226.580 83.205 226.870 83.250 ;
        RECT 227.025 83.205 227.345 83.265 ;
        RECT 220.215 83.065 222.655 83.205 ;
        RECT 216.445 82.865 216.765 82.925 ;
        RECT 209.635 82.725 216.765 82.865 ;
        RECT 181.600 82.680 181.890 82.725 ;
        RECT 184.720 82.680 185.010 82.725 ;
        RECT 186.610 82.680 186.900 82.725 ;
        RECT 194.365 82.665 194.685 82.725 ;
        RECT 216.445 82.665 216.765 82.725 ;
        RECT 222.515 82.585 222.655 83.065 ;
        RECT 226.580 83.065 227.345 83.205 ;
        RECT 228.035 83.205 228.175 83.405 ;
        RECT 230.245 83.545 230.565 83.605 ;
        RECT 233.005 83.545 233.325 83.605 ;
        RECT 230.245 83.405 233.325 83.545 ;
        RECT 230.245 83.345 230.565 83.405 ;
        RECT 233.005 83.345 233.325 83.405 ;
        RECT 233.925 83.545 234.245 83.605 ;
        RECT 240.825 83.545 241.145 83.605 ;
        RECT 242.220 83.545 242.510 83.590 ;
        RECT 233.925 83.405 242.510 83.545 ;
        RECT 233.925 83.345 234.245 83.405 ;
        RECT 240.825 83.345 241.145 83.405 ;
        RECT 242.220 83.360 242.510 83.405 ;
        RECT 242.960 83.360 243.250 83.590 ;
        RECT 234.385 83.205 234.705 83.265 ;
        RECT 241.745 83.205 242.065 83.265 ;
        RECT 228.035 83.065 231.855 83.205 ;
        RECT 226.580 83.020 226.870 83.065 ;
        RECT 227.025 83.005 227.345 83.065 ;
        RECT 225.185 82.865 225.505 82.925 ;
        RECT 228.880 82.865 229.170 82.910 ;
        RECT 230.705 82.865 231.025 82.925 ;
        RECT 225.185 82.725 231.025 82.865 ;
        RECT 225.185 82.665 225.505 82.725 ;
        RECT 228.880 82.680 229.170 82.725 ;
        RECT 230.705 82.665 231.025 82.725 ;
        RECT 189.305 82.325 189.625 82.585 ;
        RECT 222.425 82.525 222.745 82.585 ;
        RECT 227.485 82.525 227.805 82.585 ;
        RECT 231.715 82.570 231.855 83.065 ;
        RECT 234.385 83.065 242.065 83.205 ;
        RECT 234.385 83.005 234.705 83.065 ;
        RECT 241.745 83.005 242.065 83.065 ;
        RECT 236.685 82.865 237.005 82.925 ;
        RECT 243.035 82.865 243.175 83.360 ;
        RECT 243.675 83.205 243.815 83.700 ;
        RECT 244.045 83.685 244.365 83.945 ;
        RECT 244.620 83.590 244.760 84.085 ;
        RECT 245.440 84.085 248.965 84.225 ;
        RECT 245.440 84.040 245.730 84.085 ;
        RECT 248.645 84.025 248.965 84.085 ;
        RECT 258.305 84.225 258.625 84.285 ;
        RECT 260.145 84.225 260.465 84.285 ;
        RECT 266.125 84.225 266.445 84.285 ;
        RECT 258.305 84.085 260.465 84.225 ;
        RECT 258.305 84.025 258.625 84.085 ;
        RECT 260.145 84.025 260.465 84.085 ;
        RECT 262.075 84.085 266.445 84.225 ;
        RECT 248.185 83.685 248.505 83.945 ;
        RECT 258.395 83.885 258.535 84.025 ;
        RECT 248.735 83.745 258.535 83.885 ;
        RECT 244.545 83.360 244.835 83.590 ;
        RECT 245.425 83.545 245.745 83.605 ;
        RECT 246.820 83.545 247.110 83.590 ;
        RECT 245.425 83.405 247.110 83.545 ;
        RECT 244.045 83.205 244.365 83.265 ;
        RECT 243.675 83.065 244.365 83.205 ;
        RECT 244.620 83.205 244.760 83.360 ;
        RECT 245.425 83.345 245.745 83.405 ;
        RECT 246.820 83.360 247.110 83.405 ;
        RECT 247.265 83.345 247.585 83.605 ;
        RECT 247.740 83.545 248.030 83.590 ;
        RECT 248.275 83.545 248.415 83.685 ;
        RECT 247.740 83.405 248.415 83.545 ;
        RECT 247.740 83.360 248.030 83.405 ;
        RECT 244.620 83.065 247.955 83.205 ;
        RECT 244.045 83.005 244.365 83.065 ;
        RECT 247.815 82.865 247.955 83.065 ;
        RECT 248.185 83.005 248.505 83.265 ;
        RECT 248.735 82.865 248.875 83.745 ;
        RECT 251.405 83.545 251.725 83.605 ;
        RECT 262.075 83.545 262.215 84.085 ;
        RECT 266.125 84.025 266.445 84.085 ;
        RECT 277.625 84.225 277.945 84.285 ;
        RECT 293.265 84.225 293.585 84.285 ;
        RECT 295.580 84.225 295.870 84.270 ;
        RECT 277.625 84.085 282.455 84.225 ;
        RECT 277.625 84.025 277.945 84.085 ;
        RECT 282.315 83.945 282.455 84.085 ;
        RECT 293.265 84.085 295.870 84.225 ;
        RECT 293.265 84.025 293.585 84.085 ;
        RECT 295.580 84.040 295.870 84.085 ;
        RECT 300.625 84.025 300.945 84.285 ;
        RECT 262.445 83.885 262.765 83.945 ;
        RECT 277.165 83.930 277.485 83.945 ;
        RECT 266.600 83.885 266.890 83.930 ;
        RECT 262.445 83.745 266.890 83.885 ;
        RECT 262.445 83.685 262.765 83.745 ;
        RECT 266.600 83.700 266.890 83.745 ;
        RECT 276.700 83.885 277.485 83.930 ;
        RECT 280.300 83.885 280.590 83.930 ;
        RECT 276.700 83.745 280.590 83.885 ;
        RECT 276.700 83.700 277.485 83.745 ;
        RECT 277.165 83.685 277.485 83.700 ;
        RECT 280.000 83.700 280.590 83.745 ;
        RECT 262.920 83.545 263.210 83.590 ;
        RECT 251.405 83.405 263.210 83.545 ;
        RECT 251.405 83.345 251.725 83.405 ;
        RECT 262.920 83.360 263.210 83.405 ;
        RECT 263.380 83.545 263.670 83.590 ;
        RECT 265.205 83.545 265.525 83.605 ;
        RECT 263.380 83.405 265.525 83.545 ;
        RECT 263.380 83.360 263.670 83.405 ;
        RECT 265.205 83.345 265.525 83.405 ;
        RECT 265.665 83.345 265.985 83.605 ;
        RECT 273.505 83.545 273.795 83.590 ;
        RECT 275.340 83.545 275.630 83.590 ;
        RECT 278.920 83.545 279.210 83.590 ;
        RECT 273.505 83.405 279.210 83.545 ;
        RECT 273.505 83.360 273.795 83.405 ;
        RECT 275.340 83.360 275.630 83.405 ;
        RECT 278.920 83.360 279.210 83.405 ;
        RECT 280.000 83.385 280.290 83.700 ;
        RECT 282.225 83.685 282.545 83.945 ;
        RECT 292.345 83.685 292.665 83.945 ;
        RECT 294.200 83.885 294.490 83.930 ;
        RECT 296.025 83.885 296.345 83.945 ;
        RECT 294.200 83.745 296.345 83.885 ;
        RECT 294.200 83.700 294.490 83.745 ;
        RECT 296.025 83.685 296.345 83.745 ;
        RECT 297.405 83.685 297.725 83.945 ;
        RECT 300.715 83.885 300.855 84.025 ;
        RECT 303.385 83.930 303.705 83.945 ;
        RECT 299.795 83.745 300.855 83.885 ;
        RECT 303.380 83.885 304.030 83.930 ;
        RECT 306.980 83.885 307.270 83.930 ;
        RECT 303.380 83.745 307.270 83.885 ;
        RECT 288.205 83.345 288.525 83.605 ;
        RECT 299.795 83.590 299.935 83.745 ;
        RECT 303.380 83.700 304.030 83.745 ;
        RECT 306.680 83.700 307.270 83.745 ;
        RECT 303.385 83.685 303.705 83.700 ;
        RECT 299.720 83.360 300.010 83.590 ;
        RECT 300.185 83.545 300.475 83.590 ;
        RECT 302.020 83.545 302.310 83.590 ;
        RECT 305.600 83.545 305.890 83.590 ;
        RECT 300.185 83.405 305.890 83.545 ;
        RECT 300.185 83.360 300.475 83.405 ;
        RECT 302.020 83.360 302.310 83.405 ;
        RECT 305.600 83.360 305.890 83.405 ;
        RECT 306.680 83.385 306.970 83.700 ;
        RECT 252.785 83.205 253.105 83.265 ;
        RECT 261.065 83.205 261.385 83.265 ;
        RECT 252.785 83.065 261.385 83.205 ;
        RECT 252.785 83.005 253.105 83.065 ;
        RECT 261.065 83.005 261.385 83.065 ;
        RECT 261.525 83.205 261.845 83.265 ;
        RECT 262.460 83.205 262.750 83.250 ;
        RECT 261.525 83.065 262.750 83.205 ;
        RECT 261.525 83.005 261.845 83.065 ;
        RECT 262.460 83.020 262.750 83.065 ;
        RECT 263.840 83.205 264.130 83.250 ;
        RECT 267.520 83.205 267.810 83.250 ;
        RECT 263.840 83.065 267.810 83.205 ;
        RECT 263.840 83.020 264.130 83.065 ;
        RECT 267.520 83.020 267.810 83.065 ;
        RECT 273.040 83.020 273.330 83.250 ;
        RECT 236.685 82.725 244.735 82.865 ;
        RECT 247.815 82.725 248.875 82.865 ;
        RECT 249.105 82.865 249.425 82.925 ;
        RECT 272.105 82.865 272.425 82.925 ;
        RECT 249.105 82.725 272.425 82.865 ;
        RECT 236.685 82.665 237.005 82.725 ;
        RECT 244.595 82.585 244.735 82.725 ;
        RECT 249.105 82.665 249.425 82.725 ;
        RECT 272.105 82.665 272.425 82.725 ;
        RECT 227.960 82.525 228.250 82.570 ;
        RECT 222.425 82.385 228.250 82.525 ;
        RECT 222.425 82.325 222.745 82.385 ;
        RECT 227.485 82.325 227.805 82.385 ;
        RECT 227.960 82.340 228.250 82.385 ;
        RECT 231.640 82.525 231.930 82.570 ;
        RECT 233.925 82.525 234.245 82.585 ;
        RECT 231.640 82.385 234.245 82.525 ;
        RECT 231.640 82.340 231.930 82.385 ;
        RECT 233.925 82.325 234.245 82.385 ;
        RECT 237.145 82.525 237.465 82.585 ;
        RECT 243.125 82.525 243.445 82.585 ;
        RECT 237.145 82.385 243.445 82.525 ;
        RECT 237.145 82.325 237.465 82.385 ;
        RECT 243.125 82.325 243.445 82.385 ;
        RECT 244.505 82.325 244.825 82.585 ;
        RECT 245.885 82.325 246.205 82.585 ;
        RECT 249.565 82.525 249.885 82.585 ;
        RECT 258.305 82.525 258.625 82.585 ;
        RECT 249.565 82.385 258.625 82.525 ;
        RECT 249.565 82.325 249.885 82.385 ;
        RECT 258.305 82.325 258.625 82.385 ;
        RECT 264.745 82.325 265.065 82.585 ;
        RECT 272.565 82.525 272.885 82.585 ;
        RECT 273.115 82.525 273.255 83.020 ;
        RECT 274.405 83.005 274.725 83.265 ;
        RECT 286.380 83.205 286.670 83.250 ;
        RECT 294.645 83.205 294.965 83.265 ;
        RECT 279.555 83.065 294.965 83.205 ;
        RECT 273.910 82.865 274.200 82.910 ;
        RECT 275.800 82.865 276.090 82.910 ;
        RECT 278.920 82.865 279.210 82.910 ;
        RECT 273.910 82.725 279.210 82.865 ;
        RECT 273.910 82.680 274.200 82.725 ;
        RECT 275.800 82.680 276.090 82.725 ;
        RECT 278.920 82.680 279.210 82.725 ;
        RECT 274.865 82.525 275.185 82.585 ;
        RECT 279.555 82.525 279.695 83.065 ;
        RECT 286.380 83.020 286.670 83.065 ;
        RECT 294.645 83.005 294.965 83.065 ;
        RECT 296.945 83.205 297.265 83.265 ;
        RECT 297.880 83.205 298.170 83.250 ;
        RECT 296.945 83.065 298.170 83.205 ;
        RECT 296.945 83.005 297.265 83.065 ;
        RECT 297.880 83.020 298.170 83.065 ;
        RECT 298.325 83.005 298.645 83.265 ;
        RECT 301.085 83.005 301.405 83.265 ;
        RECT 281.765 82.665 282.085 82.925 ;
        RECT 300.590 82.865 300.880 82.910 ;
        RECT 302.480 82.865 302.770 82.910 ;
        RECT 305.600 82.865 305.890 82.910 ;
        RECT 300.590 82.725 305.890 82.865 ;
        RECT 300.590 82.680 300.880 82.725 ;
        RECT 302.480 82.680 302.770 82.725 ;
        RECT 305.600 82.680 305.890 82.725 ;
        RECT 272.565 82.385 279.695 82.525 ;
        RECT 286.825 82.525 287.145 82.585 ;
        RECT 287.300 82.525 287.590 82.570 ;
        RECT 286.825 82.385 287.590 82.525 ;
        RECT 272.565 82.325 272.885 82.385 ;
        RECT 274.865 82.325 275.185 82.385 ;
        RECT 286.825 82.325 287.145 82.385 ;
        RECT 287.300 82.340 287.590 82.385 ;
        RECT 301.545 82.525 301.865 82.585 ;
        RECT 307.985 82.525 308.305 82.585 ;
        RECT 308.460 82.525 308.750 82.570 ;
        RECT 301.545 82.385 308.750 82.525 ;
        RECT 301.545 82.325 301.865 82.385 ;
        RECT 307.985 82.325 308.305 82.385 ;
        RECT 308.460 82.340 308.750 82.385 ;
        RECT 162.095 81.705 311.135 82.185 ;
        RECT 188.335 81.505 188.625 81.550 ;
        RECT 189.305 81.505 189.625 81.565 ;
        RECT 188.335 81.365 189.625 81.505 ;
        RECT 188.335 81.320 188.625 81.365 ;
        RECT 189.305 81.305 189.625 81.365 ;
        RECT 195.285 81.505 195.605 81.565 ;
        RECT 195.760 81.505 196.050 81.550 ;
        RECT 195.285 81.365 196.050 81.505 ;
        RECT 195.285 81.305 195.605 81.365 ;
        RECT 195.760 81.320 196.050 81.365 ;
        RECT 208.180 81.505 208.470 81.550 ;
        RECT 210.465 81.505 210.785 81.565 ;
        RECT 208.180 81.365 210.785 81.505 ;
        RECT 208.180 81.320 208.470 81.365 ;
        RECT 174.125 81.165 174.445 81.225 ;
        RECT 170.535 81.025 174.445 81.165 ;
        RECT 170.535 80.530 170.675 81.025 ;
        RECT 174.125 80.965 174.445 81.025 ;
        RECT 175.520 80.980 175.810 81.210 ;
        RECT 187.890 81.165 188.180 81.210 ;
        RECT 189.780 81.165 190.070 81.210 ;
        RECT 192.900 81.165 193.190 81.210 ;
        RECT 187.890 81.025 193.190 81.165 ;
        RECT 187.890 80.980 188.180 81.025 ;
        RECT 189.780 80.980 190.070 81.025 ;
        RECT 192.900 80.980 193.190 81.025 ;
        RECT 175.595 80.825 175.735 80.980 ;
        RECT 193.905 80.965 194.225 81.225 ;
        RECT 195.835 81.165 195.975 81.320 ;
        RECT 210.465 81.305 210.785 81.365 ;
        RECT 215.525 81.505 215.845 81.565 ;
        RECT 237.145 81.505 237.465 81.565 ;
        RECT 215.525 81.365 238.420 81.505 ;
        RECT 215.525 81.305 215.845 81.365 ;
        RECT 237.145 81.305 237.465 81.365 ;
        RECT 230.705 81.165 231.025 81.225 ;
        RECT 233.465 81.165 233.785 81.225 ;
        RECT 195.835 81.025 228.635 81.165 ;
        RECT 171.915 80.685 175.735 80.825 ;
        RECT 171.915 80.530 172.055 80.685 ;
        RECT 178.725 80.625 179.045 80.885 ;
        RECT 186.085 80.825 186.405 80.885 ;
        RECT 187.020 80.825 187.310 80.870 ;
        RECT 193.995 80.825 194.135 80.965 ;
        RECT 186.085 80.685 194.135 80.825 ;
        RECT 186.085 80.625 186.405 80.685 ;
        RECT 187.020 80.640 187.310 80.685 ;
        RECT 215.985 80.625 216.305 80.885 ;
        RECT 219.680 80.825 219.970 80.870 ;
        RECT 223.805 80.825 224.125 80.885 ;
        RECT 219.680 80.685 224.125 80.825 ;
        RECT 219.680 80.640 219.970 80.685 ;
        RECT 223.805 80.625 224.125 80.685 ;
        RECT 170.460 80.300 170.750 80.530 ;
        RECT 171.840 80.300 172.130 80.530 ;
        RECT 173.205 80.285 173.525 80.545 ;
        RECT 177.345 80.285 177.665 80.545 ;
        RECT 185.640 80.485 185.930 80.530 ;
        RECT 187.485 80.485 187.775 80.530 ;
        RECT 189.320 80.485 189.610 80.530 ;
        RECT 192.900 80.485 193.190 80.530 ;
        RECT 185.640 80.345 187.235 80.485 ;
        RECT 185.640 80.300 185.930 80.345 ;
        RECT 176.425 80.145 176.745 80.205 ;
        RECT 187.095 80.145 187.235 80.345 ;
        RECT 187.485 80.345 193.190 80.485 ;
        RECT 187.485 80.300 187.775 80.345 ;
        RECT 189.320 80.300 189.610 80.345 ;
        RECT 192.900 80.300 193.190 80.345 ;
        RECT 188.845 80.145 189.165 80.205 ;
        RECT 193.980 80.190 194.270 80.505 ;
        RECT 209.100 80.300 209.390 80.530 ;
        RECT 210.020 80.485 210.310 80.530 ;
        RECT 211.845 80.485 212.165 80.545 ;
        RECT 210.020 80.345 212.165 80.485 ;
        RECT 216.075 80.485 216.215 80.625 ;
        RECT 220.125 80.485 220.445 80.545 ;
        RECT 216.075 80.345 220.445 80.485 ;
        RECT 210.020 80.300 210.310 80.345 ;
        RECT 190.680 80.145 191.330 80.190 ;
        RECT 193.980 80.145 194.570 80.190 ;
        RECT 176.425 80.005 178.035 80.145 ;
        RECT 187.095 80.005 189.165 80.145 ;
        RECT 176.425 79.945 176.745 80.005 ;
        RECT 177.895 79.865 178.035 80.005 ;
        RECT 188.845 79.945 189.165 80.005 ;
        RECT 190.315 80.005 194.570 80.145 ;
        RECT 209.175 80.145 209.315 80.300 ;
        RECT 211.845 80.285 212.165 80.345 ;
        RECT 220.125 80.285 220.445 80.345 ;
        RECT 221.980 80.485 222.270 80.530 ;
        RECT 224.725 80.485 225.045 80.545 ;
        RECT 227.485 80.485 227.805 80.545 ;
        RECT 228.495 80.530 228.635 81.025 ;
        RECT 230.705 81.025 233.785 81.165 ;
        RECT 230.705 80.965 231.025 81.025 ;
        RECT 233.465 80.965 233.785 81.025 ;
        RECT 236.685 80.965 237.005 81.225 ;
        RECT 236.775 80.825 236.915 80.965 ;
        RECT 238.280 80.825 238.420 81.365 ;
        RECT 238.985 81.305 239.305 81.565 ;
        RECT 248.185 81.505 248.505 81.565 ;
        RECT 261.525 81.505 261.845 81.565 ;
        RECT 242.295 81.365 261.845 81.505 ;
        RECT 236.775 80.685 237.835 80.825 ;
        RECT 238.280 80.685 238.755 80.825 ;
        RECT 227.960 80.485 228.250 80.530 ;
        RECT 221.980 80.345 223.575 80.485 ;
        RECT 221.980 80.300 222.270 80.345 ;
        RECT 223.435 80.205 223.575 80.345 ;
        RECT 224.725 80.345 228.250 80.485 ;
        RECT 224.725 80.285 225.045 80.345 ;
        RECT 227.485 80.285 227.805 80.345 ;
        RECT 227.960 80.300 228.250 80.345 ;
        RECT 228.420 80.300 228.710 80.530 ;
        RECT 228.880 80.485 229.170 80.530 ;
        RECT 229.325 80.485 229.645 80.545 ;
        RECT 228.880 80.345 229.645 80.485 ;
        RECT 228.880 80.300 229.170 80.345 ;
        RECT 229.325 80.285 229.645 80.345 ;
        RECT 229.800 80.300 230.090 80.530 ;
        RECT 231.625 80.485 231.945 80.545 ;
        RECT 236.700 80.485 236.990 80.530 ;
        RECT 231.625 80.345 236.990 80.485 ;
        RECT 237.695 80.485 237.835 80.685 ;
        RECT 238.615 80.530 238.755 80.685 ;
        RECT 238.080 80.485 238.370 80.530 ;
        RECT 237.695 80.345 238.370 80.485 ;
        RECT 213.225 80.145 213.545 80.205 ;
        RECT 209.175 80.005 213.545 80.145 ;
        RECT 169.525 79.605 169.845 79.865 ;
        RECT 170.905 79.605 171.225 79.865 ;
        RECT 174.140 79.805 174.430 79.850 ;
        RECT 176.885 79.805 177.205 79.865 ;
        RECT 174.140 79.665 177.205 79.805 ;
        RECT 174.140 79.620 174.430 79.665 ;
        RECT 176.885 79.605 177.205 79.665 ;
        RECT 177.805 79.605 178.125 79.865 ;
        RECT 186.560 79.805 186.850 79.850 ;
        RECT 187.925 79.805 188.245 79.865 ;
        RECT 186.560 79.665 188.245 79.805 ;
        RECT 186.560 79.620 186.850 79.665 ;
        RECT 187.925 79.605 188.245 79.665 ;
        RECT 188.385 79.805 188.705 79.865 ;
        RECT 190.315 79.805 190.455 80.005 ;
        RECT 190.680 79.960 191.330 80.005 ;
        RECT 194.280 79.960 194.570 80.005 ;
        RECT 213.225 79.945 213.545 80.005 ;
        RECT 222.425 79.945 222.745 80.205 ;
        RECT 223.345 79.945 223.665 80.205 ;
        RECT 229.875 80.145 230.015 80.300 ;
        RECT 231.625 80.285 231.945 80.345 ;
        RECT 236.700 80.300 236.990 80.345 ;
        RECT 238.080 80.300 238.370 80.345 ;
        RECT 238.540 80.300 238.830 80.530 ;
        RECT 239.075 80.485 239.215 81.305 ;
        RECT 242.295 81.225 242.435 81.365 ;
        RECT 248.185 81.305 248.505 81.365 ;
        RECT 261.525 81.305 261.845 81.365 ;
        RECT 274.405 81.505 274.725 81.565 ;
        RECT 275.340 81.505 275.630 81.550 ;
        RECT 274.405 81.365 275.630 81.505 ;
        RECT 274.405 81.305 274.725 81.365 ;
        RECT 275.340 81.320 275.630 81.365 ;
        RECT 288.205 81.505 288.525 81.565 ;
        RECT 294.660 81.505 294.950 81.550 ;
        RECT 288.205 81.365 294.950 81.505 ;
        RECT 288.205 81.305 288.525 81.365 ;
        RECT 294.660 81.320 294.950 81.365 ;
        RECT 301.085 81.505 301.405 81.565 ;
        RECT 304.320 81.505 304.610 81.550 ;
        RECT 301.085 81.365 304.610 81.505 ;
        RECT 301.085 81.305 301.405 81.365 ;
        RECT 304.320 81.320 304.610 81.365 ;
        RECT 304.765 81.305 305.085 81.565 ;
        RECT 239.905 81.165 240.225 81.225 ;
        RECT 239.905 81.025 241.055 81.165 ;
        RECT 239.905 80.965 240.225 81.025 ;
        RECT 239.445 80.825 239.765 80.885 ;
        RECT 239.445 80.685 240.600 80.825 ;
        RECT 239.445 80.625 239.765 80.685 ;
        RECT 240.460 80.530 240.600 80.685 ;
        RECT 239.920 80.485 240.210 80.530 ;
        RECT 239.075 80.345 240.210 80.485 ;
        RECT 239.920 80.300 240.210 80.345 ;
        RECT 240.385 80.300 240.675 80.530 ;
        RECT 228.495 80.005 230.015 80.145 ;
        RECT 237.620 80.145 237.910 80.190 ;
        RECT 240.915 80.145 241.055 81.025 ;
        RECT 242.205 80.965 242.525 81.225 ;
        RECT 243.585 80.965 243.905 81.225 ;
        RECT 244.045 81.165 244.365 81.225 ;
        RECT 245.425 81.165 245.745 81.225 ;
        RECT 270.265 81.165 270.585 81.225 ;
        RECT 285.870 81.165 286.160 81.210 ;
        RECT 287.760 81.165 288.050 81.210 ;
        RECT 290.880 81.165 291.170 81.210 ;
        RECT 244.045 81.025 283.605 81.165 ;
        RECT 244.045 80.965 244.365 81.025 ;
        RECT 245.425 80.965 245.745 81.025 ;
        RECT 270.265 80.965 270.585 81.025 ;
        RECT 243.675 80.825 243.815 80.965 ;
        RECT 241.835 80.685 243.815 80.825 ;
        RECT 247.725 80.825 248.045 80.885 ;
        RECT 251.405 80.825 251.725 80.885 ;
        RECT 247.725 80.685 251.725 80.825 ;
        RECT 241.835 80.530 241.975 80.685 ;
        RECT 247.725 80.625 248.045 80.685 ;
        RECT 251.405 80.625 251.725 80.685 ;
        RECT 253.705 80.825 254.025 80.885 ;
        RECT 265.665 80.825 265.985 80.885 ;
        RECT 253.705 80.685 265.985 80.825 ;
        RECT 253.705 80.625 254.025 80.685 ;
        RECT 265.665 80.625 265.985 80.685 ;
        RECT 241.760 80.300 242.050 80.530 ;
        RECT 242.450 80.300 242.740 80.530 ;
        RECT 237.620 80.005 241.055 80.145 ;
        RECT 228.495 79.865 228.635 80.005 ;
        RECT 237.620 79.960 237.910 80.005 ;
        RECT 240.455 79.865 240.595 80.005 ;
        RECT 241.285 79.945 241.605 80.205 ;
        RECT 242.525 80.145 242.665 80.300 ;
        RECT 243.585 80.285 243.905 80.545 ;
        RECT 244.505 80.530 244.825 80.545 ;
        RECT 244.340 80.300 244.825 80.530 ;
        RECT 244.505 80.285 244.825 80.300 ;
        RECT 245.425 80.285 245.745 80.545 ;
        RECT 246.345 80.530 246.665 80.545 ;
        RECT 246.130 80.495 246.665 80.530 ;
        RECT 246.130 80.485 247.035 80.495 ;
        RECT 251.865 80.485 252.185 80.545 ;
        RECT 245.910 80.355 252.185 80.485 ;
        RECT 245.910 80.345 246.665 80.355 ;
        RECT 246.895 80.345 252.185 80.355 ;
        RECT 246.130 80.300 246.665 80.345 ;
        RECT 246.345 80.285 246.665 80.300 ;
        RECT 251.865 80.285 252.185 80.345 ;
        RECT 257.845 80.485 258.165 80.545 ;
        RECT 257.845 80.345 258.995 80.485 ;
        RECT 257.845 80.285 258.165 80.345 ;
        RECT 241.835 80.005 242.665 80.145 ;
        RECT 244.980 80.145 245.270 80.190 ;
        RECT 248.185 80.145 248.505 80.205 ;
        RECT 244.980 80.005 248.505 80.145 ;
        RECT 258.855 80.145 258.995 80.345 ;
        RECT 259.225 80.285 259.545 80.545 ;
        RECT 259.700 80.300 259.990 80.530 ;
        RECT 260.160 80.485 260.450 80.530 ;
        RECT 260.605 80.485 260.925 80.545 ;
        RECT 260.160 80.345 260.925 80.485 ;
        RECT 260.160 80.300 260.450 80.345 ;
        RECT 259.775 80.145 259.915 80.300 ;
        RECT 260.605 80.285 260.925 80.345 ;
        RECT 261.080 80.485 261.370 80.530 ;
        RECT 268.425 80.485 268.745 80.545 ;
        RECT 261.080 80.345 268.745 80.485 ;
        RECT 261.080 80.300 261.370 80.345 ;
        RECT 268.425 80.285 268.745 80.345 ;
        RECT 274.880 80.485 275.170 80.530 ;
        RECT 275.325 80.485 275.645 80.545 ;
        RECT 274.880 80.345 275.645 80.485 ;
        RECT 274.880 80.300 275.170 80.345 ;
        RECT 275.325 80.285 275.645 80.345 ;
        RECT 276.260 80.485 276.550 80.530 ;
        RECT 278.545 80.485 278.865 80.545 ;
        RECT 276.260 80.345 278.865 80.485 ;
        RECT 283.465 80.485 283.605 81.025 ;
        RECT 285.870 81.025 291.170 81.165 ;
        RECT 285.870 80.980 286.160 81.025 ;
        RECT 287.760 80.980 288.050 81.025 ;
        RECT 290.880 80.980 291.170 81.025 ;
        RECT 296.025 81.165 296.345 81.225 ;
        RECT 298.800 81.165 299.090 81.210 ;
        RECT 296.025 81.025 299.090 81.165 ;
        RECT 296.025 80.965 296.345 81.025 ;
        RECT 298.800 80.980 299.090 81.025 ;
        RECT 284.985 80.625 285.305 80.885 ;
        RECT 286.380 80.825 286.670 80.870 ;
        RECT 286.825 80.825 287.145 80.885 ;
        RECT 286.380 80.685 287.145 80.825 ;
        RECT 286.380 80.640 286.670 80.685 ;
        RECT 286.825 80.625 287.145 80.685 ;
        RECT 290.045 80.825 290.365 80.885 ;
        RECT 297.420 80.825 297.710 80.870 ;
        RECT 290.045 80.685 297.710 80.825 ;
        RECT 290.045 80.625 290.365 80.685 ;
        RECT 297.420 80.640 297.710 80.685 ;
        RECT 298.325 80.825 298.645 80.885 ;
        RECT 301.560 80.825 301.850 80.870 ;
        RECT 298.325 80.685 301.850 80.825 ;
        RECT 298.325 80.625 298.645 80.685 ;
        RECT 301.560 80.640 301.850 80.685 ;
        RECT 285.465 80.485 285.755 80.530 ;
        RECT 287.300 80.485 287.590 80.530 ;
        RECT 290.880 80.485 291.170 80.530 ;
        RECT 283.465 80.345 285.215 80.485 ;
        RECT 276.260 80.300 276.550 80.345 ;
        RECT 278.545 80.285 278.865 80.345 ;
        RECT 258.855 80.005 259.915 80.145 ;
        RECT 277.165 80.145 277.485 80.205 ;
        RECT 284.525 80.145 284.845 80.205 ;
        RECT 277.165 80.005 284.845 80.145 ;
        RECT 241.835 79.865 241.975 80.005 ;
        RECT 244.980 79.960 245.270 80.005 ;
        RECT 248.185 79.945 248.505 80.005 ;
        RECT 277.165 79.945 277.485 80.005 ;
        RECT 284.525 79.945 284.845 80.005 ;
        RECT 188.385 79.665 190.455 79.805 ;
        RECT 194.825 79.805 195.145 79.865 ;
        RECT 214.145 79.805 214.465 79.865 ;
        RECT 194.825 79.665 214.465 79.805 ;
        RECT 188.385 79.605 188.705 79.665 ;
        RECT 194.825 79.605 195.145 79.665 ;
        RECT 214.145 79.605 214.465 79.665 ;
        RECT 227.025 79.605 227.345 79.865 ;
        RECT 228.405 79.605 228.725 79.865 ;
        RECT 239.445 79.605 239.765 79.865 ;
        RECT 240.365 79.605 240.685 79.865 ;
        RECT 241.745 79.605 242.065 79.865 ;
        RECT 243.125 79.605 243.445 79.865 ;
        RECT 246.805 79.605 247.125 79.865 ;
        RECT 258.320 79.805 258.610 79.850 ;
        RECT 260.605 79.805 260.925 79.865 ;
        RECT 258.320 79.665 260.925 79.805 ;
        RECT 258.320 79.620 258.610 79.665 ;
        RECT 260.605 79.605 260.925 79.665 ;
        RECT 273.960 79.805 274.250 79.850 ;
        RECT 274.865 79.805 275.185 79.865 ;
        RECT 273.960 79.665 275.185 79.805 ;
        RECT 285.075 79.805 285.215 80.345 ;
        RECT 285.465 80.345 291.170 80.485 ;
        RECT 285.465 80.300 285.755 80.345 ;
        RECT 287.300 80.300 287.590 80.345 ;
        RECT 290.880 80.300 291.170 80.345 ;
        RECT 291.960 80.190 292.250 80.505 ;
        RECT 293.725 80.485 294.045 80.545 ;
        RECT 296.945 80.485 297.265 80.545 ;
        RECT 293.725 80.345 297.265 80.485 ;
        RECT 293.725 80.285 294.045 80.345 ;
        RECT 296.945 80.285 297.265 80.345 ;
        RECT 300.640 80.485 300.930 80.530 ;
        RECT 304.305 80.485 304.625 80.545 ;
        RECT 304.855 80.485 304.995 81.305 ;
        RECT 300.640 80.345 304.995 80.485 ;
        RECT 300.640 80.300 300.930 80.345 ;
        RECT 304.305 80.285 304.625 80.345 ;
        RECT 305.225 80.285 305.545 80.545 ;
        RECT 288.660 80.145 289.310 80.190 ;
        RECT 291.960 80.145 292.550 80.190 ;
        RECT 292.805 80.145 293.125 80.205 ;
        RECT 303.385 80.145 303.705 80.205 ;
        RECT 288.660 80.005 303.705 80.145 ;
        RECT 288.660 79.960 289.310 80.005 ;
        RECT 292.260 79.960 292.550 80.005 ;
        RECT 292.805 79.945 293.125 80.005 ;
        RECT 303.385 79.945 303.705 80.005 ;
        RECT 293.740 79.805 294.030 79.850 ;
        RECT 296.500 79.805 296.790 79.850 ;
        RECT 285.075 79.665 296.790 79.805 ;
        RECT 273.960 79.620 274.250 79.665 ;
        RECT 274.865 79.605 275.185 79.665 ;
        RECT 293.740 79.620 294.030 79.665 ;
        RECT 296.500 79.620 296.790 79.665 ;
        RECT 301.085 79.605 301.405 79.865 ;
        RECT 162.095 78.985 311.935 79.465 ;
        RECT 187.005 78.785 187.325 78.845 ;
        RECT 168.235 78.645 187.325 78.785 ;
        RECT 168.235 78.150 168.375 78.645 ;
        RECT 187.005 78.585 187.325 78.645 ;
        RECT 188.845 78.785 189.165 78.845 ;
        RECT 198.060 78.785 198.350 78.830 ;
        RECT 188.845 78.645 198.350 78.785 ;
        RECT 188.845 78.585 189.165 78.645 ;
        RECT 198.060 78.600 198.350 78.645 ;
        RECT 199.900 78.785 200.190 78.830 ;
        RECT 200.805 78.785 201.125 78.845 ;
        RECT 215.985 78.785 216.305 78.845 ;
        RECT 199.900 78.645 216.305 78.785 ;
        RECT 199.900 78.600 200.190 78.645 ;
        RECT 200.805 78.585 201.125 78.645 ;
        RECT 215.985 78.585 216.305 78.645 ;
        RECT 219.665 78.785 219.985 78.845 ;
        RECT 221.505 78.785 221.825 78.845 ;
        RECT 219.665 78.645 221.825 78.785 ;
        RECT 219.665 78.585 219.985 78.645 ;
        RECT 221.505 78.585 221.825 78.645 ;
        RECT 222.425 78.785 222.745 78.845 ;
        RECT 223.345 78.785 223.665 78.845 ;
        RECT 227.040 78.785 227.330 78.830 ;
        RECT 222.425 78.645 223.665 78.785 ;
        RECT 222.425 78.585 222.745 78.645 ;
        RECT 223.345 78.585 223.665 78.645 ;
        RECT 224.815 78.645 227.330 78.785 ;
        RECT 169.540 78.445 169.830 78.490 ;
        RECT 170.905 78.445 171.225 78.505 ;
        RECT 169.540 78.305 171.225 78.445 ;
        RECT 169.540 78.260 169.830 78.305 ;
        RECT 170.905 78.245 171.225 78.305 ;
        RECT 171.820 78.445 172.470 78.490 ;
        RECT 172.745 78.445 173.065 78.505 ;
        RECT 175.420 78.445 175.710 78.490 ;
        RECT 171.820 78.305 175.710 78.445 ;
        RECT 171.820 78.260 172.470 78.305 ;
        RECT 172.745 78.245 173.065 78.305 ;
        RECT 175.120 78.260 175.710 78.305 ;
        RECT 176.885 78.445 177.205 78.505 ;
        RECT 179.200 78.445 179.490 78.490 ;
        RECT 176.885 78.305 179.490 78.445 ;
        RECT 168.160 77.920 168.450 78.150 ;
        RECT 168.625 78.105 168.915 78.150 ;
        RECT 170.460 78.105 170.750 78.150 ;
        RECT 174.040 78.105 174.330 78.150 ;
        RECT 168.625 77.965 174.330 78.105 ;
        RECT 168.625 77.920 168.915 77.965 ;
        RECT 170.460 77.920 170.750 77.965 ;
        RECT 174.040 77.920 174.330 77.965 ;
        RECT 175.120 77.945 175.410 78.260 ;
        RECT 176.885 78.245 177.205 78.305 ;
        RECT 179.200 78.260 179.490 78.305 ;
        RECT 179.645 78.445 179.965 78.505 ;
        RECT 181.480 78.445 182.130 78.490 ;
        RECT 185.080 78.445 185.370 78.490 ;
        RECT 179.645 78.305 185.370 78.445 ;
        RECT 179.645 78.245 179.965 78.305 ;
        RECT 181.480 78.260 182.130 78.305 ;
        RECT 184.780 78.260 185.370 78.305 ;
        RECT 178.285 78.105 178.575 78.150 ;
        RECT 180.120 78.105 180.410 78.150 ;
        RECT 183.700 78.105 183.990 78.150 ;
        RECT 178.285 77.965 183.990 78.105 ;
        RECT 178.285 77.920 178.575 77.965 ;
        RECT 180.120 77.920 180.410 77.965 ;
        RECT 183.700 77.920 183.990 77.965 ;
        RECT 184.780 77.945 185.070 78.260 ;
        RECT 187.095 78.105 187.235 78.585 ;
        RECT 187.925 78.445 188.245 78.505 ;
        RECT 189.780 78.445 190.070 78.490 ;
        RECT 187.925 78.305 190.070 78.445 ;
        RECT 187.925 78.245 188.245 78.305 ;
        RECT 189.780 78.260 190.070 78.305 ;
        RECT 192.060 78.445 192.710 78.490 ;
        RECT 195.660 78.445 195.950 78.490 ;
        RECT 192.060 78.305 195.950 78.445 ;
        RECT 192.060 78.260 192.710 78.305 ;
        RECT 195.360 78.260 195.950 78.305 ;
        RECT 196.665 78.445 196.985 78.505 ;
        RECT 200.360 78.445 200.650 78.490 ;
        RECT 196.665 78.305 200.650 78.445 ;
        RECT 187.465 78.105 187.785 78.165 ;
        RECT 188.400 78.105 188.690 78.150 ;
        RECT 187.095 77.965 188.690 78.105 ;
        RECT 187.465 77.905 187.785 77.965 ;
        RECT 188.400 77.920 188.690 77.965 ;
        RECT 188.865 78.105 189.155 78.150 ;
        RECT 190.700 78.105 190.990 78.150 ;
        RECT 194.280 78.105 194.570 78.150 ;
        RECT 188.865 77.965 194.570 78.105 ;
        RECT 188.865 77.920 189.155 77.965 ;
        RECT 190.700 77.920 190.990 77.965 ;
        RECT 194.280 77.920 194.570 77.965 ;
        RECT 194.825 77.905 195.145 78.165 ;
        RECT 195.360 77.945 195.650 78.260 ;
        RECT 196.665 78.245 196.985 78.305 ;
        RECT 200.360 78.260 200.650 78.305 ;
        RECT 206.325 78.445 206.645 78.505 ;
        RECT 207.260 78.445 207.550 78.490 ;
        RECT 206.325 78.305 207.550 78.445 ;
        RECT 200.435 78.105 200.575 78.260 ;
        RECT 206.325 78.245 206.645 78.305 ;
        RECT 207.260 78.260 207.550 78.305 ;
        RECT 207.720 78.445 208.010 78.490 ;
        RECT 207.720 78.305 224.495 78.445 ;
        RECT 207.720 78.260 208.010 78.305 ;
        RECT 200.435 77.965 206.555 78.105 ;
        RECT 177.805 77.565 178.125 77.825 ;
        RECT 186.560 77.765 186.850 77.810 ;
        RECT 194.915 77.765 195.055 77.905 ;
        RECT 186.560 77.625 195.055 77.765 ;
        RECT 186.560 77.580 186.850 77.625 ;
        RECT 169.030 77.425 169.320 77.470 ;
        RECT 170.920 77.425 171.210 77.470 ;
        RECT 174.040 77.425 174.330 77.470 ;
        RECT 169.030 77.285 174.330 77.425 ;
        RECT 169.030 77.240 169.320 77.285 ;
        RECT 170.920 77.240 171.210 77.285 ;
        RECT 174.040 77.240 174.330 77.285 ;
        RECT 176.425 77.425 176.745 77.485 ;
        RECT 176.900 77.425 177.190 77.470 ;
        RECT 176.425 77.285 177.190 77.425 ;
        RECT 176.425 77.225 176.745 77.285 ;
        RECT 176.900 77.240 177.190 77.285 ;
        RECT 178.690 77.425 178.980 77.470 ;
        RECT 180.580 77.425 180.870 77.470 ;
        RECT 183.700 77.425 183.990 77.470 ;
        RECT 178.690 77.285 183.990 77.425 ;
        RECT 178.690 77.240 178.980 77.285 ;
        RECT 180.580 77.240 180.870 77.285 ;
        RECT 183.700 77.240 183.990 77.285 ;
        RECT 178.265 77.085 178.585 77.145 ;
        RECT 186.635 77.085 186.775 77.580 ;
        RECT 189.270 77.425 189.560 77.470 ;
        RECT 191.160 77.425 191.450 77.470 ;
        RECT 194.280 77.425 194.570 77.470 ;
        RECT 189.270 77.285 194.570 77.425 ;
        RECT 189.270 77.240 189.560 77.285 ;
        RECT 191.160 77.240 191.450 77.285 ;
        RECT 194.280 77.240 194.570 77.285 ;
        RECT 195.375 77.425 195.515 77.945 ;
        RECT 197.125 77.765 197.445 77.825 ;
        RECT 200.820 77.765 201.110 77.810 ;
        RECT 202.185 77.765 202.505 77.825 ;
        RECT 197.125 77.625 202.505 77.765 ;
        RECT 197.125 77.565 197.445 77.625 ;
        RECT 200.820 77.580 201.110 77.625 ;
        RECT 202.185 77.565 202.505 77.625 ;
        RECT 195.375 77.285 200.575 77.425 ;
        RECT 178.265 76.945 186.775 77.085 ;
        RECT 188.385 77.085 188.705 77.145 ;
        RECT 195.375 77.085 195.515 77.285 ;
        RECT 188.385 76.945 195.515 77.085 ;
        RECT 196.665 77.085 196.985 77.145 ;
        RECT 197.140 77.085 197.430 77.130 ;
        RECT 196.665 76.945 197.430 77.085 ;
        RECT 200.435 77.085 200.575 77.285 ;
        RECT 205.865 77.225 206.185 77.485 ;
        RECT 200.805 77.085 201.125 77.145 ;
        RECT 200.435 76.945 201.125 77.085 ;
        RECT 206.415 77.085 206.555 77.965 ;
        RECT 206.785 77.905 207.105 78.165 ;
        RECT 206.875 77.425 207.015 77.905 ;
        RECT 207.335 77.765 207.475 78.260 ;
        RECT 223.435 78.165 223.575 78.305 ;
        RECT 208.625 77.905 208.945 78.165 ;
        RECT 209.545 77.905 209.865 78.165 ;
        RECT 210.005 78.105 210.325 78.165 ;
        RECT 210.480 78.105 210.770 78.150 ;
        RECT 210.005 77.965 210.770 78.105 ;
        RECT 210.005 77.905 210.325 77.965 ;
        RECT 210.480 77.920 210.770 77.965 ;
        RECT 214.145 77.905 214.465 78.165 ;
        RECT 218.745 77.905 219.065 78.165 ;
        RECT 219.665 78.150 219.985 78.165 ;
        RECT 219.500 77.920 219.985 78.150 ;
        RECT 219.665 77.905 219.985 77.920 ;
        RECT 220.125 77.905 220.445 78.165 ;
        RECT 221.045 78.150 221.365 78.165 ;
        RECT 220.600 77.920 220.890 78.150 ;
        RECT 221.045 78.105 221.375 78.150 ;
        RECT 221.045 77.965 221.560 78.105 ;
        RECT 221.045 77.920 221.375 77.965 ;
        RECT 210.925 77.765 211.245 77.825 ;
        RECT 207.335 77.625 211.245 77.765 ;
        RECT 214.235 77.765 214.375 77.905 ;
        RECT 220.675 77.765 220.815 77.920 ;
        RECT 221.045 77.905 221.365 77.920 ;
        RECT 222.885 77.905 223.205 78.165 ;
        RECT 223.345 77.905 223.665 78.165 ;
        RECT 224.355 78.150 224.495 78.305 ;
        RECT 223.820 77.920 224.110 78.150 ;
        RECT 224.285 77.920 224.575 78.150 ;
        RECT 214.235 77.625 220.815 77.765 ;
        RECT 222.975 77.765 223.115 77.905 ;
        RECT 223.895 77.765 224.035 77.920 ;
        RECT 222.975 77.625 224.035 77.765 ;
        RECT 210.925 77.565 211.245 77.625 ;
        RECT 224.815 77.485 224.955 78.645 ;
        RECT 227.040 78.600 227.330 78.645 ;
        RECT 228.880 78.785 229.170 78.830 ;
        RECT 234.845 78.785 235.165 78.845 ;
        RECT 239.905 78.785 240.225 78.845 ;
        RECT 243.140 78.785 243.430 78.830 ;
        RECT 245.425 78.785 245.745 78.845 ;
        RECT 247.265 78.785 247.585 78.845 ;
        RECT 228.880 78.645 235.165 78.785 ;
        RECT 228.880 78.600 229.170 78.645 ;
        RECT 225.185 78.245 225.505 78.505 ;
        RECT 228.955 78.445 229.095 78.600 ;
        RECT 234.845 78.585 235.165 78.645 ;
        RECT 236.775 78.645 239.215 78.785 ;
        RECT 226.425 78.305 229.095 78.445 ;
        RECT 231.625 78.445 231.945 78.505 ;
        RECT 236.775 78.445 236.915 78.645 ;
        RECT 231.625 78.305 236.915 78.445 ;
        RECT 226.425 78.150 226.565 78.305 ;
        RECT 231.625 78.245 231.945 78.305 ;
        RECT 237.145 78.245 237.465 78.505 ;
        RECT 238.205 78.445 238.495 78.490 ;
        RECT 238.205 78.260 238.525 78.445 ;
        RECT 225.660 77.920 225.950 78.150 ;
        RECT 226.350 77.920 226.640 78.150 ;
        RECT 225.735 77.765 225.875 77.920 ;
        RECT 227.945 77.905 228.265 78.165 ;
        RECT 228.880 78.105 229.170 78.150 ;
        RECT 229.785 78.105 230.105 78.165 ;
        RECT 232.545 78.105 232.865 78.165 ;
        RECT 234.845 78.105 235.165 78.165 ;
        RECT 228.880 77.965 232.865 78.105 ;
        RECT 228.880 77.920 229.170 77.965 ;
        RECT 229.785 77.905 230.105 77.965 ;
        RECT 232.545 77.905 232.865 77.965 ;
        RECT 233.095 77.965 235.165 78.105 ;
        RECT 237.235 78.105 237.375 78.245 ;
        RECT 237.620 78.105 237.910 78.150 ;
        RECT 237.235 77.965 237.910 78.105 ;
        RECT 238.385 78.105 238.525 78.260 ;
        RECT 238.385 77.965 238.755 78.105 ;
        RECT 233.095 77.765 233.235 77.965 ;
        RECT 234.845 77.905 235.165 77.965 ;
        RECT 237.620 77.920 237.910 77.965 ;
        RECT 238.615 77.825 238.755 77.965 ;
        RECT 225.735 77.625 233.235 77.765 ;
        RECT 233.925 77.565 234.245 77.825 ;
        RECT 235.305 77.765 235.625 77.825 ;
        RECT 235.780 77.765 236.070 77.810 ;
        RECT 236.685 77.765 237.005 77.825 ;
        RECT 235.305 77.625 237.005 77.765 ;
        RECT 235.305 77.565 235.625 77.625 ;
        RECT 235.780 77.580 236.070 77.625 ;
        RECT 236.685 77.565 237.005 77.625 ;
        RECT 237.160 77.580 237.450 77.810 ;
        RECT 213.685 77.425 214.005 77.485 ;
        RECT 206.875 77.285 214.005 77.425 ;
        RECT 213.685 77.225 214.005 77.285 ;
        RECT 221.980 77.425 222.270 77.470 ;
        RECT 223.345 77.425 223.665 77.485 ;
        RECT 221.980 77.285 223.665 77.425 ;
        RECT 221.980 77.240 222.270 77.285 ;
        RECT 223.345 77.225 223.665 77.285 ;
        RECT 224.725 77.225 225.045 77.485 ;
        RECT 232.085 77.425 232.405 77.485 ;
        RECT 234.015 77.425 234.155 77.565 ;
        RECT 237.235 77.425 237.375 77.580 ;
        RECT 238.525 77.565 238.845 77.825 ;
        RECT 239.075 77.765 239.215 78.645 ;
        RECT 239.905 78.645 241.975 78.785 ;
        RECT 239.905 78.585 240.225 78.645 ;
        RECT 241.835 78.490 241.975 78.645 ;
        RECT 243.140 78.645 245.745 78.785 ;
        RECT 243.140 78.600 243.430 78.645 ;
        RECT 245.425 78.585 245.745 78.645 ;
        RECT 245.975 78.645 247.585 78.785 ;
        RECT 241.760 78.260 242.050 78.490 ;
        RECT 245.975 78.445 246.115 78.645 ;
        RECT 247.265 78.585 247.585 78.645 ;
        RECT 247.725 78.785 248.045 78.845 ;
        RECT 256.005 78.785 256.325 78.845 ;
        RECT 247.725 78.645 256.325 78.785 ;
        RECT 247.725 78.585 248.045 78.645 ;
        RECT 256.005 78.585 256.325 78.645 ;
        RECT 259.685 78.785 260.005 78.845 ;
        RECT 274.865 78.785 275.185 78.845 ;
        RECT 259.685 78.645 260.375 78.785 ;
        RECT 259.685 78.585 260.005 78.645 ;
        RECT 244.595 78.305 246.115 78.445 ;
        RECT 246.345 78.445 246.665 78.505 ;
        RECT 246.345 78.305 247.955 78.445 ;
        RECT 239.905 77.905 240.225 78.165 ;
        RECT 242.665 78.150 242.985 78.165 ;
        RECT 240.385 77.920 240.675 78.150 ;
        RECT 241.300 78.105 241.590 78.150 ;
        RECT 240.915 77.965 241.590 78.105 ;
        RECT 240.460 77.765 240.600 77.920 ;
        RECT 239.075 77.625 240.600 77.765 ;
        RECT 238.065 77.425 238.385 77.485 ;
        RECT 232.085 77.285 236.915 77.425 ;
        RECT 237.235 77.285 238.385 77.425 ;
        RECT 232.085 77.225 232.405 77.285 ;
        RECT 236.225 77.085 236.545 77.145 ;
        RECT 206.415 76.945 236.545 77.085 ;
        RECT 236.775 77.085 236.915 77.285 ;
        RECT 238.065 77.225 238.385 77.285 ;
        RECT 238.985 77.225 239.305 77.485 ;
        RECT 240.915 77.085 241.055 77.965 ;
        RECT 241.300 77.920 241.590 77.965 ;
        RECT 242.440 77.920 242.985 78.150 ;
        RECT 243.600 78.105 243.890 78.150 ;
        RECT 244.045 78.105 244.365 78.165 ;
        RECT 244.595 78.150 244.735 78.305 ;
        RECT 246.345 78.245 246.665 78.305 ;
        RECT 243.600 77.965 244.365 78.105 ;
        RECT 243.600 77.920 243.890 77.965 ;
        RECT 242.665 77.905 242.985 77.920 ;
        RECT 244.045 77.905 244.365 77.965 ;
        RECT 244.520 77.920 244.810 78.150 ;
        RECT 244.980 77.920 245.270 78.150 ;
        RECT 236.775 76.945 241.055 77.085 ;
        RECT 242.205 77.085 242.525 77.145 ;
        RECT 244.505 77.085 244.825 77.145 ;
        RECT 245.055 77.085 245.195 77.920 ;
        RECT 245.425 77.905 245.745 78.165 ;
        RECT 247.815 78.150 247.955 78.305 ;
        RECT 248.645 78.245 248.965 78.505 ;
        RECT 258.305 78.445 258.625 78.505 ;
        RECT 258.305 78.305 258.805 78.445 ;
        RECT 258.305 78.245 258.625 78.305 ;
        RECT 246.820 77.920 247.110 78.150 ;
        RECT 247.740 77.920 248.030 78.150 ;
        RECT 246.895 77.765 247.035 77.920 ;
        RECT 248.735 77.765 248.875 78.245 ;
        RECT 256.465 77.905 256.785 78.165 ;
        RECT 256.945 77.920 257.235 78.150 ;
        RECT 257.385 78.105 257.705 78.165 ;
        RECT 260.235 78.150 260.375 78.645 ;
        RECT 274.035 78.645 275.185 78.785 ;
        RECT 261.065 78.445 261.385 78.505 ;
        RECT 261.540 78.445 261.830 78.490 ;
        RECT 261.065 78.305 261.830 78.445 ;
        RECT 261.065 78.245 261.385 78.305 ;
        RECT 261.540 78.260 261.830 78.305 ;
        RECT 261.985 78.245 262.305 78.505 ;
        RECT 274.035 78.490 274.175 78.645 ;
        RECT 274.865 78.585 275.185 78.645 ;
        RECT 284.525 78.785 284.845 78.845 ;
        RECT 295.105 78.785 295.425 78.845 ;
        RECT 284.525 78.645 291.195 78.785 ;
        RECT 284.525 78.585 284.845 78.645 ;
        RECT 273.960 78.260 274.250 78.490 ;
        RECT 276.240 78.445 276.890 78.490 ;
        RECT 277.165 78.445 277.485 78.505 ;
        RECT 279.840 78.445 280.130 78.490 ;
        RECT 276.240 78.305 280.130 78.445 ;
        RECT 276.240 78.260 276.890 78.305 ;
        RECT 277.165 78.245 277.485 78.305 ;
        RECT 279.540 78.260 280.130 78.305 ;
        RECT 282.225 78.445 282.545 78.505 ;
        RECT 284.985 78.445 285.305 78.505 ;
        RECT 289.600 78.445 289.890 78.490 ;
        RECT 282.225 78.305 283.605 78.445 ;
        RECT 257.860 78.105 258.150 78.150 ;
        RECT 257.385 77.965 258.150 78.105 ;
        RECT 246.895 77.625 248.875 77.765 ;
        RECT 250.485 77.765 250.805 77.825 ;
        RECT 257.015 77.765 257.155 77.920 ;
        RECT 257.385 77.905 257.705 77.965 ;
        RECT 257.860 77.920 258.150 77.965 ;
        RECT 258.805 77.920 259.095 78.150 ;
        RECT 260.160 77.920 260.450 78.150 ;
        RECT 260.625 78.105 260.915 78.150 ;
        RECT 262.485 78.105 262.775 78.150 ;
        RECT 264.285 78.105 264.605 78.165 ;
        RECT 260.625 77.965 262.215 78.105 ;
        RECT 260.625 77.920 260.915 77.965 ;
        RECT 250.485 77.625 257.155 77.765 ;
        RECT 250.485 77.565 250.805 77.625 ;
        RECT 258.855 77.145 258.995 77.920 ;
        RECT 261.065 77.765 261.385 77.825 ;
        RECT 262.075 77.765 262.215 77.965 ;
        RECT 262.485 77.965 264.605 78.105 ;
        RECT 262.485 77.920 262.775 77.965 ;
        RECT 264.285 77.905 264.605 77.965 ;
        RECT 270.265 78.105 270.585 78.165 ;
        RECT 272.565 78.105 272.885 78.165 ;
        RECT 270.265 77.965 272.885 78.105 ;
        RECT 270.265 77.905 270.585 77.965 ;
        RECT 272.565 77.905 272.885 77.965 ;
        RECT 273.045 78.105 273.335 78.150 ;
        RECT 274.880 78.105 275.170 78.150 ;
        RECT 278.460 78.105 278.750 78.150 ;
        RECT 273.045 77.965 278.750 78.105 ;
        RECT 273.045 77.920 273.335 77.965 ;
        RECT 274.880 77.920 275.170 77.965 ;
        RECT 278.460 77.920 278.750 77.965 ;
        RECT 279.540 77.945 279.830 78.260 ;
        RECT 282.225 78.245 282.545 78.305 ;
        RECT 283.465 78.105 283.605 78.305 ;
        RECT 284.985 78.305 289.890 78.445 ;
        RECT 284.985 78.245 285.305 78.305 ;
        RECT 289.600 78.260 289.890 78.305 ;
        RECT 291.055 78.165 291.195 78.645 ;
        RECT 295.105 78.645 296.255 78.785 ;
        RECT 295.105 78.585 295.425 78.645 ;
        RECT 296.115 78.490 296.255 78.645 ;
        RECT 296.040 78.260 296.330 78.490 ;
        RECT 298.320 78.445 298.970 78.490 ;
        RECT 301.920 78.445 302.210 78.490 ;
        RECT 303.385 78.445 303.705 78.505 ;
        RECT 298.320 78.305 303.705 78.445 ;
        RECT 298.320 78.260 298.970 78.305 ;
        RECT 301.620 78.260 302.210 78.305 ;
        RECT 285.905 78.105 286.225 78.165 ;
        RECT 283.465 77.965 286.225 78.105 ;
        RECT 285.905 77.905 286.225 77.965 ;
        RECT 290.965 77.905 291.285 78.165 ;
        RECT 294.645 77.905 294.965 78.165 ;
        RECT 295.125 78.105 295.415 78.150 ;
        RECT 296.960 78.105 297.250 78.150 ;
        RECT 300.540 78.105 300.830 78.150 ;
        RECT 295.125 77.965 300.830 78.105 ;
        RECT 295.125 77.920 295.415 77.965 ;
        RECT 296.960 77.920 297.250 77.965 ;
        RECT 300.540 77.920 300.830 77.965 ;
        RECT 301.620 77.945 301.910 78.260 ;
        RECT 303.385 78.245 303.705 78.305 ;
        RECT 297.865 77.765 298.185 77.825 ;
        RECT 259.790 77.625 260.835 77.765 ;
        RECT 259.790 77.470 259.930 77.625 ;
        RECT 259.700 77.240 259.990 77.470 ;
        RECT 260.695 77.425 260.835 77.625 ;
        RECT 261.065 77.625 298.185 77.765 ;
        RECT 261.065 77.565 261.385 77.625 ;
        RECT 297.865 77.565 298.185 77.625 ;
        RECT 303.400 77.765 303.690 77.810 ;
        RECT 305.685 77.765 306.005 77.825 ;
        RECT 303.400 77.625 306.005 77.765 ;
        RECT 303.400 77.580 303.690 77.625 ;
        RECT 305.685 77.565 306.005 77.625 ;
        RECT 261.985 77.425 262.305 77.485 ;
        RECT 260.695 77.285 262.305 77.425 ;
        RECT 261.985 77.225 262.305 77.285 ;
        RECT 273.450 77.425 273.740 77.470 ;
        RECT 275.340 77.425 275.630 77.470 ;
        RECT 278.460 77.425 278.750 77.470 ;
        RECT 273.450 77.285 278.750 77.425 ;
        RECT 273.450 77.240 273.740 77.285 ;
        RECT 275.340 77.240 275.630 77.285 ;
        RECT 278.460 77.240 278.750 77.285 ;
        RECT 295.530 77.425 295.820 77.470 ;
        RECT 297.420 77.425 297.710 77.470 ;
        RECT 300.540 77.425 300.830 77.470 ;
        RECT 295.530 77.285 300.830 77.425 ;
        RECT 295.530 77.240 295.820 77.285 ;
        RECT 297.420 77.240 297.710 77.285 ;
        RECT 300.540 77.240 300.830 77.285 ;
        RECT 242.205 76.945 245.195 77.085 ;
        RECT 246.360 77.085 246.650 77.130 ;
        RECT 246.820 77.085 247.110 77.130 ;
        RECT 246.360 76.945 247.110 77.085 ;
        RECT 178.265 76.885 178.585 76.945 ;
        RECT 188.385 76.885 188.705 76.945 ;
        RECT 196.665 76.885 196.985 76.945 ;
        RECT 197.140 76.900 197.430 76.945 ;
        RECT 200.805 76.885 201.125 76.945 ;
        RECT 236.225 76.885 236.545 76.945 ;
        RECT 242.205 76.885 242.525 76.945 ;
        RECT 244.505 76.885 244.825 76.945 ;
        RECT 246.360 76.900 246.650 76.945 ;
        RECT 246.820 76.900 247.110 76.945 ;
        RECT 248.645 76.885 248.965 77.145 ;
        RECT 258.765 76.885 259.085 77.145 ;
        RECT 262.905 77.085 263.225 77.145 ;
        RECT 263.380 77.085 263.670 77.130 ;
        RECT 262.905 76.945 263.670 77.085 ;
        RECT 262.905 76.885 263.225 76.945 ;
        RECT 263.380 76.900 263.670 76.945 ;
        RECT 276.245 77.085 276.565 77.145 ;
        RECT 281.320 77.085 281.610 77.130 ;
        RECT 276.245 76.945 281.610 77.085 ;
        RECT 276.245 76.885 276.565 76.945 ;
        RECT 281.320 76.900 281.610 76.945 ;
        RECT 162.095 76.265 311.135 76.745 ;
        RECT 172.745 75.865 173.065 76.125 ;
        RECT 173.205 76.065 173.525 76.125 ;
        RECT 175.980 76.065 176.270 76.110 ;
        RECT 173.205 75.925 176.270 76.065 ;
        RECT 173.205 75.865 173.525 75.925 ;
        RECT 175.980 75.880 176.270 75.925 ;
        RECT 194.365 76.065 194.685 76.125 ;
        RECT 195.300 76.065 195.590 76.110 ;
        RECT 194.365 75.925 195.590 76.065 ;
        RECT 194.365 75.865 194.685 75.925 ;
        RECT 195.300 75.880 195.590 75.925 ;
        RECT 196.205 76.065 196.525 76.125 ;
        RECT 200.805 76.065 201.125 76.125 ;
        RECT 202.200 76.065 202.490 76.110 ;
        RECT 196.205 75.925 199.195 76.065 ;
        RECT 196.205 75.865 196.525 75.925 ;
        RECT 166.270 75.725 166.560 75.770 ;
        RECT 168.160 75.725 168.450 75.770 ;
        RECT 171.280 75.725 171.570 75.770 ;
        RECT 172.835 75.725 172.975 75.865 ;
        RECT 179.185 75.725 179.505 75.785 ;
        RECT 166.270 75.585 171.570 75.725 ;
        RECT 166.270 75.540 166.560 75.585 ;
        RECT 168.160 75.540 168.450 75.585 ;
        RECT 171.280 75.540 171.570 75.585 ;
        RECT 172.375 75.585 179.505 75.725 ;
        RECT 166.780 75.385 167.070 75.430 ;
        RECT 169.525 75.385 169.845 75.445 ;
        RECT 166.780 75.245 169.845 75.385 ;
        RECT 166.780 75.200 167.070 75.245 ;
        RECT 169.525 75.185 169.845 75.245 ;
        RECT 165.385 74.845 165.705 75.105 ;
        RECT 165.865 75.045 166.155 75.090 ;
        RECT 167.700 75.045 167.990 75.090 ;
        RECT 171.280 75.045 171.570 75.090 ;
        RECT 172.375 75.065 172.515 75.585 ;
        RECT 179.185 75.525 179.505 75.585 ;
        RECT 186.510 75.725 186.800 75.770 ;
        RECT 188.400 75.725 188.690 75.770 ;
        RECT 191.520 75.725 191.810 75.770 ;
        RECT 186.510 75.585 191.810 75.725 ;
        RECT 186.510 75.540 186.800 75.585 ;
        RECT 188.400 75.540 188.690 75.585 ;
        RECT 191.520 75.540 191.810 75.585 ;
        RECT 196.665 75.725 196.985 75.785 ;
        RECT 199.055 75.725 199.195 75.925 ;
        RECT 200.805 75.925 202.490 76.065 ;
        RECT 200.805 75.865 201.125 75.925 ;
        RECT 202.200 75.880 202.490 75.925 ;
        RECT 208.625 75.865 208.945 76.125 ;
        RECT 213.685 76.065 214.005 76.125 ;
        RECT 215.065 76.065 215.385 76.125 ;
        RECT 213.685 75.925 215.385 76.065 ;
        RECT 213.685 75.865 214.005 75.925 ;
        RECT 215.065 75.865 215.385 75.925 ;
        RECT 219.205 75.865 219.525 76.125 ;
        RECT 227.025 75.865 227.345 76.125 ;
        RECT 227.485 76.065 227.805 76.125 ;
        RECT 237.160 76.065 237.450 76.110 ;
        RECT 239.905 76.065 240.225 76.125 ;
        RECT 227.485 75.925 236.915 76.065 ;
        RECT 227.485 75.865 227.805 75.925 ;
        RECT 196.665 75.585 198.275 75.725 ;
        RECT 199.055 75.585 201.495 75.725 ;
        RECT 196.665 75.525 196.985 75.585 ;
        RECT 177.805 75.185 178.125 75.445 ;
        RECT 178.265 75.185 178.585 75.445 ;
        RECT 178.725 75.185 179.045 75.445 ;
        RECT 179.275 75.385 179.415 75.525 ;
        RECT 179.275 75.245 185.395 75.385 ;
        RECT 165.865 74.905 171.570 75.045 ;
        RECT 165.865 74.860 166.155 74.905 ;
        RECT 167.700 74.860 167.990 74.905 ;
        RECT 171.280 74.860 171.570 74.905 ;
        RECT 172.360 74.750 172.650 75.065 ;
        RECT 177.895 75.045 178.035 75.185 ;
        RECT 181.040 75.045 181.330 75.090 ;
        RECT 181.945 75.045 182.265 75.105 ;
        RECT 177.895 74.905 182.265 75.045 ;
        RECT 185.255 75.045 185.395 75.245 ;
        RECT 185.625 75.185 185.945 75.445 ;
        RECT 187.005 75.185 187.325 75.445 ;
        RECT 192.065 75.385 192.385 75.445 ;
        RECT 192.065 75.245 193.675 75.385 ;
        RECT 192.065 75.185 192.385 75.245 ;
        RECT 186.105 75.045 186.395 75.090 ;
        RECT 187.940 75.045 188.230 75.090 ;
        RECT 191.520 75.045 191.810 75.090 ;
        RECT 185.255 74.905 185.855 75.045 ;
        RECT 181.040 74.860 181.330 74.905 ;
        RECT 181.945 74.845 182.265 74.905 ;
        RECT 169.060 74.705 169.710 74.750 ;
        RECT 172.360 74.705 172.950 74.750 ;
        RECT 179.185 74.705 179.505 74.765 ;
        RECT 169.060 74.565 172.950 74.705 ;
        RECT 169.060 74.520 169.710 74.565 ;
        RECT 172.660 74.520 172.950 74.565 ;
        RECT 174.215 74.565 179.505 74.705 ;
        RECT 174.215 74.410 174.355 74.565 ;
        RECT 179.185 74.505 179.505 74.565 ;
        RECT 185.180 74.520 185.470 74.750 ;
        RECT 185.715 74.705 185.855 74.905 ;
        RECT 186.105 74.905 191.810 75.045 ;
        RECT 186.105 74.860 186.395 74.905 ;
        RECT 187.940 74.860 188.230 74.905 ;
        RECT 191.520 74.860 191.810 74.905 ;
        RECT 188.385 74.705 188.705 74.765 ;
        RECT 192.600 74.750 192.890 75.065 ;
        RECT 189.300 74.705 189.950 74.750 ;
        RECT 192.600 74.705 193.190 74.750 ;
        RECT 185.715 74.565 193.190 74.705 ;
        RECT 193.535 74.705 193.675 75.245 ;
        RECT 195.285 75.185 195.605 75.445 ;
        RECT 198.135 75.430 198.275 75.585 ;
        RECT 198.060 75.200 198.350 75.430 ;
        RECT 195.375 75.045 195.515 75.185 ;
        RECT 201.355 75.105 201.495 75.585 ;
        RECT 208.715 75.385 208.855 75.865 ;
        RECT 210.020 75.725 210.310 75.770 ;
        RECT 223.345 75.725 223.665 75.785 ;
        RECT 226.120 75.725 226.410 75.770 ;
        RECT 227.575 75.725 227.715 75.865 ;
        RECT 210.020 75.585 221.505 75.725 ;
        RECT 210.020 75.540 210.310 75.585 ;
        RECT 206.875 75.245 208.855 75.385 ;
        RECT 211.845 75.385 212.165 75.445 ;
        RECT 216.000 75.385 216.290 75.430 ;
        RECT 220.125 75.385 220.445 75.445 ;
        RECT 211.845 75.245 220.445 75.385 ;
        RECT 221.365 75.385 221.505 75.585 ;
        RECT 223.345 75.585 225.875 75.725 ;
        RECT 223.345 75.525 223.665 75.585 ;
        RECT 221.365 75.245 224.495 75.385 ;
        RECT 197.600 75.045 197.890 75.090 ;
        RECT 195.375 74.905 197.890 75.045 ;
        RECT 197.600 74.860 197.890 74.905 ;
        RECT 197.675 74.705 197.815 74.860 ;
        RECT 200.345 74.845 200.665 75.105 ;
        RECT 201.265 75.045 201.585 75.105 ;
        RECT 206.875 75.090 207.015 75.245 ;
        RECT 211.845 75.185 212.165 75.245 ;
        RECT 216.000 75.200 216.290 75.245 ;
        RECT 220.125 75.185 220.445 75.245 ;
        RECT 209.085 75.090 209.405 75.105 ;
        RECT 201.740 75.045 202.030 75.090 ;
        RECT 201.265 74.905 202.030 75.045 ;
        RECT 201.265 74.845 201.585 74.905 ;
        RECT 201.740 74.860 202.030 74.905 ;
        RECT 206.800 74.860 207.090 75.090 ;
        RECT 207.265 74.860 207.555 75.090 ;
        RECT 209.085 75.045 209.415 75.090 ;
        RECT 209.085 74.905 209.600 75.045 ;
        RECT 209.085 74.860 209.415 74.905 ;
        RECT 193.535 74.565 197.355 74.705 ;
        RECT 197.675 74.565 201.495 74.705 ;
        RECT 174.140 74.180 174.430 74.410 ;
        RECT 177.805 74.165 178.125 74.425 ;
        RECT 185.255 74.365 185.395 74.520 ;
        RECT 188.385 74.505 188.705 74.565 ;
        RECT 189.300 74.520 189.950 74.565 ;
        RECT 192.900 74.520 193.190 74.565 ;
        RECT 197.215 74.425 197.355 74.565 ;
        RECT 193.445 74.365 193.765 74.425 ;
        RECT 185.255 74.225 193.765 74.365 ;
        RECT 193.445 74.165 193.765 74.225 ;
        RECT 194.365 74.165 194.685 74.425 ;
        RECT 197.125 74.165 197.445 74.425 ;
        RECT 198.045 74.365 198.365 74.425 ;
        RECT 199.440 74.365 199.730 74.410 ;
        RECT 198.045 74.225 199.730 74.365 ;
        RECT 201.355 74.365 201.495 74.565 ;
        RECT 207.335 74.365 207.475 74.860 ;
        RECT 209.085 74.845 209.405 74.860 ;
        RECT 214.145 74.845 214.465 75.105 ;
        RECT 216.445 75.045 216.765 75.105 ;
        RECT 217.380 75.045 217.670 75.090 ;
        RECT 216.445 74.905 217.670 75.045 ;
        RECT 216.445 74.845 216.765 74.905 ;
        RECT 217.380 74.860 217.670 74.905 ;
        RECT 219.680 74.860 219.970 75.090 ;
        RECT 208.180 74.520 208.470 74.750 ;
        RECT 208.640 74.705 208.930 74.750 ;
        RECT 214.235 74.705 214.375 74.845 ;
        RECT 208.640 74.565 214.375 74.705 ;
        RECT 214.620 74.705 214.910 74.750 ;
        RECT 218.425 74.705 218.715 74.750 ;
        RECT 219.205 74.705 219.525 74.765 ;
        RECT 214.620 74.565 219.525 74.705 ;
        RECT 219.755 74.705 219.895 74.860 ;
        RECT 221.965 74.845 222.285 75.105 ;
        RECT 223.360 75.045 223.650 75.090 ;
        RECT 223.805 75.045 224.125 75.105 ;
        RECT 223.360 74.905 224.125 75.045 ;
        RECT 223.360 74.860 223.650 74.905 ;
        RECT 222.425 74.705 222.745 74.765 ;
        RECT 219.755 74.565 222.745 74.705 ;
        RECT 208.640 74.520 208.930 74.565 ;
        RECT 214.620 74.520 214.910 74.565 ;
        RECT 218.425 74.520 218.715 74.565 ;
        RECT 201.355 74.225 207.475 74.365 ;
        RECT 208.255 74.365 208.395 74.520 ;
        RECT 219.205 74.505 219.525 74.565 ;
        RECT 222.425 74.505 222.745 74.565 ;
        RECT 210.005 74.365 210.325 74.425 ;
        RECT 208.255 74.225 210.325 74.365 ;
        RECT 198.045 74.165 198.365 74.225 ;
        RECT 199.440 74.180 199.730 74.225 ;
        RECT 210.005 74.165 210.325 74.225 ;
        RECT 215.065 74.365 215.385 74.425 ;
        RECT 215.985 74.365 216.305 74.425 ;
        RECT 215.065 74.225 216.305 74.365 ;
        RECT 215.065 74.165 215.385 74.225 ;
        RECT 215.985 74.165 216.305 74.225 ;
        RECT 217.840 74.365 218.130 74.410 ;
        RECT 223.435 74.365 223.575 74.860 ;
        RECT 223.805 74.845 224.125 74.905 ;
        RECT 224.355 74.705 224.495 75.245 ;
        RECT 224.725 75.185 225.045 75.445 ;
        RECT 225.735 75.385 225.875 75.585 ;
        RECT 226.120 75.585 227.715 75.725 ;
        RECT 228.880 75.725 229.170 75.770 ;
        RECT 235.305 75.725 235.625 75.785 ;
        RECT 228.880 75.585 235.625 75.725 ;
        RECT 236.775 75.725 236.915 75.925 ;
        RECT 237.160 75.925 240.225 76.065 ;
        RECT 237.160 75.880 237.450 75.925 ;
        RECT 239.905 75.865 240.225 75.925 ;
        RECT 243.125 75.865 243.445 76.125 ;
        RECT 250.945 76.065 251.265 76.125 ;
        RECT 261.065 76.065 261.385 76.125 ;
        RECT 250.945 75.925 261.385 76.065 ;
        RECT 250.945 75.865 251.265 75.925 ;
        RECT 261.065 75.865 261.385 75.925 ;
        RECT 261.540 76.065 261.830 76.110 ;
        RECT 261.985 76.065 262.305 76.125 ;
        RECT 261.540 75.925 262.305 76.065 ;
        RECT 261.540 75.880 261.830 75.925 ;
        RECT 261.985 75.865 262.305 75.925 ;
        RECT 262.920 75.880 263.210 76.110 ;
        RECT 273.960 76.065 274.250 76.110 ;
        RECT 275.325 76.065 275.645 76.125 ;
        RECT 273.960 75.925 275.645 76.065 ;
        RECT 273.960 75.880 274.250 75.925 ;
        RECT 245.425 75.725 245.745 75.785 ;
        RECT 259.225 75.725 259.545 75.785 ;
        RECT 236.775 75.585 259.545 75.725 ;
        RECT 226.120 75.540 226.410 75.585 ;
        RECT 228.880 75.540 229.170 75.585 ;
        RECT 235.305 75.525 235.625 75.585 ;
        RECT 245.425 75.525 245.745 75.585 ;
        RECT 259.225 75.525 259.545 75.585 ;
        RECT 260.160 75.725 260.450 75.770 ;
        RECT 262.995 75.725 263.135 75.880 ;
        RECT 275.325 75.865 275.645 75.925 ;
        RECT 278.545 75.865 278.865 76.125 ;
        RECT 280.845 76.065 281.165 76.125 ;
        RECT 304.320 76.065 304.610 76.110 ;
        RECT 305.225 76.065 305.545 76.125 ;
        RECT 280.845 75.925 285.675 76.065 ;
        RECT 280.845 75.865 281.165 75.925 ;
        RECT 280.935 75.725 281.075 75.865 ;
        RECT 260.160 75.585 263.135 75.725 ;
        RECT 269.665 75.585 281.075 75.725 ;
        RECT 260.160 75.540 260.450 75.585 ;
        RECT 227.500 75.385 227.790 75.430 ;
        RECT 233.925 75.385 234.245 75.445 ;
        RECT 225.735 75.245 227.790 75.385 ;
        RECT 227.500 75.200 227.790 75.245 ;
        RECT 228.035 75.245 234.245 75.385 ;
        RECT 224.815 75.045 224.955 75.185 ;
        RECT 228.035 75.105 228.175 75.245 ;
        RECT 233.925 75.185 234.245 75.245 ;
        RECT 237.145 75.185 237.465 75.445 ;
        RECT 239.445 75.385 239.765 75.445 ;
        RECT 242.680 75.385 242.970 75.430 ;
        RECT 246.805 75.385 247.125 75.445 ;
        RECT 269.665 75.385 269.805 75.585 ;
        RECT 239.445 75.245 242.435 75.385 ;
        RECT 239.445 75.185 239.765 75.245 ;
        RECT 227.040 75.045 227.330 75.090 ;
        RECT 224.815 74.905 227.330 75.045 ;
        RECT 227.040 74.860 227.330 74.905 ;
        RECT 227.945 74.845 228.265 75.105 ;
        RECT 232.545 75.045 232.865 75.105 ;
        RECT 235.320 75.045 235.610 75.090 ;
        RECT 232.545 74.905 235.610 75.045 ;
        RECT 232.545 74.845 232.865 74.905 ;
        RECT 235.320 74.860 235.610 74.905 ;
        RECT 236.365 75.045 236.655 75.090 ;
        RECT 237.235 75.045 237.375 75.185 ;
        RECT 236.365 74.905 237.375 75.045 ;
        RECT 236.365 74.860 236.655 74.905 ;
        RECT 238.985 74.845 239.305 75.105 ;
        RECT 242.295 75.090 242.435 75.245 ;
        RECT 242.680 75.245 247.125 75.385 ;
        RECT 242.680 75.200 242.970 75.245 ;
        RECT 246.805 75.185 247.125 75.245 ;
        RECT 257.475 75.245 269.805 75.385 ;
        RECT 275.325 75.385 275.645 75.445 ;
        RECT 276.720 75.385 277.010 75.430 ;
        RECT 281.320 75.385 281.610 75.430 ;
        RECT 275.325 75.245 281.610 75.385 ;
        RECT 242.220 74.860 242.510 75.090 ;
        RECT 243.585 74.845 243.905 75.105 ;
        RECT 245.885 75.045 246.205 75.105 ;
        RECT 248.645 75.045 248.965 75.105 ;
        RECT 245.885 74.905 248.965 75.045 ;
        RECT 245.885 74.845 246.205 74.905 ;
        RECT 248.645 74.845 248.965 74.905 ;
        RECT 253.705 75.045 254.025 75.105 ;
        RECT 257.475 75.090 257.615 75.245 ;
        RECT 275.325 75.185 275.645 75.245 ;
        RECT 276.720 75.200 277.010 75.245 ;
        RECT 281.320 75.200 281.610 75.245 ;
        RECT 281.765 75.185 282.085 75.445 ;
        RECT 257.400 75.045 257.690 75.090 ;
        RECT 253.705 74.905 257.690 75.045 ;
        RECT 253.705 74.845 254.025 74.905 ;
        RECT 257.400 74.860 257.690 74.905 ;
        RECT 259.225 74.845 259.545 75.105 ;
        RECT 260.605 74.845 260.925 75.105 ;
        RECT 261.065 74.845 261.385 75.105 ;
        RECT 262.905 74.845 263.225 75.105 ;
        RECT 263.380 74.860 263.670 75.090 ;
        RECT 233.465 74.705 233.785 74.765 ;
        RECT 235.780 74.705 236.070 74.750 ;
        RECT 237.605 74.705 237.925 74.765 ;
        RECT 224.355 74.565 229.555 74.705 ;
        RECT 229.415 74.425 229.555 74.565 ;
        RECT 233.465 74.565 237.925 74.705 ;
        RECT 239.075 74.705 239.215 74.845 ;
        RECT 243.675 74.705 243.815 74.845 ;
        RECT 239.075 74.565 243.815 74.705 ;
        RECT 247.265 74.705 247.585 74.765 ;
        RECT 256.925 74.705 257.245 74.765 ;
        RECT 258.320 74.705 258.610 74.750 ;
        RECT 247.265 74.565 258.610 74.705 ;
        RECT 233.465 74.505 233.785 74.565 ;
        RECT 235.780 74.520 236.070 74.565 ;
        RECT 237.605 74.505 237.925 74.565 ;
        RECT 247.265 74.505 247.585 74.565 ;
        RECT 256.925 74.505 257.245 74.565 ;
        RECT 258.320 74.520 258.610 74.565 ;
        RECT 258.765 74.505 259.085 74.765 ;
        RECT 263.455 74.705 263.595 74.860 ;
        RECT 275.785 74.845 276.105 75.105 ;
        RECT 276.245 74.845 276.565 75.105 ;
        RECT 280.860 75.045 281.150 75.090 ;
        RECT 281.855 75.045 281.995 75.185 ;
        RECT 280.860 74.905 281.995 75.045 ;
        RECT 280.860 74.860 281.150 74.905 ;
        RECT 284.985 74.845 285.305 75.105 ;
        RECT 285.535 75.045 285.675 75.925 ;
        RECT 304.320 75.925 305.545 76.065 ;
        RECT 304.320 75.880 304.610 75.925 ;
        RECT 305.225 75.865 305.545 75.925 ;
        RECT 285.920 75.540 286.210 75.770 ;
        RECT 289.240 75.725 289.530 75.770 ;
        RECT 292.360 75.725 292.650 75.770 ;
        RECT 294.250 75.725 294.540 75.770 ;
        RECT 289.240 75.585 294.540 75.725 ;
        RECT 289.240 75.540 289.530 75.585 ;
        RECT 292.360 75.540 292.650 75.585 ;
        RECT 294.250 75.540 294.540 75.585 ;
        RECT 285.995 75.385 286.135 75.540 ;
        RECT 299.705 75.525 300.025 75.785 ;
        RECT 293.740 75.385 294.030 75.430 ;
        RECT 285.995 75.245 294.030 75.385 ;
        RECT 293.740 75.200 294.030 75.245 ;
        RECT 296.500 75.385 296.790 75.430 ;
        RECT 298.325 75.385 298.645 75.445 ;
        RECT 307.080 75.385 307.370 75.430 ;
        RECT 296.500 75.245 307.370 75.385 ;
        RECT 296.500 75.200 296.790 75.245 ;
        RECT 285.535 74.905 286.595 75.045 ;
        RECT 259.315 74.565 263.595 74.705 ;
        RECT 275.875 74.705 276.015 74.845 ;
        RECT 284.065 74.705 284.385 74.765 ;
        RECT 275.875 74.565 284.385 74.705 ;
        RECT 217.840 74.225 223.575 74.365 ;
        RECT 217.840 74.180 218.130 74.225 ;
        RECT 229.325 74.165 229.645 74.425 ;
        RECT 236.685 74.365 237.005 74.425 ;
        RECT 238.985 74.365 239.305 74.425 ;
        RECT 236.685 74.225 239.305 74.365 ;
        RECT 236.685 74.165 237.005 74.225 ;
        RECT 238.985 74.165 239.305 74.225 ;
        RECT 239.445 74.365 239.765 74.425 ;
        RECT 240.825 74.365 241.145 74.425 ;
        RECT 239.445 74.225 241.145 74.365 ;
        RECT 239.445 74.165 239.765 74.225 ;
        RECT 240.825 74.165 241.145 74.225 ;
        RECT 244.045 74.165 244.365 74.425 ;
        RECT 248.645 74.365 248.965 74.425 ;
        RECT 259.315 74.365 259.455 74.565 ;
        RECT 284.065 74.505 284.385 74.565 ;
        RECT 248.645 74.225 259.455 74.365 ;
        RECT 248.645 74.165 248.965 74.225 ;
        RECT 262.445 74.165 262.765 74.425 ;
        RECT 262.905 74.365 263.225 74.425 ;
        RECT 264.760 74.365 265.050 74.410 ;
        RECT 262.905 74.225 265.050 74.365 ;
        RECT 262.905 74.165 263.225 74.225 ;
        RECT 264.760 74.180 265.050 74.225 ;
        RECT 280.400 74.365 280.690 74.410 ;
        RECT 284.525 74.365 284.845 74.425 ;
        RECT 286.455 74.410 286.595 74.905 ;
        RECT 288.160 74.750 288.450 75.065 ;
        RECT 289.240 75.045 289.530 75.090 ;
        RECT 292.820 75.045 293.110 75.090 ;
        RECT 294.655 75.045 294.945 75.090 ;
        RECT 289.240 74.905 294.945 75.045 ;
        RECT 289.240 74.860 289.530 74.905 ;
        RECT 292.820 74.860 293.110 74.905 ;
        RECT 294.655 74.860 294.945 74.905 ;
        RECT 295.120 74.860 295.410 75.090 ;
        RECT 287.860 74.705 288.450 74.750 ;
        RECT 290.965 74.750 291.285 74.765 ;
        RECT 290.965 74.705 291.750 74.750 ;
        RECT 295.195 74.705 295.335 74.860 ;
        RECT 287.860 74.565 291.750 74.705 ;
        RECT 287.860 74.520 288.150 74.565 ;
        RECT 290.965 74.520 291.750 74.565 ;
        RECT 294.275 74.565 295.335 74.705 ;
        RECT 290.965 74.505 291.285 74.520 ;
        RECT 294.275 74.425 294.415 74.565 ;
        RECT 280.400 74.225 284.845 74.365 ;
        RECT 280.400 74.180 280.690 74.225 ;
        RECT 284.525 74.165 284.845 74.225 ;
        RECT 286.380 74.365 286.670 74.410 ;
        RECT 288.665 74.365 288.985 74.425 ;
        RECT 286.380 74.225 288.985 74.365 ;
        RECT 286.380 74.180 286.670 74.225 ;
        RECT 288.665 74.165 288.985 74.225 ;
        RECT 294.185 74.165 294.505 74.425 ;
        RECT 294.645 74.365 294.965 74.425 ;
        RECT 296.575 74.365 296.715 75.200 ;
        RECT 298.325 75.185 298.645 75.245 ;
        RECT 307.080 75.200 307.370 75.245 ;
        RECT 299.705 75.045 300.025 75.105 ;
        RECT 301.100 75.045 301.390 75.090 ;
        RECT 299.705 74.905 301.390 75.045 ;
        RECT 299.705 74.845 300.025 74.905 ;
        RECT 301.100 74.860 301.390 74.905 ;
        RECT 301.545 75.045 301.865 75.105 ;
        RECT 306.160 75.045 306.450 75.090 ;
        RECT 301.545 74.905 306.450 75.045 ;
        RECT 301.545 74.845 301.865 74.905 ;
        RECT 306.160 74.860 306.450 74.905 ;
        RECT 297.865 74.705 298.185 74.765 ;
        RECT 304.765 74.705 305.085 74.765 ;
        RECT 297.865 74.565 305.085 74.705 ;
        RECT 297.865 74.505 298.185 74.565 ;
        RECT 304.765 74.505 305.085 74.565 ;
        RECT 294.645 74.225 296.715 74.365 ;
        RECT 294.645 74.165 294.965 74.225 ;
        RECT 297.405 74.165 297.725 74.425 ;
        RECT 298.325 74.365 298.645 74.425 ;
        RECT 300.180 74.365 300.470 74.410 ;
        RECT 298.325 74.225 300.470 74.365 ;
        RECT 298.325 74.165 298.645 74.225 ;
        RECT 300.180 74.180 300.470 74.225 ;
        RECT 306.605 74.165 306.925 74.425 ;
        RECT 162.095 73.545 311.935 74.025 ;
        RECT 174.125 73.345 174.445 73.405 ;
        RECT 177.360 73.345 177.650 73.390 ;
        RECT 174.125 73.205 177.650 73.345 ;
        RECT 174.125 73.145 174.445 73.205 ;
        RECT 177.360 73.160 177.650 73.205 ;
        RECT 179.185 73.145 179.505 73.405 ;
        RECT 184.705 73.345 185.025 73.405 ;
        RECT 185.180 73.345 185.470 73.390 ;
        RECT 192.065 73.345 192.385 73.405 ;
        RECT 184.705 73.205 185.470 73.345 ;
        RECT 184.705 73.145 185.025 73.205 ;
        RECT 185.180 73.160 185.470 73.205 ;
        RECT 187.095 73.205 192.385 73.345 ;
        RECT 177.805 73.005 178.125 73.065 ;
        RECT 187.095 73.005 187.235 73.205 ;
        RECT 192.065 73.145 192.385 73.205 ;
        RECT 197.125 73.345 197.445 73.405 ;
        RECT 219.665 73.345 219.985 73.405 ;
        RECT 221.965 73.345 222.285 73.405 ;
        RECT 232.085 73.345 232.405 73.405 ;
        RECT 243.140 73.345 243.430 73.390 ;
        RECT 248.645 73.345 248.965 73.405 ;
        RECT 197.125 73.205 219.985 73.345 ;
        RECT 197.125 73.145 197.445 73.205 ;
        RECT 219.665 73.145 219.985 73.205 ;
        RECT 220.675 73.205 227.255 73.345 ;
        RECT 175.135 72.865 177.575 73.005 ;
        RECT 175.135 72.725 175.275 72.865 ;
        RECT 170.920 72.665 171.210 72.710 ;
        RECT 170.920 72.525 173.435 72.665 ;
        RECT 170.920 72.480 171.210 72.525 ;
        RECT 173.295 72.030 173.435 72.525 ;
        RECT 175.045 72.465 175.365 72.725 ;
        RECT 175.505 72.465 175.825 72.725 ;
        RECT 177.435 72.665 177.575 72.865 ;
        RECT 177.805 72.865 187.235 73.005 ;
        RECT 187.465 73.005 187.785 73.065 ;
        RECT 188.860 73.005 189.150 73.050 ;
        RECT 187.465 72.865 189.150 73.005 ;
        RECT 177.805 72.805 178.125 72.865 ;
        RECT 187.465 72.805 187.785 72.865 ;
        RECT 188.860 72.820 189.150 72.865 ;
        RECT 193.000 73.005 193.290 73.050 ;
        RECT 193.445 73.005 193.765 73.065 ;
        RECT 194.825 73.005 195.145 73.065 ;
        RECT 220.675 73.050 220.815 73.205 ;
        RECT 221.965 73.145 222.285 73.205 ;
        RECT 227.115 73.065 227.255 73.205 ;
        RECT 232.085 73.205 241.515 73.345 ;
        RECT 232.085 73.145 232.405 73.205 ;
        RECT 222.425 73.050 222.745 73.065 ;
        RECT 193.000 72.865 195.145 73.005 ;
        RECT 193.000 72.820 193.290 72.865 ;
        RECT 193.445 72.805 193.765 72.865 ;
        RECT 194.825 72.805 195.145 72.865 ;
        RECT 197.580 73.005 198.230 73.050 ;
        RECT 201.180 73.005 201.470 73.050 ;
        RECT 197.580 72.865 201.470 73.005 ;
        RECT 197.580 72.820 198.230 72.865 ;
        RECT 200.880 72.820 201.470 72.865 ;
        RECT 220.600 72.820 220.890 73.050 ;
        RECT 222.425 73.005 222.775 73.050 ;
        RECT 222.425 72.865 222.940 73.005 ;
        RECT 222.425 72.820 222.775 72.865 ;
        RECT 200.880 72.725 201.170 72.820 ;
        RECT 222.425 72.805 222.745 72.820 ;
        RECT 227.025 72.805 227.345 73.065 ;
        RECT 230.245 73.005 230.565 73.065 ;
        RECT 241.375 73.050 241.515 73.205 ;
        RECT 243.140 73.205 248.965 73.345 ;
        RECT 243.140 73.160 243.430 73.205 ;
        RECT 248.645 73.145 248.965 73.205 ;
        RECT 258.320 73.345 258.610 73.390 ;
        RECT 261.065 73.345 261.385 73.405 ;
        RECT 258.320 73.205 261.385 73.345 ;
        RECT 258.320 73.160 258.610 73.205 ;
        RECT 261.065 73.145 261.385 73.205 ;
        RECT 271.645 73.345 271.965 73.405 ;
        RECT 284.525 73.345 284.845 73.405 ;
        RECT 286.365 73.345 286.685 73.405 ;
        RECT 293.725 73.345 294.045 73.405 ;
        RECT 271.645 73.205 277.855 73.345 ;
        RECT 271.645 73.145 271.965 73.205 ;
        RECT 241.300 73.005 241.590 73.050 ;
        RECT 256.480 73.005 256.770 73.050 ;
        RECT 230.245 72.865 240.600 73.005 ;
        RECT 230.245 72.805 230.565 72.865 ;
        RECT 233.555 72.725 233.695 72.865 ;
        RECT 185.640 72.665 185.930 72.710 ;
        RECT 192.525 72.665 192.845 72.725 ;
        RECT 177.435 72.525 192.845 72.665 ;
        RECT 185.640 72.480 185.930 72.525 ;
        RECT 192.525 72.465 192.845 72.525 ;
        RECT 193.905 72.465 194.225 72.725 ;
        RECT 194.385 72.665 194.675 72.710 ;
        RECT 196.220 72.665 196.510 72.710 ;
        RECT 199.800 72.665 200.090 72.710 ;
        RECT 194.385 72.525 200.090 72.665 ;
        RECT 194.385 72.480 194.675 72.525 ;
        RECT 196.220 72.480 196.510 72.525 ;
        RECT 199.800 72.480 200.090 72.525 ;
        RECT 200.805 72.505 201.170 72.725 ;
        RECT 204.500 72.665 204.790 72.710 ;
        RECT 205.405 72.665 205.725 72.725 ;
        RECT 204.500 72.525 205.725 72.665 ;
        RECT 200.805 72.465 201.125 72.505 ;
        RECT 204.500 72.480 204.790 72.525 ;
        RECT 205.405 72.465 205.725 72.525 ;
        RECT 205.880 72.665 206.170 72.710 ;
        RECT 207.245 72.665 207.565 72.725 ;
        RECT 223.820 72.665 224.110 72.710 ;
        RECT 229.785 72.665 230.105 72.725 ;
        RECT 205.880 72.525 223.575 72.665 ;
        RECT 205.880 72.480 206.170 72.525 ;
        RECT 176.425 72.125 176.745 72.385 ;
        RECT 177.345 72.325 177.665 72.385 ;
        RECT 178.265 72.325 178.585 72.385 ;
        RECT 179.660 72.325 179.950 72.370 ;
        RECT 177.345 72.185 179.950 72.325 ;
        RECT 177.345 72.125 177.665 72.185 ;
        RECT 178.265 72.125 178.585 72.185 ;
        RECT 179.660 72.140 179.950 72.185 ;
        RECT 180.120 72.140 180.410 72.370 ;
        RECT 184.720 72.325 185.010 72.370 ;
        RECT 193.445 72.325 193.765 72.385 ;
        RECT 184.720 72.185 193.765 72.325 ;
        RECT 184.720 72.140 185.010 72.185 ;
        RECT 173.220 71.800 173.510 72.030 ;
        RECT 180.195 71.985 180.335 72.140 ;
        RECT 193.445 72.125 193.765 72.185 ;
        RECT 195.300 72.325 195.590 72.370 ;
        RECT 198.045 72.325 198.365 72.385 ;
        RECT 202.645 72.325 202.965 72.385 ;
        RECT 195.300 72.185 198.365 72.325 ;
        RECT 195.300 72.140 195.590 72.185 ;
        RECT 198.045 72.125 198.365 72.185 ;
        RECT 200.435 72.185 202.965 72.325 ;
        RECT 178.815 71.845 180.335 71.985 ;
        RECT 194.790 71.985 195.080 72.030 ;
        RECT 196.680 71.985 196.970 72.030 ;
        RECT 199.800 71.985 200.090 72.030 ;
        RECT 194.790 71.845 200.090 71.985 ;
        RECT 178.815 71.705 178.955 71.845 ;
        RECT 194.790 71.800 195.080 71.845 ;
        RECT 196.680 71.800 196.970 71.845 ;
        RECT 199.800 71.800 200.090 71.845 ;
        RECT 169.985 71.445 170.305 71.705 ;
        RECT 178.725 71.445 179.045 71.705 ;
        RECT 187.465 71.445 187.785 71.705 ;
        RECT 195.745 71.645 196.065 71.705 ;
        RECT 197.585 71.645 197.905 71.705 ;
        RECT 200.435 71.645 200.575 72.185 ;
        RECT 202.645 72.125 202.965 72.185 ;
        RECT 204.025 72.325 204.345 72.385 ;
        RECT 205.955 72.325 206.095 72.480 ;
        RECT 207.245 72.465 207.565 72.525 ;
        RECT 204.025 72.185 206.095 72.325 ;
        RECT 223.435 72.325 223.575 72.525 ;
        RECT 223.820 72.525 230.105 72.665 ;
        RECT 223.820 72.480 224.110 72.525 ;
        RECT 229.785 72.465 230.105 72.525 ;
        RECT 233.465 72.465 233.785 72.725 ;
        RECT 235.765 72.665 236.085 72.725 ;
        RECT 237.605 72.665 237.925 72.725 ;
        RECT 235.765 72.525 237.925 72.665 ;
        RECT 235.765 72.465 236.085 72.525 ;
        RECT 237.605 72.465 237.925 72.525 ;
        RECT 239.905 72.465 240.225 72.725 ;
        RECT 240.460 72.710 240.600 72.865 ;
        RECT 241.300 72.865 256.770 73.005 ;
        RECT 241.300 72.820 241.590 72.865 ;
        RECT 256.480 72.820 256.770 72.865 ;
        RECT 256.940 73.005 257.230 73.050 ;
        RECT 260.605 73.005 260.925 73.065 ;
        RECT 277.165 73.005 277.485 73.065 ;
        RECT 256.940 72.865 277.485 73.005 ;
        RECT 277.715 73.005 277.855 73.205 ;
        RECT 284.525 73.205 294.045 73.345 ;
        RECT 284.525 73.145 284.845 73.205 ;
        RECT 286.365 73.145 286.685 73.205 ;
        RECT 293.725 73.145 294.045 73.205 ;
        RECT 294.660 73.345 294.950 73.390 ;
        RECT 303.860 73.345 304.150 73.390 ;
        RECT 304.305 73.345 304.625 73.405 ;
        RECT 294.660 73.205 296.715 73.345 ;
        RECT 294.660 73.160 294.950 73.205 ;
        RECT 285.445 73.005 285.765 73.065 ;
        RECT 296.025 73.005 296.345 73.065 ;
        RECT 296.575 73.050 296.715 73.205 ;
        RECT 303.860 73.205 304.625 73.345 ;
        RECT 303.860 73.160 304.150 73.205 ;
        RECT 277.715 72.865 285.765 73.005 ;
        RECT 256.940 72.820 257.230 72.865 ;
        RECT 260.605 72.805 260.925 72.865 ;
        RECT 277.165 72.805 277.485 72.865 ;
        RECT 285.445 72.805 285.765 72.865 ;
        RECT 293.815 72.865 296.345 73.005 ;
        RECT 240.385 72.480 240.675 72.710 ;
        RECT 241.745 72.465 242.065 72.725 ;
        RECT 242.665 72.710 242.985 72.725 ;
        RECT 242.450 72.480 242.985 72.710 ;
        RECT 242.665 72.465 242.985 72.480 ;
        RECT 243.125 72.665 243.445 72.725 ;
        RECT 256.005 72.710 256.325 72.725 ;
        RECT 255.100 72.665 255.390 72.710 ;
        RECT 243.125 72.525 255.390 72.665 ;
        RECT 243.125 72.465 243.445 72.525 ;
        RECT 255.100 72.480 255.390 72.525 ;
        RECT 255.840 72.480 256.325 72.710 ;
        RECT 256.005 72.465 256.325 72.480 ;
        RECT 257.385 72.710 257.705 72.725 ;
        RECT 257.385 72.665 257.715 72.710 ;
        RECT 278.085 72.665 278.405 72.725 ;
        RECT 279.020 72.665 279.310 72.710 ;
        RECT 257.385 72.525 257.900 72.665 ;
        RECT 278.085 72.525 279.310 72.665 ;
        RECT 257.385 72.480 257.715 72.525 ;
        RECT 257.385 72.465 257.705 72.480 ;
        RECT 278.085 72.465 278.405 72.525 ;
        RECT 279.020 72.480 279.310 72.525 ;
        RECT 279.465 72.665 279.785 72.725 ;
        RECT 279.940 72.665 280.230 72.710 ;
        RECT 279.465 72.525 280.230 72.665 ;
        RECT 279.465 72.465 279.785 72.525 ;
        RECT 279.940 72.480 280.230 72.525 ;
        RECT 285.905 72.465 286.225 72.725 ;
        RECT 293.815 72.710 293.955 72.865 ;
        RECT 296.025 72.805 296.345 72.865 ;
        RECT 296.500 72.820 296.790 73.050 ;
        RECT 298.780 73.005 299.430 73.050 ;
        RECT 302.380 73.005 302.670 73.050 ;
        RECT 303.385 73.005 303.705 73.065 ;
        RECT 298.780 72.865 303.705 73.005 ;
        RECT 298.780 72.820 299.430 72.865 ;
        RECT 302.080 72.820 302.670 72.865 ;
        RECT 293.740 72.480 294.030 72.710 ;
        RECT 295.585 72.665 295.875 72.710 ;
        RECT 297.420 72.665 297.710 72.710 ;
        RECT 301.000 72.665 301.290 72.710 ;
        RECT 295.585 72.525 301.290 72.665 ;
        RECT 295.585 72.480 295.875 72.525 ;
        RECT 297.420 72.480 297.710 72.525 ;
        RECT 301.000 72.480 301.290 72.525 ;
        RECT 302.080 72.505 302.370 72.820 ;
        RECT 303.385 72.805 303.705 72.865 ;
        RECT 278.545 72.325 278.865 72.385 ;
        RECT 223.435 72.185 278.865 72.325 ;
        RECT 204.025 72.125 204.345 72.185 ;
        RECT 278.545 72.125 278.865 72.185 ;
        RECT 280.385 72.325 280.705 72.385 ;
        RECT 289.600 72.325 289.890 72.370 ;
        RECT 294.185 72.325 294.505 72.385 ;
        RECT 295.120 72.325 295.410 72.370 ;
        RECT 280.385 72.185 295.410 72.325 ;
        RECT 280.385 72.125 280.705 72.185 ;
        RECT 289.600 72.140 289.890 72.185 ;
        RECT 294.185 72.125 294.505 72.185 ;
        RECT 295.120 72.140 295.410 72.185 ;
        RECT 219.205 71.985 219.525 72.045 ;
        RECT 221.505 71.985 221.825 72.045 ;
        RECT 219.205 71.845 221.825 71.985 ;
        RECT 219.205 71.785 219.525 71.845 ;
        RECT 221.505 71.785 221.825 71.845 ;
        RECT 224.725 71.985 225.045 72.045 ;
        RECT 238.525 71.985 238.845 72.045 ;
        RECT 243.585 71.985 243.905 72.045 ;
        RECT 224.725 71.845 243.905 71.985 ;
        RECT 224.725 71.785 225.045 71.845 ;
        RECT 238.525 71.785 238.845 71.845 ;
        RECT 243.585 71.785 243.905 71.845 ;
        RECT 267.045 71.985 267.365 72.045 ;
        RECT 268.425 71.985 268.745 72.045 ;
        RECT 280.860 71.985 281.150 72.030 ;
        RECT 294.645 71.985 294.965 72.045 ;
        RECT 267.045 71.845 280.615 71.985 ;
        RECT 267.045 71.785 267.365 71.845 ;
        RECT 268.425 71.785 268.745 71.845 ;
        RECT 195.745 71.505 200.575 71.645 ;
        RECT 200.805 71.645 201.125 71.705 ;
        RECT 203.580 71.645 203.870 71.690 ;
        RECT 200.805 71.505 203.870 71.645 ;
        RECT 195.745 71.445 196.065 71.505 ;
        RECT 197.585 71.445 197.905 71.505 ;
        RECT 200.805 71.445 201.125 71.505 ;
        RECT 203.580 71.460 203.870 71.505 ;
        RECT 205.420 71.645 205.710 71.690 ;
        RECT 211.845 71.645 212.165 71.705 ;
        RECT 205.420 71.505 212.165 71.645 ;
        RECT 205.420 71.460 205.710 71.505 ;
        RECT 211.845 71.445 212.165 71.505 ;
        RECT 222.420 71.645 222.710 71.690 ;
        RECT 223.805 71.645 224.125 71.705 ;
        RECT 222.420 71.505 224.125 71.645 ;
        RECT 222.420 71.460 222.710 71.505 ;
        RECT 223.805 71.445 224.125 71.505 ;
        RECT 253.245 71.645 253.565 71.705 ;
        RECT 258.765 71.645 259.085 71.705 ;
        RECT 253.245 71.505 259.085 71.645 ;
        RECT 280.475 71.645 280.615 71.845 ;
        RECT 280.860 71.845 294.965 71.985 ;
        RECT 280.860 71.800 281.150 71.845 ;
        RECT 294.645 71.785 294.965 71.845 ;
        RECT 295.990 71.985 296.280 72.030 ;
        RECT 297.880 71.985 298.170 72.030 ;
        RECT 301.000 71.985 301.290 72.030 ;
        RECT 295.990 71.845 301.290 71.985 ;
        RECT 295.990 71.800 296.280 71.845 ;
        RECT 297.880 71.800 298.170 71.845 ;
        RECT 301.000 71.800 301.290 71.845 ;
        RECT 303.935 71.645 304.075 73.160 ;
        RECT 304.305 73.145 304.625 73.205 ;
        RECT 280.475 71.505 304.075 71.645 ;
        RECT 253.245 71.445 253.565 71.505 ;
        RECT 258.765 71.445 259.085 71.505 ;
        RECT 162.095 70.825 311.135 71.305 ;
        RECT 174.140 70.625 174.430 70.670 ;
        RECT 175.505 70.625 175.825 70.685 ;
        RECT 174.140 70.485 175.825 70.625 ;
        RECT 174.140 70.440 174.430 70.485 ;
        RECT 175.505 70.425 175.825 70.485 ;
        RECT 194.380 70.625 194.670 70.670 ;
        RECT 196.205 70.625 196.525 70.685 ;
        RECT 194.380 70.485 196.525 70.625 ;
        RECT 194.380 70.440 194.670 70.485 ;
        RECT 196.205 70.425 196.525 70.485 ;
        RECT 201.725 70.625 202.045 70.685 ;
        RECT 215.985 70.625 216.305 70.685 ;
        RECT 232.560 70.625 232.850 70.670 ;
        RECT 236.225 70.625 236.545 70.685 ;
        RECT 201.725 70.485 220.815 70.625 ;
        RECT 201.725 70.425 202.045 70.485 ;
        RECT 215.985 70.425 216.305 70.485 ;
        RECT 166.270 70.285 166.560 70.330 ;
        RECT 168.160 70.285 168.450 70.330 ;
        RECT 171.280 70.285 171.570 70.330 ;
        RECT 166.270 70.145 171.570 70.285 ;
        RECT 166.270 70.100 166.560 70.145 ;
        RECT 168.160 70.100 168.450 70.145 ;
        RECT 171.280 70.100 171.570 70.145 ;
        RECT 187.925 70.285 188.245 70.345 ;
        RECT 188.400 70.285 188.690 70.330 ;
        RECT 201.265 70.285 201.585 70.345 ;
        RECT 208.165 70.285 208.485 70.345 ;
        RECT 187.925 70.145 188.690 70.285 ;
        RECT 187.925 70.085 188.245 70.145 ;
        RECT 188.400 70.100 188.690 70.145 ;
        RECT 188.935 70.145 197.355 70.285 ;
        RECT 166.780 69.945 167.070 69.990 ;
        RECT 169.985 69.945 170.305 70.005 ;
        RECT 166.780 69.805 170.305 69.945 ;
        RECT 166.780 69.760 167.070 69.805 ;
        RECT 169.985 69.745 170.305 69.805 ;
        RECT 176.425 69.945 176.745 70.005 ;
        RECT 179.185 69.945 179.505 70.005 ;
        RECT 179.660 69.945 179.950 69.990 ;
        RECT 183.325 69.945 183.645 70.005 ;
        RECT 188.935 69.945 189.075 70.145 ;
        RECT 176.425 69.805 183.645 69.945 ;
        RECT 176.425 69.745 176.745 69.805 ;
        RECT 179.185 69.745 179.505 69.805 ;
        RECT 179.660 69.760 179.950 69.805 ;
        RECT 183.325 69.745 183.645 69.805 ;
        RECT 187.095 69.805 189.075 69.945 ;
        RECT 165.385 69.405 165.705 69.665 ;
        RECT 165.865 69.605 166.155 69.650 ;
        RECT 167.700 69.605 167.990 69.650 ;
        RECT 171.280 69.605 171.570 69.650 ;
        RECT 165.865 69.465 171.570 69.605 ;
        RECT 165.865 69.420 166.155 69.465 ;
        RECT 167.700 69.420 167.990 69.465 ;
        RECT 171.280 69.420 171.570 69.465 ;
        RECT 172.285 69.625 172.605 69.665 ;
        RECT 172.285 69.405 172.650 69.625 ;
        RECT 187.095 69.605 187.235 69.805 ;
        RECT 192.540 69.760 192.830 69.990 ;
        RECT 193.445 69.945 193.765 70.005 ;
        RECT 196.665 69.945 196.985 70.005 ;
        RECT 193.445 69.805 196.985 69.945 ;
        RECT 172.360 69.310 172.650 69.405 ;
        RECT 178.355 69.465 187.235 69.605 ;
        RECT 187.465 69.605 187.785 69.665 ;
        RECT 189.320 69.605 189.610 69.650 ;
        RECT 187.465 69.465 189.610 69.605 ;
        RECT 169.060 69.265 169.710 69.310 ;
        RECT 172.360 69.265 172.950 69.310 ;
        RECT 177.345 69.265 177.665 69.325 ;
        RECT 178.355 69.310 178.495 69.465 ;
        RECT 187.465 69.405 187.785 69.465 ;
        RECT 189.320 69.420 189.610 69.465 ;
        RECT 192.065 69.405 192.385 69.665 ;
        RECT 178.280 69.265 178.570 69.310 ;
        RECT 169.060 69.125 172.950 69.265 ;
        RECT 169.060 69.080 169.710 69.125 ;
        RECT 172.660 69.080 172.950 69.125 ;
        RECT 173.755 69.125 176.655 69.265 ;
        RECT 171.365 68.925 171.685 68.985 ;
        RECT 173.755 68.925 173.895 69.125 ;
        RECT 176.515 68.970 176.655 69.125 ;
        RECT 177.345 69.125 178.570 69.265 ;
        RECT 177.345 69.065 177.665 69.125 ;
        RECT 178.280 69.080 178.570 69.125 ;
        RECT 179.185 69.265 179.505 69.325 ;
        RECT 192.615 69.265 192.755 69.760 ;
        RECT 193.445 69.745 193.765 69.805 ;
        RECT 196.665 69.745 196.985 69.805 ;
        RECT 195.285 69.650 195.605 69.665 ;
        RECT 195.265 69.420 195.605 69.650 ;
        RECT 197.215 69.605 197.355 70.145 ;
        RECT 201.265 70.145 208.485 70.285 ;
        RECT 201.265 70.085 201.585 70.145 ;
        RECT 208.165 70.085 208.485 70.145 ;
        RECT 208.625 70.285 208.945 70.345 ;
        RECT 210.465 70.285 210.785 70.345 ;
        RECT 208.625 70.145 210.785 70.285 ;
        RECT 220.675 70.285 220.815 70.485 ;
        RECT 222.055 70.485 227.255 70.625 ;
        RECT 222.055 70.285 222.195 70.485 ;
        RECT 220.675 70.145 222.195 70.285 ;
        RECT 223.805 70.285 224.125 70.345 ;
        RECT 226.565 70.285 226.885 70.345 ;
        RECT 223.805 70.145 226.885 70.285 ;
        RECT 227.115 70.285 227.255 70.485 ;
        RECT 232.560 70.485 236.545 70.625 ;
        RECT 232.560 70.440 232.850 70.485 ;
        RECT 236.225 70.425 236.545 70.485 ;
        RECT 237.160 70.625 237.450 70.670 ;
        RECT 239.905 70.625 240.225 70.685 ;
        RECT 237.160 70.485 240.225 70.625 ;
        RECT 237.160 70.440 237.450 70.485 ;
        RECT 239.905 70.425 240.225 70.485 ;
        RECT 240.365 70.625 240.685 70.685 ;
        RECT 257.845 70.625 258.165 70.685 ;
        RECT 240.365 70.485 258.165 70.625 ;
        RECT 240.365 70.425 240.685 70.485 ;
        RECT 257.845 70.425 258.165 70.485 ;
        RECT 258.305 70.625 258.625 70.685 ;
        RECT 276.705 70.625 277.025 70.685 ;
        RECT 258.305 70.485 277.025 70.625 ;
        RECT 258.305 70.425 258.625 70.485 ;
        RECT 276.705 70.425 277.025 70.485 ;
        RECT 279.020 70.625 279.310 70.670 ;
        RECT 279.925 70.625 280.245 70.685 ;
        RECT 279.020 70.485 280.245 70.625 ;
        RECT 279.020 70.440 279.310 70.485 ;
        RECT 261.065 70.285 261.385 70.345 ;
        RECT 279.095 70.285 279.235 70.440 ;
        RECT 279.925 70.425 280.245 70.485 ;
        RECT 284.985 70.625 285.305 70.685 ;
        RECT 286.840 70.625 287.130 70.670 ;
        RECT 284.985 70.485 287.130 70.625 ;
        RECT 284.985 70.425 285.305 70.485 ;
        RECT 286.840 70.440 287.130 70.485 ;
        RECT 288.205 70.625 288.525 70.685 ;
        RECT 301.085 70.625 301.405 70.685 ;
        RECT 288.205 70.485 301.405 70.625 ;
        RECT 288.205 70.425 288.525 70.485 ;
        RECT 301.085 70.425 301.405 70.485 ;
        RECT 302.940 70.625 303.230 70.670 ;
        RECT 304.765 70.625 305.085 70.685 ;
        RECT 302.940 70.485 305.085 70.625 ;
        RECT 302.940 70.440 303.230 70.485 ;
        RECT 304.765 70.425 305.085 70.485 ;
        RECT 282.700 70.285 282.990 70.330 ;
        RECT 227.115 70.145 260.835 70.285 ;
        RECT 208.625 70.085 208.945 70.145 ;
        RECT 210.465 70.085 210.785 70.145 ;
        RECT 223.805 70.085 224.125 70.145 ;
        RECT 226.565 70.085 226.885 70.145 ;
        RECT 197.585 69.745 197.905 70.005 ;
        RECT 202.185 69.945 202.505 70.005 ;
        RECT 209.085 69.945 209.405 70.005 ;
        RECT 221.965 69.945 222.285 70.005 ;
        RECT 202.185 69.805 204.715 69.945 ;
        RECT 202.185 69.745 202.505 69.805 ;
        RECT 201.725 69.605 202.045 69.665 ;
        RECT 197.215 69.585 198.275 69.605 ;
        RECT 198.595 69.585 202.045 69.605 ;
        RECT 197.215 69.465 202.045 69.585 ;
        RECT 195.285 69.405 195.605 69.420 ;
        RECT 198.135 69.445 198.735 69.465 ;
        RECT 197.125 69.265 197.445 69.325 ;
        RECT 179.185 69.125 197.445 69.265 ;
        RECT 179.185 69.065 179.505 69.125 ;
        RECT 197.125 69.065 197.445 69.125 ;
        RECT 171.365 68.785 173.895 68.925 ;
        RECT 171.365 68.725 171.685 68.785 ;
        RECT 176.440 68.740 176.730 68.970 ;
        RECT 178.740 68.925 179.030 68.970 ;
        RECT 180.565 68.925 180.885 68.985 ;
        RECT 178.740 68.785 180.885 68.925 ;
        RECT 178.740 68.740 179.030 68.785 ;
        RECT 180.565 68.725 180.885 68.785 ;
        RECT 189.765 68.725 190.085 68.985 ;
        RECT 191.620 68.925 191.910 68.970 ;
        RECT 196.665 68.925 196.985 68.985 ;
        RECT 198.135 68.970 198.275 69.445 ;
        RECT 201.725 69.405 202.045 69.465 ;
        RECT 203.565 69.405 203.885 69.665 ;
        RECT 204.025 69.405 204.345 69.665 ;
        RECT 203.120 69.080 203.410 69.310 ;
        RECT 204.575 69.265 204.715 69.805 ;
        RECT 205.035 69.805 212.995 69.945 ;
        RECT 205.035 69.650 205.175 69.805 ;
        RECT 209.085 69.745 209.405 69.805 ;
        RECT 204.960 69.420 205.250 69.650 ;
        RECT 206.800 69.605 207.090 69.650 ;
        RECT 205.495 69.465 207.090 69.605 ;
        RECT 205.495 69.265 205.635 69.465 ;
        RECT 206.800 69.420 207.090 69.465 ;
        RECT 207.245 69.405 207.565 69.665 ;
        RECT 208.180 69.605 208.470 69.650 ;
        RECT 209.545 69.605 209.865 69.665 ;
        RECT 212.855 69.650 212.995 69.805 ;
        RECT 221.965 69.805 227.720 69.945 ;
        RECT 221.965 69.745 222.285 69.805 ;
        RECT 208.180 69.465 209.865 69.605 ;
        RECT 208.180 69.420 208.470 69.465 ;
        RECT 209.545 69.405 209.865 69.465 ;
        RECT 212.780 69.420 213.070 69.650 ;
        RECT 224.265 69.605 224.585 69.665 ;
        RECT 226.565 69.605 226.885 69.665 ;
        RECT 227.580 69.650 227.720 69.805 ;
        RECT 228.955 69.805 235.075 69.945 ;
        RECT 228.955 69.650 229.095 69.805 ;
        RECT 234.935 69.665 235.075 69.805 ;
        RECT 235.765 69.745 236.085 70.005 ;
        RECT 247.265 69.945 247.585 70.005 ;
        RECT 236.440 69.805 247.585 69.945 ;
        RECT 236.440 69.665 236.580 69.805 ;
        RECT 247.265 69.745 247.585 69.805 ;
        RECT 251.865 69.945 252.185 70.005 ;
        RECT 257.400 69.945 257.690 69.990 ;
        RECT 259.685 69.945 260.005 70.005 ;
        RECT 251.865 69.805 255.340 69.945 ;
        RECT 251.865 69.745 252.185 69.805 ;
        RECT 227.040 69.605 227.330 69.650 ;
        RECT 224.265 69.465 227.330 69.605 ;
        RECT 224.265 69.405 224.585 69.465 ;
        RECT 226.565 69.405 226.885 69.465 ;
        RECT 227.040 69.420 227.330 69.465 ;
        RECT 227.505 69.420 227.795 69.650 ;
        RECT 228.880 69.420 229.170 69.650 ;
        RECT 229.570 69.605 229.860 69.650 ;
        RECT 230.705 69.605 231.025 69.665 ;
        RECT 229.570 69.465 231.025 69.605 ;
        RECT 229.570 69.420 229.860 69.465 ;
        RECT 230.705 69.405 231.025 69.465 ;
        RECT 232.085 69.605 232.405 69.665 ;
        RECT 233.925 69.605 234.245 69.665 ;
        RECT 232.085 69.465 234.245 69.605 ;
        RECT 232.085 69.405 232.405 69.465 ;
        RECT 233.925 69.405 234.245 69.465 ;
        RECT 234.845 69.405 235.165 69.665 ;
        RECT 236.225 69.650 236.580 69.665 ;
        RECT 236.225 69.420 236.655 69.650 ;
        RECT 238.065 69.605 238.385 69.665 ;
        RECT 245.900 69.605 246.190 69.650 ;
        RECT 252.800 69.605 253.090 69.650 ;
        RECT 238.065 69.465 244.735 69.605 ;
        RECT 236.225 69.405 236.545 69.420 ;
        RECT 238.065 69.405 238.385 69.465 ;
        RECT 244.595 69.325 244.735 69.465 ;
        RECT 245.900 69.465 253.090 69.605 ;
        RECT 245.900 69.420 246.190 69.465 ;
        RECT 252.800 69.420 253.090 69.465 ;
        RECT 253.245 69.605 253.565 69.665 ;
        RECT 253.245 69.465 253.760 69.605 ;
        RECT 253.245 69.405 253.565 69.465 ;
        RECT 254.625 69.405 254.945 69.665 ;
        RECT 255.200 69.650 255.340 69.805 ;
        RECT 257.400 69.805 260.005 69.945 ;
        RECT 257.400 69.760 257.690 69.805 ;
        RECT 259.685 69.745 260.005 69.805 ;
        RECT 255.125 69.585 255.415 69.650 ;
        RECT 257.845 69.605 258.165 69.665 ;
        RECT 255.865 69.585 258.165 69.605 ;
        RECT 255.125 69.465 258.165 69.585 ;
        RECT 255.125 69.445 256.005 69.465 ;
        RECT 255.125 69.420 255.415 69.445 ;
        RECT 257.845 69.405 258.165 69.465 ;
        RECT 258.320 69.420 258.610 69.650 ;
        RECT 204.575 69.125 205.635 69.265 ;
        RECT 206.340 69.080 206.630 69.310 ;
        RECT 207.705 69.265 208.025 69.325 ;
        RECT 210.020 69.265 210.310 69.310 ;
        RECT 207.705 69.125 210.310 69.265 ;
        RECT 191.620 68.785 196.985 68.925 ;
        RECT 191.620 68.740 191.910 68.785 ;
        RECT 196.665 68.725 196.985 68.785 ;
        RECT 198.060 68.740 198.350 68.970 ;
        RECT 199.885 68.725 200.205 68.985 ;
        RECT 203.195 68.925 203.335 69.080 ;
        RECT 205.405 68.925 205.725 68.985 ;
        RECT 206.415 68.925 206.555 69.080 ;
        RECT 207.705 69.065 208.025 69.125 ;
        RECT 210.020 69.080 210.310 69.125 ;
        RECT 211.845 69.265 212.165 69.325 ;
        RECT 228.420 69.265 228.710 69.310 ;
        RECT 232.545 69.265 232.865 69.325 ;
        RECT 235.320 69.265 235.610 69.310 ;
        RECT 241.285 69.265 241.605 69.325 ;
        RECT 211.845 69.125 230.935 69.265 ;
        RECT 211.845 69.065 212.165 69.125 ;
        RECT 228.420 69.080 228.710 69.125 ;
        RECT 203.195 68.785 206.555 68.925 ;
        RECT 213.240 68.925 213.530 68.970 ;
        RECT 229.785 68.925 230.105 68.985 ;
        RECT 213.240 68.785 230.105 68.925 ;
        RECT 205.405 68.725 205.725 68.785 ;
        RECT 213.240 68.740 213.530 68.785 ;
        RECT 229.785 68.725 230.105 68.785 ;
        RECT 230.245 68.725 230.565 68.985 ;
        RECT 230.795 68.925 230.935 69.125 ;
        RECT 232.545 69.125 241.605 69.265 ;
        RECT 232.545 69.065 232.865 69.125 ;
        RECT 235.320 69.080 235.610 69.125 ;
        RECT 241.285 69.065 241.605 69.125 ;
        RECT 243.140 69.265 243.430 69.310 ;
        RECT 243.585 69.265 243.905 69.325 ;
        RECT 243.140 69.125 243.905 69.265 ;
        RECT 243.140 69.080 243.430 69.125 ;
        RECT 243.585 69.065 243.905 69.125 ;
        RECT 244.505 69.065 244.825 69.325 ;
        RECT 244.980 69.265 245.270 69.310 ;
        RECT 248.185 69.265 248.505 69.325 ;
        RECT 254.180 69.265 254.470 69.310 ;
        RECT 258.395 69.265 258.535 69.420 ;
        RECT 244.980 69.125 247.955 69.265 ;
        RECT 244.980 69.080 245.270 69.125 ;
        RECT 238.065 68.925 238.385 68.985 ;
        RECT 230.795 68.785 238.385 68.925 ;
        RECT 238.065 68.725 238.385 68.785 ;
        RECT 238.985 68.925 239.305 68.985 ;
        RECT 244.060 68.925 244.350 68.970 ;
        RECT 246.345 68.925 246.665 68.985 ;
        RECT 238.985 68.785 246.665 68.925 ;
        RECT 247.815 68.925 247.955 69.125 ;
        RECT 248.185 69.125 258.535 69.265 ;
        RECT 260.695 69.265 260.835 70.145 ;
        RECT 261.065 70.145 279.235 70.285 ;
        RECT 280.475 70.145 282.990 70.285 ;
        RECT 261.065 70.085 261.385 70.145 ;
        RECT 263.365 69.945 263.685 70.005 ;
        RECT 268.885 69.945 269.205 70.005 ;
        RECT 274.880 69.945 275.170 69.990 ;
        RECT 263.365 69.805 275.170 69.945 ;
        RECT 263.365 69.745 263.685 69.805 ;
        RECT 268.885 69.745 269.205 69.805 ;
        RECT 274.880 69.760 275.170 69.805 ;
        RECT 275.325 69.745 275.645 70.005 ;
        RECT 278.545 69.405 278.865 69.665 ;
        RECT 279.465 69.605 279.785 69.665 ;
        RECT 279.940 69.605 280.230 69.650 ;
        RECT 279.465 69.465 280.230 69.605 ;
        RECT 280.475 69.605 280.615 70.145 ;
        RECT 282.700 70.100 282.990 70.145 ;
        RECT 295.070 70.285 295.360 70.330 ;
        RECT 296.960 70.285 297.250 70.330 ;
        RECT 300.080 70.285 300.370 70.330 ;
        RECT 295.070 70.145 300.370 70.285 ;
        RECT 295.070 70.100 295.360 70.145 ;
        RECT 296.960 70.100 297.250 70.145 ;
        RECT 300.080 70.100 300.370 70.145 ;
        RECT 303.845 70.285 304.165 70.345 ;
        RECT 305.240 70.285 305.530 70.330 ;
        RECT 303.845 70.145 305.530 70.285 ;
        RECT 303.845 70.085 304.165 70.145 ;
        RECT 305.240 70.100 305.530 70.145 ;
        RECT 280.860 69.945 281.150 69.990 ;
        RECT 285.920 69.945 286.210 69.990 ;
        RECT 290.045 69.945 290.365 70.005 ;
        RECT 280.860 69.805 290.365 69.945 ;
        RECT 280.860 69.760 281.150 69.805 ;
        RECT 285.920 69.760 286.210 69.805 ;
        RECT 290.045 69.745 290.365 69.805 ;
        RECT 294.185 69.745 294.505 70.005 ;
        RECT 295.580 69.945 295.870 69.990 ;
        RECT 298.325 69.945 298.645 70.005 ;
        RECT 310.745 69.945 311.065 70.005 ;
        RECT 295.580 69.805 298.645 69.945 ;
        RECT 295.580 69.760 295.870 69.805 ;
        RECT 298.325 69.745 298.645 69.805 ;
        RECT 309.455 69.805 311.065 69.945 ;
        RECT 282.240 69.605 282.530 69.650 ;
        RECT 280.475 69.465 282.530 69.605 ;
        RECT 279.465 69.405 279.785 69.465 ;
        RECT 279.940 69.420 280.230 69.465 ;
        RECT 282.240 69.420 282.530 69.465 ;
        RECT 284.525 69.405 284.845 69.665 ;
        RECT 288.665 69.405 288.985 69.665 ;
        RECT 294.665 69.605 294.955 69.650 ;
        RECT 296.500 69.605 296.790 69.650 ;
        RECT 300.080 69.605 300.370 69.650 ;
        RECT 294.665 69.465 300.370 69.605 ;
        RECT 294.665 69.420 294.955 69.465 ;
        RECT 296.500 69.420 296.790 69.465 ;
        RECT 300.080 69.420 300.370 69.465 ;
        RECT 301.160 69.605 301.450 69.625 ;
        RECT 303.385 69.605 303.705 69.665 ;
        RECT 301.160 69.465 303.705 69.605 ;
        RECT 301.160 69.310 301.450 69.465 ;
        RECT 303.385 69.405 303.705 69.465 ;
        RECT 304.305 69.405 304.625 69.665 ;
        RECT 309.455 69.650 309.595 69.805 ;
        RECT 310.745 69.745 311.065 69.805 ;
        RECT 309.380 69.420 309.670 69.650 ;
        RECT 274.420 69.265 274.710 69.310 ;
        RECT 297.860 69.265 298.510 69.310 ;
        RECT 301.160 69.265 301.750 69.310 ;
        RECT 260.695 69.125 289.355 69.265 ;
        RECT 248.185 69.065 248.505 69.125 ;
        RECT 254.180 69.080 254.470 69.125 ;
        RECT 274.420 69.080 274.710 69.125 ;
        RECT 250.945 68.925 251.265 68.985 ;
        RECT 247.815 68.785 251.265 68.925 ;
        RECT 238.985 68.725 239.305 68.785 ;
        RECT 244.060 68.740 244.350 68.785 ;
        RECT 246.345 68.725 246.665 68.785 ;
        RECT 250.945 68.725 251.265 68.785 ;
        RECT 253.245 68.925 253.565 68.985 ;
        RECT 256.020 68.925 256.310 68.970 ;
        RECT 253.245 68.785 256.310 68.925 ;
        RECT 253.245 68.725 253.565 68.785 ;
        RECT 256.020 68.740 256.310 68.785 ;
        RECT 259.225 68.725 259.545 68.985 ;
        RECT 269.805 68.925 270.125 68.985 ;
        RECT 272.580 68.925 272.870 68.970 ;
        RECT 269.805 68.785 272.870 68.925 ;
        RECT 269.805 68.725 270.125 68.785 ;
        RECT 272.580 68.740 272.870 68.785 ;
        RECT 281.305 68.725 281.625 68.985 ;
        RECT 285.000 68.925 285.290 68.970 ;
        RECT 288.205 68.925 288.525 68.985 ;
        RECT 289.215 68.970 289.355 69.125 ;
        RECT 297.860 69.125 301.750 69.265 ;
        RECT 297.860 69.080 298.510 69.125 ;
        RECT 301.460 69.080 301.750 69.125 ;
        RECT 285.000 68.785 288.525 68.925 ;
        RECT 285.000 68.740 285.290 68.785 ;
        RECT 288.205 68.725 288.525 68.785 ;
        RECT 289.140 68.925 289.430 68.970 ;
        RECT 297.405 68.925 297.725 68.985 ;
        RECT 289.140 68.785 297.725 68.925 ;
        RECT 289.140 68.740 289.430 68.785 ;
        RECT 297.405 68.725 297.725 68.785 ;
        RECT 305.685 68.925 306.005 68.985 ;
        RECT 308.460 68.925 308.750 68.970 ;
        RECT 305.685 68.785 308.750 68.925 ;
        RECT 305.685 68.725 306.005 68.785 ;
        RECT 308.460 68.740 308.750 68.785 ;
        RECT 162.095 68.105 311.935 68.585 ;
        RECT 171.380 67.720 171.670 67.950 ;
        RECT 172.285 67.905 172.605 67.965 ;
        RECT 198.060 67.905 198.350 67.950 ;
        RECT 172.285 67.765 175.275 67.905 ;
        RECT 171.455 67.565 171.595 67.720 ;
        RECT 172.285 67.705 172.605 67.765 ;
        RECT 173.220 67.565 173.510 67.610 ;
        RECT 171.455 67.425 173.510 67.565 ;
        RECT 175.135 67.565 175.275 67.765 ;
        RECT 185.255 67.765 198.350 67.905 ;
        RECT 175.500 67.565 176.150 67.610 ;
        RECT 179.100 67.565 179.390 67.610 ;
        RECT 175.135 67.425 179.390 67.565 ;
        RECT 173.220 67.380 173.510 67.425 ;
        RECT 175.500 67.380 176.150 67.425 ;
        RECT 178.800 67.380 179.390 67.425 ;
        RECT 169.985 67.025 170.305 67.285 ;
        RECT 170.460 67.225 170.750 67.270 ;
        RECT 171.365 67.225 171.685 67.285 ;
        RECT 170.460 67.085 171.685 67.225 ;
        RECT 170.460 67.040 170.750 67.085 ;
        RECT 171.365 67.025 171.685 67.085 ;
        RECT 172.305 67.225 172.595 67.270 ;
        RECT 174.140 67.225 174.430 67.270 ;
        RECT 177.720 67.225 178.010 67.270 ;
        RECT 172.305 67.085 178.010 67.225 ;
        RECT 172.305 67.040 172.595 67.085 ;
        RECT 174.140 67.040 174.430 67.085 ;
        RECT 177.720 67.040 178.010 67.085 ;
        RECT 178.800 67.065 179.090 67.380 ;
        RECT 185.255 67.270 185.395 67.765 ;
        RECT 198.060 67.720 198.350 67.765 ;
        RECT 199.900 67.905 200.190 67.950 ;
        RECT 200.345 67.905 200.665 67.965 ;
        RECT 199.900 67.765 200.665 67.905 ;
        RECT 199.900 67.720 200.190 67.765 ;
        RECT 200.345 67.705 200.665 67.765 ;
        RECT 202.645 67.905 202.965 67.965 ;
        RECT 204.025 67.905 204.345 67.965 ;
        RECT 202.645 67.765 204.345 67.905 ;
        RECT 202.645 67.705 202.965 67.765 ;
        RECT 204.025 67.705 204.345 67.765 ;
        RECT 208.180 67.905 208.470 67.950 ;
        RECT 209.085 67.905 209.405 67.965 ;
        RECT 208.180 67.765 209.405 67.905 ;
        RECT 208.180 67.720 208.470 67.765 ;
        RECT 209.085 67.705 209.405 67.765 ;
        RECT 209.545 67.905 209.865 67.965 ;
        RECT 211.860 67.905 212.150 67.950 ;
        RECT 209.545 67.765 212.150 67.905 ;
        RECT 209.545 67.705 209.865 67.765 ;
        RECT 211.860 67.720 212.150 67.765 ;
        RECT 216.000 67.905 216.290 67.950 ;
        RECT 224.740 67.905 225.030 67.950 ;
        RECT 225.185 67.905 225.505 67.965 ;
        RECT 216.000 67.765 224.500 67.905 ;
        RECT 216.000 67.720 216.290 67.765 ;
        RECT 189.765 67.565 190.085 67.625 ;
        RECT 186.635 67.425 190.085 67.565 ;
        RECT 186.635 67.270 186.775 67.425 ;
        RECT 189.765 67.365 190.085 67.425 ;
        RECT 192.060 67.565 192.710 67.610 ;
        RECT 195.660 67.565 195.950 67.610 ;
        RECT 196.205 67.565 196.525 67.625 ;
        RECT 192.060 67.425 196.525 67.565 ;
        RECT 192.060 67.380 192.710 67.425 ;
        RECT 195.360 67.380 195.950 67.425 ;
        RECT 185.180 67.040 185.470 67.270 ;
        RECT 186.560 67.040 186.850 67.270 ;
        RECT 188.865 67.225 189.155 67.270 ;
        RECT 190.700 67.225 190.990 67.270 ;
        RECT 194.280 67.225 194.570 67.270 ;
        RECT 188.865 67.085 194.570 67.225 ;
        RECT 188.865 67.040 189.155 67.085 ;
        RECT 190.700 67.040 190.990 67.085 ;
        RECT 194.280 67.040 194.570 67.085 ;
        RECT 195.360 67.065 195.650 67.380 ;
        RECT 196.205 67.365 196.525 67.425 ;
        RECT 197.125 67.565 197.445 67.625 ;
        RECT 200.805 67.565 201.125 67.625 ;
        RECT 197.125 67.425 201.125 67.565 ;
        RECT 197.125 67.365 197.445 67.425 ;
        RECT 200.805 67.365 201.125 67.425 ;
        RECT 201.265 67.565 201.585 67.625 ;
        RECT 210.005 67.565 210.325 67.625 ;
        RECT 201.265 67.425 210.325 67.565 ;
        RECT 201.265 67.365 201.585 67.425 ;
        RECT 210.005 67.365 210.325 67.425 ;
        RECT 171.840 66.885 172.130 66.930 ;
        RECT 181.945 66.885 182.265 66.945 ;
        RECT 186.085 66.885 186.405 66.945 ;
        RECT 188.400 66.885 188.690 66.930 ;
        RECT 189.780 66.885 190.070 66.930 ;
        RECT 171.840 66.745 188.690 66.885 ;
        RECT 171.840 66.700 172.130 66.745 ;
        RECT 165.385 66.545 165.705 66.605 ;
        RECT 171.915 66.545 172.055 66.700 ;
        RECT 181.945 66.685 182.265 66.745 ;
        RECT 186.085 66.685 186.405 66.745 ;
        RECT 188.400 66.700 188.690 66.745 ;
        RECT 188.935 66.745 190.070 66.885 ;
        RECT 165.385 66.405 172.055 66.545 ;
        RECT 172.710 66.545 173.000 66.590 ;
        RECT 174.600 66.545 174.890 66.590 ;
        RECT 177.720 66.545 178.010 66.590 ;
        RECT 172.710 66.405 178.010 66.545 ;
        RECT 165.385 66.345 165.705 66.405 ;
        RECT 172.710 66.360 173.000 66.405 ;
        RECT 174.600 66.360 174.890 66.405 ;
        RECT 177.720 66.360 178.010 66.405 ;
        RECT 180.565 66.345 180.885 66.605 ;
        RECT 188.935 66.545 189.075 66.745 ;
        RECT 189.780 66.700 190.070 66.745 ;
        RECT 197.140 66.885 197.430 66.930 ;
        RECT 199.885 66.885 200.205 66.945 ;
        RECT 197.140 66.745 200.205 66.885 ;
        RECT 197.140 66.700 197.430 66.745 ;
        RECT 199.885 66.685 200.205 66.745 ;
        RECT 200.345 66.685 200.665 66.945 ;
        RECT 200.895 66.930 201.035 67.365 ;
        RECT 204.025 67.225 204.345 67.285 ;
        RECT 204.500 67.225 204.790 67.270 ;
        RECT 204.025 67.085 204.790 67.225 ;
        RECT 204.025 67.025 204.345 67.085 ;
        RECT 204.500 67.040 204.790 67.085 ;
        RECT 207.245 67.025 207.565 67.285 ;
        RECT 208.165 67.025 208.485 67.285 ;
        RECT 209.085 67.025 209.405 67.285 ;
        RECT 210.925 67.025 211.245 67.285 ;
        RECT 211.935 67.225 212.075 67.720 ;
        RECT 223.345 67.565 223.665 67.625 ;
        RECT 213.315 67.425 223.665 67.565 ;
        RECT 224.360 67.565 224.500 67.765 ;
        RECT 224.740 67.765 225.505 67.905 ;
        RECT 224.740 67.720 225.030 67.765 ;
        RECT 225.185 67.705 225.505 67.765 ;
        RECT 226.105 67.705 226.425 67.965 ;
        RECT 227.960 67.720 228.250 67.950 ;
        RECT 229.785 67.905 230.105 67.965 ;
        RECT 236.685 67.905 237.005 67.965 ;
        RECT 240.825 67.905 241.145 67.965 ;
        RECT 257.845 67.905 258.165 67.965 ;
        RECT 229.785 67.765 249.105 67.905 ;
        RECT 226.195 67.565 226.335 67.705 ;
        RECT 228.035 67.565 228.175 67.720 ;
        RECT 229.785 67.705 230.105 67.765 ;
        RECT 236.685 67.705 237.005 67.765 ;
        RECT 240.825 67.705 241.145 67.765 ;
        RECT 239.905 67.565 240.225 67.625 ;
        RECT 224.360 67.425 227.255 67.565 ;
        RECT 228.035 67.425 230.475 67.565 ;
        RECT 212.305 67.225 212.625 67.285 ;
        RECT 213.315 67.270 213.455 67.425 ;
        RECT 223.345 67.365 223.665 67.425 ;
        RECT 211.935 67.085 212.625 67.225 ;
        RECT 212.305 67.025 212.625 67.085 ;
        RECT 213.240 67.040 213.530 67.270 ;
        RECT 200.820 66.700 201.110 66.930 ;
        RECT 204.945 66.885 205.265 66.945 ;
        RECT 205.865 66.885 206.185 66.945 ;
        RECT 213.315 66.885 213.455 67.040 ;
        RECT 214.605 67.025 214.925 67.285 ;
        RECT 221.965 67.225 222.285 67.285 ;
        RECT 223.820 67.225 224.110 67.270 ;
        RECT 221.965 67.085 224.110 67.225 ;
        RECT 221.965 67.025 222.285 67.085 ;
        RECT 223.820 67.040 224.110 67.085 ;
        RECT 224.725 67.025 225.045 67.285 ;
        RECT 225.200 67.225 225.490 67.270 ;
        RECT 225.645 67.225 225.965 67.285 ;
        RECT 227.115 67.270 227.255 67.425 ;
        RECT 225.200 67.085 225.965 67.225 ;
        RECT 225.200 67.040 225.490 67.085 ;
        RECT 225.645 67.025 225.965 67.085 ;
        RECT 226.120 67.040 226.410 67.270 ;
        RECT 226.580 67.040 226.870 67.270 ;
        RECT 227.040 67.040 227.330 67.270 ;
        RECT 204.945 66.745 213.455 66.885 ;
        RECT 221.505 66.885 221.825 66.945 ;
        RECT 222.885 66.885 223.205 66.945 ;
        RECT 221.505 66.745 223.205 66.885 ;
        RECT 204.945 66.685 205.265 66.745 ;
        RECT 205.865 66.685 206.185 66.745 ;
        RECT 221.505 66.685 221.825 66.745 ;
        RECT 222.885 66.685 223.205 66.745 ;
        RECT 223.360 66.885 223.650 66.930 ;
        RECT 224.815 66.885 224.955 67.025 ;
        RECT 226.195 66.885 226.335 67.040 ;
        RECT 223.360 66.745 224.035 66.885 ;
        RECT 224.815 66.745 226.335 66.885 ;
        RECT 226.655 66.885 226.795 67.040 ;
        RECT 228.405 67.025 228.725 67.285 ;
        RECT 229.325 67.025 229.645 67.285 ;
        RECT 230.335 67.270 230.475 67.425 ;
        RECT 236.315 67.425 240.225 67.565 ;
        RECT 248.965 67.565 249.105 67.765 ;
        RECT 257.845 67.765 260.375 67.905 ;
        RECT 257.845 67.705 258.165 67.765 ;
        RECT 255.560 67.565 255.850 67.610 ;
        RECT 248.965 67.425 255.850 67.565 ;
        RECT 236.315 67.285 236.455 67.425 ;
        RECT 239.905 67.365 240.225 67.425 ;
        RECT 255.560 67.380 255.850 67.425 ;
        RECT 256.005 67.365 256.325 67.625 ;
        RECT 258.305 67.565 258.625 67.625 ;
        RECT 259.700 67.565 259.990 67.610 ;
        RECT 258.305 67.425 259.990 67.565 ;
        RECT 258.305 67.365 258.625 67.425 ;
        RECT 259.700 67.380 259.990 67.425 ;
        RECT 260.235 67.285 260.375 67.765 ;
        RECT 260.605 67.705 260.925 67.965 ;
        RECT 284.985 67.905 285.305 67.965 ;
        RECT 289.140 67.905 289.430 67.950 ;
        RECT 263.915 67.765 278.315 67.905 ;
        RECT 230.260 67.040 230.550 67.270 ;
        RECT 236.225 67.025 236.545 67.285 ;
        RECT 236.685 67.225 237.005 67.285 ;
        RECT 237.160 67.225 237.450 67.270 ;
        RECT 236.685 67.085 237.450 67.225 ;
        RECT 236.685 67.025 237.005 67.085 ;
        RECT 237.160 67.040 237.450 67.085 ;
        RECT 237.620 67.040 237.910 67.270 ;
        RECT 238.065 67.225 238.385 67.285 ;
        RECT 240.365 67.225 240.685 67.285 ;
        RECT 238.065 67.085 240.685 67.225 ;
        RECT 228.495 66.885 228.635 67.025 ;
        RECT 233.465 66.885 233.785 66.945 ;
        RECT 237.695 66.885 237.835 67.040 ;
        RECT 238.065 67.025 238.385 67.085 ;
        RECT 240.365 67.025 240.685 67.085 ;
        RECT 248.645 67.025 248.965 67.285 ;
        RECT 250.485 67.225 250.805 67.285 ;
        RECT 254.640 67.225 254.930 67.270 ;
        RECT 250.485 67.085 254.930 67.225 ;
        RECT 250.485 67.025 250.805 67.085 ;
        RECT 254.640 67.040 254.930 67.085 ;
        RECT 256.480 67.225 256.770 67.270 ;
        RECT 257.385 67.225 257.705 67.285 ;
        RECT 256.480 67.085 257.705 67.225 ;
        RECT 256.480 67.040 256.770 67.085 ;
        RECT 257.385 67.025 257.705 67.085 ;
        RECT 259.010 67.040 259.300 67.270 ;
        RECT 226.655 66.745 228.635 66.885 ;
        RECT 230.335 66.745 237.835 66.885 ;
        RECT 252.325 66.885 252.645 66.945 ;
        RECT 259.085 66.885 259.225 67.040 ;
        RECT 260.145 67.025 260.465 67.285 ;
        RECT 260.695 67.270 260.835 67.705 ;
        RECT 263.915 67.610 264.055 67.765 ;
        RECT 278.175 67.625 278.315 67.765 ;
        RECT 284.985 67.765 289.430 67.905 ;
        RECT 284.985 67.705 285.305 67.765 ;
        RECT 289.140 67.720 289.430 67.765 ;
        RECT 303.845 67.905 304.165 67.965 ;
        RECT 303.845 67.765 306.835 67.905 ;
        RECT 303.845 67.705 304.165 67.765 ;
        RECT 263.380 67.565 263.670 67.610 ;
        RECT 262.075 67.425 263.670 67.565 ;
        RECT 260.695 67.085 261.090 67.270 ;
        RECT 260.800 67.040 261.090 67.085 ;
        RECT 261.540 67.040 261.830 67.270 ;
        RECT 252.325 66.745 259.225 66.885 ;
        RECT 259.685 66.885 260.005 66.945 ;
        RECT 261.615 66.885 261.755 67.040 ;
        RECT 259.685 66.745 261.755 66.885 ;
        RECT 223.360 66.700 223.650 66.745 ;
        RECT 223.895 66.605 224.035 66.745 ;
        RECT 186.175 66.405 189.075 66.545 ;
        RECT 189.270 66.545 189.560 66.590 ;
        RECT 191.160 66.545 191.450 66.590 ;
        RECT 194.280 66.545 194.570 66.590 ;
        RECT 189.270 66.405 194.570 66.545 ;
        RECT 169.065 66.005 169.385 66.265 ;
        RECT 186.175 66.250 186.315 66.405 ;
        RECT 189.270 66.360 189.560 66.405 ;
        RECT 191.160 66.360 191.450 66.405 ;
        RECT 194.280 66.360 194.570 66.405 ;
        RECT 196.665 66.545 196.985 66.605 ;
        RECT 219.205 66.545 219.525 66.605 ;
        RECT 196.665 66.405 219.525 66.545 ;
        RECT 196.665 66.345 196.985 66.405 ;
        RECT 219.205 66.345 219.525 66.405 ;
        RECT 223.805 66.345 224.125 66.605 ;
        RECT 228.405 66.345 228.725 66.605 ;
        RECT 230.335 66.545 230.475 66.745 ;
        RECT 233.465 66.685 233.785 66.745 ;
        RECT 252.325 66.685 252.645 66.745 ;
        RECT 259.685 66.685 260.005 66.745 ;
        RECT 229.875 66.405 230.475 66.545 ;
        RECT 186.100 66.020 186.390 66.250 ;
        RECT 187.465 66.005 187.785 66.265 ;
        RECT 197.585 66.205 197.905 66.265 ;
        RECT 229.875 66.205 230.015 66.405 ;
        RECT 242.205 66.345 242.525 66.605 ;
        RECT 242.665 66.545 242.985 66.605 ;
        RECT 256.005 66.545 256.325 66.605 ;
        RECT 262.075 66.545 262.215 67.425 ;
        RECT 263.380 67.380 263.670 67.425 ;
        RECT 263.840 67.380 264.130 67.610 ;
        RECT 268.425 67.565 268.745 67.625 ;
        RECT 271.185 67.565 271.505 67.625 ;
        RECT 264.375 67.425 268.745 67.565 ;
        RECT 264.375 67.285 264.515 67.425 ;
        RECT 268.425 67.365 268.745 67.425 ;
        RECT 269.665 67.425 271.505 67.565 ;
        RECT 262.920 67.225 263.210 67.270 ;
        RECT 264.285 67.225 264.605 67.285 ;
        RECT 262.920 67.085 264.605 67.225 ;
        RECT 262.920 67.040 263.210 67.085 ;
        RECT 264.285 67.025 264.605 67.085 ;
        RECT 264.760 67.225 265.050 67.270 ;
        RECT 267.045 67.225 267.365 67.285 ;
        RECT 264.760 67.085 267.365 67.225 ;
        RECT 264.760 67.040 265.050 67.085 ;
        RECT 267.045 67.025 267.365 67.085 ;
        RECT 268.900 67.225 269.190 67.270 ;
        RECT 269.665 67.225 269.805 67.425 ;
        RECT 271.185 67.365 271.505 67.425 ;
        RECT 273.025 67.565 273.345 67.625 ;
        RECT 273.940 67.565 274.590 67.610 ;
        RECT 277.540 67.565 277.830 67.610 ;
        RECT 273.025 67.425 277.830 67.565 ;
        RECT 273.025 67.365 273.345 67.425 ;
        RECT 273.940 67.380 274.590 67.425 ;
        RECT 277.240 67.380 277.830 67.425 ;
        RECT 268.900 67.085 269.805 67.225 ;
        RECT 268.900 67.040 269.190 67.085 ;
        RECT 270.265 67.025 270.585 67.285 ;
        RECT 270.745 67.225 271.035 67.270 ;
        RECT 272.580 67.225 272.870 67.270 ;
        RECT 276.160 67.225 276.450 67.270 ;
        RECT 270.745 67.085 276.450 67.225 ;
        RECT 270.745 67.040 271.035 67.085 ;
        RECT 272.580 67.040 272.870 67.085 ;
        RECT 276.160 67.040 276.450 67.085 ;
        RECT 276.705 67.025 277.025 67.285 ;
        RECT 277.240 67.065 277.530 67.380 ;
        RECT 278.085 67.365 278.405 67.625 ;
        RECT 281.305 67.565 281.625 67.625 ;
        RECT 281.780 67.565 282.070 67.610 ;
        RECT 281.305 67.425 282.070 67.565 ;
        RECT 281.305 67.365 281.625 67.425 ;
        RECT 281.780 67.380 282.070 67.425 ;
        RECT 284.060 67.565 284.710 67.610 ;
        RECT 287.660 67.565 287.950 67.610 ;
        RECT 290.965 67.565 291.285 67.625 ;
        RECT 284.060 67.425 291.285 67.565 ;
        RECT 284.060 67.380 284.710 67.425 ;
        RECT 287.360 67.380 287.950 67.425 ;
        RECT 280.865 67.225 281.155 67.270 ;
        RECT 282.700 67.225 282.990 67.270 ;
        RECT 286.280 67.225 286.570 67.270 ;
        RECT 280.865 67.085 286.570 67.225 ;
        RECT 280.865 67.040 281.155 67.085 ;
        RECT 282.700 67.040 282.990 67.085 ;
        RECT 286.280 67.040 286.570 67.085 ;
        RECT 287.360 67.065 287.650 67.380 ;
        RECT 290.965 67.365 291.285 67.425 ;
        RECT 298.780 67.565 299.430 67.610 ;
        RECT 302.380 67.565 302.670 67.610 ;
        RECT 303.385 67.565 303.705 67.625 ;
        RECT 306.695 67.610 306.835 67.765 ;
        RECT 304.780 67.565 305.070 67.610 ;
        RECT 298.780 67.425 305.070 67.565 ;
        RECT 298.780 67.380 299.430 67.425 ;
        RECT 302.080 67.380 302.670 67.425 ;
        RECT 293.725 67.025 294.045 67.285 ;
        RECT 294.185 67.225 294.505 67.285 ;
        RECT 295.120 67.225 295.410 67.270 ;
        RECT 294.185 67.085 295.410 67.225 ;
        RECT 294.185 67.025 294.505 67.085 ;
        RECT 295.120 67.040 295.410 67.085 ;
        RECT 295.585 67.225 295.875 67.270 ;
        RECT 297.420 67.225 297.710 67.270 ;
        RECT 301.000 67.225 301.290 67.270 ;
        RECT 295.585 67.085 301.290 67.225 ;
        RECT 295.585 67.040 295.875 67.085 ;
        RECT 297.420 67.040 297.710 67.085 ;
        RECT 301.000 67.040 301.290 67.085 ;
        RECT 302.080 67.065 302.370 67.380 ;
        RECT 303.385 67.365 303.705 67.425 ;
        RECT 304.780 67.380 305.070 67.425 ;
        RECT 306.620 67.380 306.910 67.610 ;
        RECT 271.660 66.885 271.950 66.930 ;
        RECT 269.895 66.745 271.950 66.885 ;
        RECT 265.205 66.545 265.525 66.605 ;
        RECT 269.895 66.590 270.035 66.745 ;
        RECT 271.660 66.700 271.950 66.745 ;
        RECT 274.865 66.885 275.185 66.945 ;
        RECT 276.795 66.885 276.935 67.025 ;
        RECT 274.865 66.745 276.935 66.885 ;
        RECT 274.865 66.685 275.185 66.745 ;
        RECT 242.665 66.405 256.325 66.545 ;
        RECT 242.665 66.345 242.985 66.405 ;
        RECT 256.005 66.345 256.325 66.405 ;
        RECT 257.015 66.405 258.995 66.545 ;
        RECT 197.585 66.065 230.015 66.205 ;
        RECT 197.585 66.005 197.905 66.065 ;
        RECT 230.245 66.005 230.565 66.265 ;
        RECT 238.985 66.005 239.305 66.265 ;
        RECT 249.565 66.205 249.885 66.265 ;
        RECT 257.015 66.205 257.155 66.405 ;
        RECT 249.565 66.065 257.155 66.205 ;
        RECT 249.565 66.005 249.885 66.065 ;
        RECT 257.385 66.005 257.705 66.265 ;
        RECT 258.305 66.005 258.625 66.265 ;
        RECT 258.855 66.205 258.995 66.405 ;
        RECT 261.615 66.405 265.525 66.545 ;
        RECT 261.615 66.205 261.755 66.405 ;
        RECT 265.205 66.345 265.525 66.405 ;
        RECT 269.820 66.360 270.110 66.590 ;
        RECT 271.150 66.545 271.440 66.590 ;
        RECT 273.040 66.545 273.330 66.590 ;
        RECT 276.160 66.545 276.450 66.590 ;
        RECT 271.150 66.405 276.450 66.545 ;
        RECT 276.795 66.545 276.935 66.745 ;
        RECT 277.625 66.885 277.945 66.945 ;
        RECT 280.385 66.885 280.705 66.945 ;
        RECT 296.500 66.885 296.790 66.930 ;
        RECT 277.625 66.745 280.705 66.885 ;
        RECT 277.625 66.685 277.945 66.745 ;
        RECT 280.385 66.685 280.705 66.745 ;
        RECT 294.735 66.745 296.790 66.885 ;
        RECT 294.735 66.590 294.875 66.745 ;
        RECT 296.500 66.700 296.790 66.745 ;
        RECT 279.020 66.545 279.310 66.590 ;
        RECT 276.795 66.405 279.310 66.545 ;
        RECT 271.150 66.360 271.440 66.405 ;
        RECT 273.040 66.360 273.330 66.405 ;
        RECT 276.160 66.360 276.450 66.405 ;
        RECT 279.020 66.360 279.310 66.405 ;
        RECT 281.270 66.545 281.560 66.590 ;
        RECT 283.160 66.545 283.450 66.590 ;
        RECT 286.280 66.545 286.570 66.590 ;
        RECT 281.270 66.405 286.570 66.545 ;
        RECT 281.270 66.360 281.560 66.405 ;
        RECT 283.160 66.360 283.450 66.405 ;
        RECT 286.280 66.360 286.570 66.405 ;
        RECT 294.660 66.360 294.950 66.590 ;
        RECT 295.990 66.545 296.280 66.590 ;
        RECT 297.880 66.545 298.170 66.590 ;
        RECT 301.000 66.545 301.290 66.590 ;
        RECT 295.990 66.405 301.290 66.545 ;
        RECT 295.990 66.360 296.280 66.405 ;
        RECT 297.880 66.360 298.170 66.405 ;
        RECT 301.000 66.360 301.290 66.405 ;
        RECT 258.855 66.065 261.755 66.205 ;
        RECT 261.985 66.005 262.305 66.265 ;
        RECT 263.365 66.205 263.685 66.265 ;
        RECT 279.465 66.205 279.785 66.265 ;
        RECT 263.365 66.065 279.785 66.205 ;
        RECT 263.365 66.005 263.685 66.065 ;
        RECT 279.465 66.005 279.785 66.065 ;
        RECT 303.845 66.005 304.165 66.265 ;
        RECT 162.095 65.385 311.135 65.865 ;
        RECT 169.985 65.185 170.305 65.245 ;
        RECT 175.520 65.185 175.810 65.230 ;
        RECT 169.985 65.045 175.810 65.185 ;
        RECT 169.985 64.985 170.305 65.045 ;
        RECT 175.520 65.000 175.810 65.045 ;
        RECT 177.345 64.985 177.665 65.245 ;
        RECT 197.585 65.185 197.905 65.245 ;
        RECT 185.715 65.045 197.905 65.185 ;
        RECT 166.270 64.845 166.560 64.890 ;
        RECT 168.160 64.845 168.450 64.890 ;
        RECT 171.280 64.845 171.570 64.890 ;
        RECT 166.270 64.705 171.570 64.845 ;
        RECT 166.270 64.660 166.560 64.705 ;
        RECT 168.160 64.660 168.450 64.705 ;
        RECT 171.280 64.660 171.570 64.705 ;
        RECT 177.435 64.845 177.575 64.985 ;
        RECT 181.945 64.845 182.265 64.905 ;
        RECT 177.435 64.705 182.265 64.845 ;
        RECT 166.780 64.505 167.070 64.550 ;
        RECT 169.065 64.505 169.385 64.565 ;
        RECT 166.780 64.365 169.385 64.505 ;
        RECT 166.780 64.320 167.070 64.365 ;
        RECT 169.065 64.305 169.385 64.365 ;
        RECT 174.140 64.320 174.430 64.550 ;
        RECT 177.435 64.505 177.575 64.705 ;
        RECT 181.945 64.645 182.265 64.705 ;
        RECT 177.820 64.505 178.110 64.550 ;
        RECT 177.435 64.365 178.110 64.505 ;
        RECT 177.820 64.320 178.110 64.365 ;
        RECT 165.385 63.965 165.705 64.225 ;
        RECT 165.865 64.165 166.155 64.210 ;
        RECT 167.700 64.165 167.990 64.210 ;
        RECT 171.280 64.165 171.570 64.210 ;
        RECT 165.865 64.025 171.570 64.165 ;
        RECT 165.865 63.980 166.155 64.025 ;
        RECT 167.700 63.980 167.990 64.025 ;
        RECT 171.280 63.980 171.570 64.025 ;
        RECT 172.285 64.185 172.605 64.225 ;
        RECT 172.285 63.965 172.650 64.185 ;
        RECT 174.215 64.165 174.355 64.320 ;
        RECT 178.725 64.305 179.045 64.565 ;
        RECT 177.360 64.165 177.650 64.210 ;
        RECT 185.715 64.165 185.855 65.045 ;
        RECT 197.585 64.985 197.905 65.045 ;
        RECT 205.420 65.000 205.710 65.230 ;
        RECT 206.340 65.185 206.630 65.230 ;
        RECT 207.705 65.185 208.025 65.245 ;
        RECT 206.340 65.045 208.025 65.185 ;
        RECT 206.340 65.000 206.630 65.045 ;
        RECT 186.970 64.845 187.260 64.890 ;
        RECT 188.860 64.845 189.150 64.890 ;
        RECT 191.980 64.845 192.270 64.890 ;
        RECT 186.970 64.705 192.270 64.845 ;
        RECT 186.970 64.660 187.260 64.705 ;
        RECT 188.860 64.660 189.150 64.705 ;
        RECT 191.980 64.660 192.270 64.705 ;
        RECT 192.525 64.645 192.845 64.905 ;
        RECT 194.840 64.845 195.130 64.890 ;
        RECT 196.665 64.845 196.985 64.905 ;
        RECT 194.840 64.705 196.985 64.845 ;
        RECT 194.840 64.660 195.130 64.705 ;
        RECT 196.665 64.645 196.985 64.705 ;
        RECT 186.085 64.305 186.405 64.565 ;
        RECT 187.465 64.305 187.785 64.565 ;
        RECT 192.615 64.505 192.755 64.645 ;
        RECT 200.345 64.505 200.665 64.565 ;
        RECT 192.615 64.365 200.665 64.505 ;
        RECT 205.495 64.505 205.635 65.000 ;
        RECT 207.705 64.985 208.025 65.045 ;
        RECT 208.625 65.185 208.945 65.245 ;
        RECT 213.240 65.185 213.530 65.230 ;
        RECT 208.625 65.045 213.530 65.185 ;
        RECT 208.625 64.985 208.945 65.045 ;
        RECT 213.240 65.000 213.530 65.045 ;
        RECT 214.160 65.185 214.450 65.230 ;
        RECT 214.605 65.185 214.925 65.245 ;
        RECT 221.505 65.185 221.825 65.245 ;
        RECT 214.160 65.045 214.925 65.185 ;
        RECT 214.160 65.000 214.450 65.045 ;
        RECT 214.605 64.985 214.925 65.045 ;
        RECT 215.155 65.045 221.825 65.185 ;
        RECT 206.785 64.845 207.105 64.905 ;
        RECT 211.400 64.845 211.690 64.890 ;
        RECT 206.785 64.705 211.690 64.845 ;
        RECT 206.785 64.645 207.105 64.705 ;
        RECT 211.400 64.660 211.690 64.705 ;
        RECT 211.845 64.845 212.165 64.905 ;
        RECT 215.155 64.845 215.295 65.045 ;
        RECT 221.505 64.985 221.825 65.045 ;
        RECT 222.885 65.185 223.205 65.245 ;
        RECT 224.725 65.185 225.045 65.245 ;
        RECT 231.165 65.185 231.485 65.245 ;
        RECT 222.885 65.045 231.485 65.185 ;
        RECT 222.885 64.985 223.205 65.045 ;
        RECT 224.725 64.985 225.045 65.045 ;
        RECT 231.165 64.985 231.485 65.045 ;
        RECT 238.985 65.185 239.305 65.245 ;
        RECT 250.040 65.185 250.330 65.230 ;
        RECT 257.385 65.185 257.705 65.245 ;
        RECT 258.320 65.185 258.610 65.230 ;
        RECT 238.985 65.045 250.330 65.185 ;
        RECT 238.985 64.985 239.305 65.045 ;
        RECT 250.040 65.000 250.330 65.045 ;
        RECT 250.575 65.045 253.475 65.185 ;
        RECT 211.845 64.705 215.295 64.845 ;
        RECT 216.905 64.845 217.225 64.905 ;
        RECT 230.245 64.845 230.565 64.905 ;
        RECT 239.445 64.845 239.765 64.905 ;
        RECT 216.905 64.705 239.765 64.845 ;
        RECT 211.845 64.645 212.165 64.705 ;
        RECT 216.905 64.645 217.225 64.705 ;
        RECT 230.245 64.645 230.565 64.705 ;
        RECT 239.445 64.645 239.765 64.705 ;
        RECT 243.125 64.645 243.445 64.905 ;
        RECT 250.575 64.845 250.715 65.045 ;
        RECT 243.675 64.705 250.715 64.845 ;
        RECT 208.625 64.505 208.945 64.565 ;
        RECT 205.495 64.365 208.945 64.505 ;
        RECT 200.345 64.305 200.665 64.365 ;
        RECT 208.625 64.305 208.945 64.365 ;
        RECT 210.020 64.505 210.310 64.550 ;
        RECT 221.060 64.505 221.350 64.550 ;
        RECT 223.805 64.505 224.125 64.565 ;
        RECT 225.200 64.505 225.490 64.550 ;
        RECT 243.675 64.505 243.815 64.705 ;
        RECT 252.800 64.660 253.090 64.890 ;
        RECT 253.335 64.845 253.475 65.045 ;
        RECT 257.385 65.045 258.610 65.185 ;
        RECT 257.385 64.985 257.705 65.045 ;
        RECT 258.320 65.000 258.610 65.045 ;
        RECT 258.780 65.185 259.070 65.230 ;
        RECT 259.225 65.185 259.545 65.245 ;
        RECT 258.780 65.045 259.545 65.185 ;
        RECT 258.780 65.000 259.070 65.045 ;
        RECT 259.225 64.985 259.545 65.045 ;
        RECT 263.365 64.985 263.685 65.245 ;
        RECT 293.725 65.185 294.045 65.245 ;
        RECT 294.200 65.185 294.490 65.230 ;
        RECT 293.725 65.045 294.490 65.185 ;
        RECT 293.725 64.985 294.045 65.045 ;
        RECT 294.200 65.000 294.490 65.045 ;
        RECT 263.455 64.845 263.595 64.985 ;
        RECT 253.335 64.705 263.595 64.845 ;
        RECT 267.980 64.845 268.270 64.890 ;
        RECT 271.760 64.845 272.050 64.890 ;
        RECT 274.880 64.845 275.170 64.890 ;
        RECT 276.770 64.845 277.060 64.890 ;
        RECT 267.980 64.705 269.805 64.845 ;
        RECT 267.980 64.660 268.270 64.705 ;
        RECT 252.875 64.505 253.015 64.660 ;
        RECT 210.020 64.365 215.755 64.505 ;
        RECT 210.020 64.320 210.310 64.365 ;
        RECT 174.215 64.025 185.855 64.165 ;
        RECT 186.565 64.165 186.855 64.210 ;
        RECT 188.400 64.165 188.690 64.210 ;
        RECT 191.980 64.165 192.270 64.210 ;
        RECT 186.565 64.025 192.270 64.165 ;
        RECT 177.360 63.980 177.650 64.025 ;
        RECT 186.565 63.980 186.855 64.025 ;
        RECT 188.400 63.980 188.690 64.025 ;
        RECT 191.980 63.980 192.270 64.025 ;
        RECT 193.060 64.165 193.350 64.185 ;
        RECT 196.205 64.165 196.525 64.225 ;
        RECT 193.060 64.025 196.525 64.165 ;
        RECT 172.360 63.870 172.650 63.965 ;
        RECT 193.060 63.870 193.350 64.025 ;
        RECT 196.205 63.965 196.525 64.025 ;
        RECT 203.565 64.165 203.885 64.225 ;
        RECT 208.165 64.165 208.485 64.225 ;
        RECT 203.565 64.025 211.155 64.165 ;
        RECT 203.565 63.965 203.885 64.025 ;
        RECT 208.165 63.965 208.485 64.025 ;
        RECT 169.060 63.825 169.710 63.870 ;
        RECT 172.360 63.825 172.950 63.870 ;
        RECT 169.060 63.685 172.950 63.825 ;
        RECT 169.060 63.640 169.710 63.685 ;
        RECT 172.660 63.640 172.950 63.685 ;
        RECT 189.760 63.825 190.410 63.870 ;
        RECT 193.060 63.825 193.650 63.870 ;
        RECT 206.785 63.825 207.105 63.885 ;
        RECT 207.720 63.825 208.010 63.870 ;
        RECT 189.760 63.685 193.650 63.825 ;
        RECT 189.760 63.640 190.410 63.685 ;
        RECT 193.360 63.640 193.650 63.685 ;
        RECT 205.495 63.685 208.010 63.825 ;
        RECT 197.585 63.485 197.905 63.545 ;
        RECT 204.025 63.485 204.345 63.545 ;
        RECT 205.495 63.530 205.635 63.685 ;
        RECT 206.785 63.625 207.105 63.685 ;
        RECT 207.720 63.640 208.010 63.685 ;
        RECT 208.625 63.825 208.945 63.885 ;
        RECT 210.480 63.825 210.770 63.870 ;
        RECT 208.625 63.685 210.770 63.825 ;
        RECT 211.015 63.825 211.155 64.025 ;
        RECT 213.240 63.825 213.530 63.870 ;
        RECT 211.015 63.685 213.530 63.825 ;
        RECT 208.625 63.625 208.945 63.685 ;
        RECT 210.480 63.640 210.770 63.685 ;
        RECT 213.240 63.640 213.530 63.685 ;
        RECT 205.420 63.485 205.710 63.530 ;
        RECT 197.585 63.345 205.710 63.485 ;
        RECT 215.615 63.485 215.755 64.365 ;
        RECT 221.060 64.365 225.490 64.505 ;
        RECT 221.060 64.320 221.350 64.365 ;
        RECT 223.805 64.305 224.125 64.365 ;
        RECT 225.200 64.320 225.490 64.365 ;
        RECT 238.155 64.365 243.815 64.505 ;
        RECT 250.115 64.365 253.015 64.505 ;
        RECT 220.585 64.165 220.905 64.225 ;
        RECT 221.520 64.165 221.810 64.210 ;
        RECT 223.355 64.165 223.645 64.210 ;
        RECT 220.585 64.025 221.810 64.165 ;
        RECT 223.250 64.025 223.645 64.165 ;
        RECT 220.585 63.965 220.905 64.025 ;
        RECT 221.520 63.980 221.810 64.025 ;
        RECT 223.355 63.980 223.645 64.025 ;
        RECT 224.265 64.165 224.585 64.225 ;
        RECT 224.740 64.165 225.030 64.210 ;
        RECT 224.265 64.025 225.030 64.165 ;
        RECT 219.205 63.825 219.525 63.885 ;
        RECT 223.435 63.825 223.575 63.980 ;
        RECT 224.265 63.965 224.585 64.025 ;
        RECT 224.740 63.980 225.030 64.025 ;
        RECT 225.660 64.165 225.950 64.210 ;
        RECT 230.705 64.165 231.025 64.225 ;
        RECT 225.660 64.025 231.025 64.165 ;
        RECT 225.660 63.980 225.950 64.025 ;
        RECT 230.705 63.965 231.025 64.025 ;
        RECT 238.155 63.825 238.295 64.365 ;
        RECT 239.920 63.980 240.210 64.210 ;
        RECT 219.205 63.685 238.295 63.825 ;
        RECT 219.205 63.625 219.525 63.685 ;
        RECT 222.885 63.485 223.205 63.545 ;
        RECT 215.615 63.345 223.205 63.485 ;
        RECT 197.585 63.285 197.905 63.345 ;
        RECT 204.025 63.285 204.345 63.345 ;
        RECT 205.420 63.300 205.710 63.345 ;
        RECT 222.885 63.285 223.205 63.345 ;
        RECT 223.805 63.285 224.125 63.545 ;
        RECT 232.085 63.485 232.405 63.545 ;
        RECT 239.995 63.485 240.135 63.980 ;
        RECT 240.365 63.965 240.685 64.225 ;
        RECT 241.285 63.965 241.605 64.225 ;
        RECT 242.345 64.165 242.635 64.210 ;
        RECT 249.565 64.165 249.885 64.225 ;
        RECT 250.115 64.210 250.255 64.365 ;
        RECT 253.245 64.305 253.565 64.565 ;
        RECT 259.240 64.505 259.530 64.550 ;
        RECT 261.985 64.505 262.305 64.565 ;
        RECT 268.885 64.505 269.205 64.565 ;
        RECT 254.255 64.365 258.995 64.505 ;
        RECT 242.345 64.025 249.885 64.165 ;
        RECT 242.345 63.980 242.635 64.025 ;
        RECT 249.565 63.965 249.885 64.025 ;
        RECT 250.040 63.980 250.330 64.210 ;
        RECT 250.960 64.165 251.250 64.210 ;
        RECT 253.335 64.165 253.475 64.305 ;
        RECT 254.255 64.210 254.395 64.365 ;
        RECT 250.960 64.025 253.475 64.165 ;
        RECT 250.960 63.980 251.250 64.025 ;
        RECT 253.695 63.980 253.985 64.210 ;
        RECT 254.180 63.980 254.470 64.210 ;
        RECT 240.455 63.825 240.595 63.965 ;
        RECT 241.760 63.825 242.050 63.870 ;
        RECT 240.455 63.685 242.050 63.825 ;
        RECT 241.760 63.640 242.050 63.685 ;
        RECT 252.325 63.625 252.645 63.885 ;
        RECT 253.770 63.825 253.910 63.980 ;
        RECT 254.625 63.965 254.945 64.225 ;
        RECT 255.545 64.165 255.865 64.225 ;
        RECT 255.350 64.025 255.865 64.165 ;
        RECT 255.545 63.965 255.865 64.025 ;
        RECT 256.020 63.980 256.310 64.210 ;
        RECT 257.400 64.165 257.690 64.210 ;
        RECT 258.305 64.165 258.625 64.225 ;
        RECT 257.400 64.025 258.625 64.165 ;
        RECT 258.855 64.165 258.995 64.365 ;
        RECT 259.240 64.365 262.305 64.505 ;
        RECT 259.240 64.320 259.530 64.365 ;
        RECT 261.985 64.305 262.305 64.365 ;
        RECT 263.915 64.365 269.205 64.505 ;
        RECT 269.665 64.505 269.805 64.705 ;
        RECT 271.760 64.705 277.060 64.845 ;
        RECT 271.760 64.660 272.050 64.705 ;
        RECT 274.880 64.660 275.170 64.705 ;
        RECT 276.770 64.660 277.060 64.705 ;
        RECT 284.065 64.845 284.385 64.905 ;
        RECT 284.065 64.705 297.175 64.845 ;
        RECT 284.065 64.645 284.385 64.705 ;
        RECT 276.260 64.505 276.550 64.550 ;
        RECT 269.665 64.365 276.550 64.505 ;
        RECT 263.915 64.165 264.055 64.365 ;
        RECT 268.885 64.305 269.205 64.365 ;
        RECT 276.260 64.320 276.550 64.365 ;
        RECT 277.625 64.305 277.945 64.565 ;
        RECT 290.965 64.305 291.285 64.565 ;
        RECT 291.975 64.550 292.115 64.705 ;
        RECT 291.900 64.320 292.190 64.550 ;
        RECT 296.485 64.305 296.805 64.565 ;
        RECT 297.035 64.550 297.175 64.705 ;
        RECT 296.960 64.505 297.250 64.550 ;
        RECT 306.605 64.505 306.925 64.565 ;
        RECT 296.960 64.365 306.925 64.505 ;
        RECT 296.960 64.320 297.250 64.365 ;
        RECT 306.605 64.305 306.925 64.365 ;
        RECT 258.855 64.025 264.055 64.165 ;
        RECT 267.060 64.165 267.350 64.210 ;
        RECT 269.805 64.165 270.125 64.225 ;
        RECT 267.060 64.025 270.125 64.165 ;
        RECT 257.400 63.980 257.690 64.025 ;
        RECT 253.340 63.685 253.910 63.825 ;
        RECT 256.095 63.825 256.235 63.980 ;
        RECT 258.305 63.965 258.625 64.025 ;
        RECT 267.060 63.980 267.350 64.025 ;
        RECT 269.805 63.965 270.125 64.025 ;
        RECT 259.685 63.825 260.005 63.885 ;
        RECT 270.680 63.870 270.970 64.185 ;
        RECT 271.760 64.165 272.050 64.210 ;
        RECT 275.340 64.165 275.630 64.210 ;
        RECT 277.175 64.165 277.465 64.210 ;
        RECT 271.760 64.025 277.465 64.165 ;
        RECT 271.760 63.980 272.050 64.025 ;
        RECT 275.340 63.980 275.630 64.025 ;
        RECT 277.175 63.980 277.465 64.025 ;
        RECT 283.605 64.165 283.925 64.225 ;
        RECT 284.985 64.165 285.305 64.225 ;
        RECT 283.605 64.025 285.305 64.165 ;
        RECT 283.605 63.965 283.925 64.025 ;
        RECT 284.985 63.965 285.305 64.025 ;
        RECT 285.445 64.165 285.765 64.225 ;
        RECT 292.360 64.165 292.650 64.210 ;
        RECT 303.845 64.165 304.165 64.225 ;
        RECT 285.445 64.025 304.165 64.165 ;
        RECT 285.445 63.965 285.765 64.025 ;
        RECT 292.360 63.980 292.650 64.025 ;
        RECT 303.845 63.965 304.165 64.025 ;
        RECT 256.095 63.685 260.005 63.825 ;
        RECT 232.085 63.345 240.135 63.485 ;
        RECT 232.085 63.285 232.405 63.345 ;
        RECT 251.865 63.285 252.185 63.545 ;
        RECT 252.415 63.485 252.555 63.625 ;
        RECT 253.340 63.485 253.480 63.685 ;
        RECT 259.685 63.625 260.005 63.685 ;
        RECT 270.380 63.825 270.970 63.870 ;
        RECT 272.565 63.825 272.885 63.885 ;
        RECT 273.620 63.825 274.270 63.870 ;
        RECT 270.380 63.685 274.270 63.825 ;
        RECT 270.380 63.640 270.670 63.685 ;
        RECT 272.565 63.625 272.885 63.685 ;
        RECT 273.620 63.640 274.270 63.685 ;
        RECT 284.525 63.825 284.845 63.885 ;
        RECT 286.365 63.825 286.685 63.885 ;
        RECT 284.525 63.685 286.685 63.825 ;
        RECT 284.525 63.625 284.845 63.685 ;
        RECT 286.365 63.625 286.685 63.685 ;
        RECT 252.415 63.345 253.480 63.485 ;
        RECT 256.925 63.485 257.245 63.545 ;
        RECT 257.860 63.485 258.150 63.530 ;
        RECT 256.925 63.345 258.150 63.485 ;
        RECT 256.925 63.285 257.245 63.345 ;
        RECT 257.860 63.300 258.150 63.345 ;
        RECT 258.765 63.485 259.085 63.545 ;
        RECT 264.285 63.485 264.605 63.545 ;
        RECT 258.765 63.345 264.605 63.485 ;
        RECT 258.765 63.285 259.085 63.345 ;
        RECT 264.285 63.285 264.605 63.345 ;
        RECT 265.205 63.485 265.525 63.545 ;
        RECT 283.145 63.485 283.465 63.545 ;
        RECT 265.205 63.345 283.465 63.485 ;
        RECT 265.205 63.285 265.525 63.345 ;
        RECT 283.145 63.285 283.465 63.345 ;
        RECT 284.065 63.485 284.385 63.545 ;
        RECT 288.205 63.485 288.525 63.545 ;
        RECT 284.065 63.345 288.525 63.485 ;
        RECT 284.065 63.285 284.385 63.345 ;
        RECT 288.205 63.285 288.525 63.345 ;
        RECT 297.420 63.485 297.710 63.530 ;
        RECT 298.325 63.485 298.645 63.545 ;
        RECT 297.420 63.345 298.645 63.485 ;
        RECT 297.420 63.300 297.710 63.345 ;
        RECT 298.325 63.285 298.645 63.345 ;
        RECT 299.245 63.285 299.565 63.545 ;
        RECT 162.095 62.665 311.935 63.145 ;
        RECT 172.300 62.280 172.590 62.510 ;
        RECT 174.140 62.465 174.430 62.510 ;
        RECT 175.045 62.465 175.365 62.525 ;
        RECT 174.140 62.325 175.365 62.465 ;
        RECT 174.140 62.280 174.430 62.325 ;
        RECT 164.940 61.600 165.230 61.830 ;
        RECT 169.540 61.785 169.830 61.830 ;
        RECT 172.375 61.785 172.515 62.280 ;
        RECT 175.045 62.265 175.365 62.325 ;
        RECT 178.265 62.265 178.585 62.525 ;
        RECT 184.245 62.465 184.565 62.525 ;
        RECT 205.865 62.465 206.185 62.525 ;
        RECT 184.245 62.325 206.185 62.465 ;
        RECT 184.245 62.265 184.565 62.325 ;
        RECT 205.865 62.265 206.185 62.325 ;
        RECT 206.785 62.465 207.105 62.525 ;
        RECT 208.640 62.465 208.930 62.510 ;
        RECT 206.785 62.325 208.930 62.465 ;
        RECT 206.785 62.265 207.105 62.325 ;
        RECT 208.640 62.280 208.930 62.325 ;
        RECT 209.560 62.465 209.850 62.510 ;
        RECT 215.525 62.465 215.845 62.525 ;
        RECT 218.285 62.465 218.605 62.525 ;
        RECT 209.560 62.325 215.845 62.465 ;
        RECT 209.560 62.280 209.850 62.325 ;
        RECT 203.565 62.125 203.885 62.185 ;
        RECT 207.720 62.125 208.010 62.170 ;
        RECT 203.565 61.985 208.010 62.125 ;
        RECT 208.715 62.125 208.855 62.280 ;
        RECT 215.525 62.265 215.845 62.325 ;
        RECT 216.075 62.325 218.605 62.465 ;
        RECT 210.940 62.125 211.230 62.170 ;
        RECT 216.075 62.125 216.215 62.325 ;
        RECT 218.285 62.265 218.605 62.325 ;
        RECT 218.760 62.465 219.050 62.510 ;
        RECT 219.665 62.465 219.985 62.525 ;
        RECT 218.760 62.325 219.985 62.465 ;
        RECT 218.760 62.280 219.050 62.325 ;
        RECT 219.665 62.265 219.985 62.325 ;
        RECT 223.805 62.465 224.125 62.525 ;
        RECT 271.185 62.465 271.505 62.525 ;
        RECT 272.580 62.465 272.870 62.510 ;
        RECT 223.805 62.325 269.805 62.465 ;
        RECT 223.805 62.265 224.125 62.325 ;
        RECT 233.925 62.125 234.245 62.185 ;
        RECT 257.400 62.125 257.690 62.170 ;
        RECT 262.445 62.125 262.765 62.185 ;
        RECT 208.715 61.985 211.230 62.125 ;
        RECT 203.565 61.925 203.885 61.985 ;
        RECT 207.720 61.940 208.010 61.985 ;
        RECT 210.940 61.940 211.230 61.985 ;
        RECT 211.475 61.985 216.215 62.125 ;
        RECT 226.195 61.985 233.235 62.125 ;
        RECT 193.000 61.785 193.290 61.830 ;
        RECT 198.045 61.785 198.365 61.845 ;
        RECT 169.540 61.645 172.515 61.785 ;
        RECT 173.065 61.645 192.755 61.785 ;
        RECT 169.540 61.600 169.830 61.645 ;
        RECT 165.015 61.445 165.155 61.600 ;
        RECT 173.065 61.445 173.205 61.645 ;
        RECT 165.015 61.305 173.205 61.445 ;
        RECT 174.125 61.445 174.445 61.505 ;
        RECT 174.600 61.445 174.890 61.490 ;
        RECT 174.125 61.305 174.890 61.445 ;
        RECT 174.125 61.245 174.445 61.305 ;
        RECT 174.600 61.260 174.890 61.305 ;
        RECT 175.520 61.260 175.810 61.490 ;
        RECT 175.965 61.445 176.285 61.505 ;
        RECT 178.725 61.445 179.045 61.505 ;
        RECT 175.965 61.305 179.045 61.445 ;
        RECT 175.595 61.105 175.735 61.260 ;
        RECT 175.965 61.245 176.285 61.305 ;
        RECT 178.725 61.245 179.045 61.305 ;
        RECT 179.185 61.245 179.505 61.505 ;
        RECT 192.615 61.445 192.755 61.645 ;
        RECT 193.000 61.645 198.365 61.785 ;
        RECT 193.000 61.600 193.290 61.645 ;
        RECT 198.045 61.585 198.365 61.645 ;
        RECT 202.660 61.785 202.950 61.830 ;
        RECT 202.660 61.645 204.255 61.785 ;
        RECT 202.660 61.600 202.950 61.645 ;
        RECT 197.585 61.445 197.905 61.505 ;
        RECT 203.580 61.445 203.870 61.490 ;
        RECT 192.615 61.305 197.905 61.445 ;
        RECT 197.585 61.245 197.905 61.305 ;
        RECT 202.735 61.305 203.870 61.445 ;
        RECT 204.115 61.445 204.255 61.645 ;
        RECT 204.485 61.585 204.805 61.845 ;
        RECT 205.405 61.445 205.725 61.505 ;
        RECT 211.475 61.445 211.615 61.985 ;
        RECT 212.765 61.785 213.085 61.845 ;
        RECT 214.160 61.785 214.450 61.830 ;
        RECT 212.765 61.645 214.450 61.785 ;
        RECT 212.765 61.585 213.085 61.645 ;
        RECT 214.160 61.600 214.450 61.645 ;
        RECT 215.080 61.785 215.370 61.830 ;
        RECT 217.840 61.785 218.130 61.830 ;
        RECT 220.585 61.785 220.905 61.845 ;
        RECT 215.080 61.775 217.595 61.785 ;
        RECT 217.735 61.775 220.905 61.785 ;
        RECT 215.080 61.645 220.905 61.775 ;
        RECT 215.080 61.600 215.370 61.645 ;
        RECT 215.615 61.505 215.755 61.645 ;
        RECT 217.455 61.635 218.130 61.645 ;
        RECT 217.840 61.600 218.130 61.635 ;
        RECT 220.585 61.585 220.905 61.645 ;
        RECT 204.115 61.305 211.615 61.445 ;
        RECT 179.275 61.105 179.415 61.245 ;
        RECT 202.735 61.165 202.875 61.305 ;
        RECT 203.580 61.260 203.870 61.305 ;
        RECT 205.405 61.245 205.725 61.305 ;
        RECT 215.525 61.245 215.845 61.505 ;
        RECT 215.985 61.245 216.305 61.505 ;
        RECT 216.905 61.245 217.225 61.505 ;
        RECT 219.680 61.445 219.970 61.490 ;
        RECT 220.125 61.445 220.445 61.505 ;
        RECT 219.680 61.305 220.445 61.445 ;
        RECT 219.680 61.260 219.970 61.305 ;
        RECT 220.125 61.245 220.445 61.305 ;
        RECT 175.595 60.965 179.415 61.105 ;
        RECT 202.645 61.105 202.965 61.165 ;
        RECT 204.025 61.105 204.345 61.165 ;
        RECT 202.645 60.965 204.345 61.105 ;
        RECT 202.645 60.905 202.965 60.965 ;
        RECT 204.025 60.905 204.345 60.965 ;
        RECT 205.865 61.105 206.185 61.165 ;
        RECT 214.605 61.105 214.925 61.165 ;
        RECT 216.995 61.105 217.135 61.245 ;
        RECT 226.195 61.105 226.335 61.985 ;
        RECT 229.875 61.830 230.015 61.985 ;
        RECT 228.880 61.600 229.170 61.830 ;
        RECT 229.800 61.600 230.090 61.830 ;
        RECT 231.180 61.785 231.470 61.830 ;
        RECT 230.335 61.645 231.470 61.785 ;
        RECT 205.865 60.965 212.075 61.105 ;
        RECT 205.865 60.905 206.185 60.965 ;
        RECT 164.005 60.565 164.325 60.825 ;
        RECT 168.605 60.565 168.925 60.825 ;
        RECT 175.045 60.765 175.365 60.825 ;
        RECT 176.440 60.765 176.730 60.810 ;
        RECT 175.045 60.625 176.730 60.765 ;
        RECT 175.045 60.565 175.365 60.625 ;
        RECT 176.440 60.580 176.730 60.625 ;
        RECT 192.065 60.565 192.385 60.825 ;
        RECT 192.525 60.765 192.845 60.825 ;
        RECT 203.120 60.765 203.410 60.810 ;
        RECT 192.525 60.625 203.410 60.765 ;
        RECT 192.525 60.565 192.845 60.625 ;
        RECT 203.120 60.580 203.410 60.625 ;
        RECT 208.625 60.565 208.945 60.825 ;
        RECT 210.925 60.765 211.245 60.825 ;
        RECT 211.400 60.765 211.690 60.810 ;
        RECT 210.925 60.625 211.690 60.765 ;
        RECT 211.935 60.765 212.075 60.965 ;
        RECT 214.605 60.965 217.135 61.105 ;
        RECT 217.455 60.965 226.335 61.105 ;
        RECT 226.565 61.105 226.885 61.165 ;
        RECT 228.955 61.105 229.095 61.600 ;
        RECT 229.325 61.445 229.645 61.505 ;
        RECT 230.335 61.445 230.475 61.645 ;
        RECT 231.180 61.600 231.470 61.645 ;
        RECT 231.625 61.785 231.945 61.845 ;
        RECT 232.100 61.785 232.390 61.830 ;
        RECT 231.625 61.645 232.390 61.785 ;
        RECT 231.625 61.585 231.945 61.645 ;
        RECT 232.100 61.600 232.390 61.645 ;
        RECT 232.545 61.585 232.865 61.845 ;
        RECT 233.095 61.830 233.235 61.985 ;
        RECT 233.925 61.985 254.395 62.125 ;
        RECT 233.925 61.925 234.245 61.985 ;
        RECT 233.020 61.600 233.310 61.830 ;
        RECT 235.305 61.785 235.625 61.845 ;
        RECT 236.240 61.785 236.530 61.830 ;
        RECT 235.305 61.645 236.530 61.785 ;
        RECT 235.305 61.585 235.625 61.645 ;
        RECT 236.240 61.600 236.530 61.645 ;
        RECT 236.685 61.785 237.005 61.845 ;
        RECT 250.485 61.785 250.805 61.845 ;
        RECT 253.705 61.785 254.025 61.845 ;
        RECT 236.685 61.645 254.025 61.785 ;
        RECT 236.685 61.585 237.005 61.645 ;
        RECT 250.485 61.585 250.805 61.645 ;
        RECT 253.705 61.585 254.025 61.645 ;
        RECT 229.325 61.305 230.475 61.445 ;
        RECT 230.720 61.445 231.010 61.490 ;
        RECT 235.780 61.445 236.070 61.490 ;
        RECT 230.720 61.305 236.070 61.445 ;
        RECT 229.325 61.245 229.645 61.305 ;
        RECT 230.720 61.260 231.010 61.305 ;
        RECT 235.780 61.260 236.070 61.305 ;
        RECT 237.145 61.445 237.465 61.505 ;
        RECT 241.745 61.445 242.065 61.505 ;
        RECT 237.145 61.305 242.065 61.445 ;
        RECT 237.145 61.245 237.465 61.305 ;
        RECT 241.745 61.245 242.065 61.305 ;
        RECT 250.025 61.445 250.345 61.505 ;
        RECT 252.340 61.445 252.630 61.490 ;
        RECT 250.025 61.305 252.630 61.445 ;
        RECT 254.255 61.445 254.395 61.985 ;
        RECT 257.400 61.985 262.765 62.125 ;
        RECT 269.665 62.125 269.805 62.325 ;
        RECT 271.185 62.325 272.870 62.465 ;
        RECT 271.185 62.265 271.505 62.325 ;
        RECT 272.580 62.280 272.870 62.325 ;
        RECT 274.865 62.265 275.185 62.525 ;
        RECT 275.325 62.265 275.645 62.525 ;
        RECT 284.080 62.465 284.370 62.510 ;
        RECT 284.985 62.465 285.305 62.525 ;
        RECT 288.220 62.465 288.510 62.510 ;
        RECT 284.080 62.325 284.755 62.465 ;
        RECT 284.080 62.280 284.370 62.325 ;
        RECT 275.415 62.125 275.555 62.265 ;
        RECT 283.605 62.125 283.925 62.185 ;
        RECT 269.665 61.985 275.555 62.125 ;
        RECT 278.175 61.985 283.925 62.125 ;
        RECT 284.615 62.125 284.755 62.325 ;
        RECT 284.985 62.325 288.510 62.465 ;
        RECT 284.985 62.265 285.305 62.325 ;
        RECT 288.220 62.280 288.510 62.325 ;
        RECT 293.740 62.465 294.030 62.510 ;
        RECT 296.025 62.465 296.345 62.525 ;
        RECT 302.940 62.465 303.230 62.510 ;
        RECT 293.740 62.325 295.795 62.465 ;
        RECT 293.740 62.280 294.030 62.325 ;
        RECT 289.125 62.125 289.445 62.185 ;
        RECT 295.655 62.170 295.795 62.325 ;
        RECT 296.025 62.325 303.230 62.465 ;
        RECT 296.025 62.265 296.345 62.325 ;
        RECT 302.940 62.280 303.230 62.325 ;
        RECT 284.615 61.985 289.445 62.125 ;
        RECT 257.400 61.940 257.690 61.985 ;
        RECT 262.445 61.925 262.765 61.985 ;
        RECT 254.640 61.785 254.930 61.830 ;
        RECT 256.940 61.785 257.230 61.830 ;
        RECT 254.640 61.645 257.230 61.785 ;
        RECT 254.640 61.600 254.930 61.645 ;
        RECT 256.940 61.600 257.230 61.645 ;
        RECT 258.320 61.785 258.610 61.830 ;
        RECT 261.525 61.785 261.845 61.845 ;
        RECT 274.420 61.785 274.710 61.830 ;
        RECT 278.175 61.785 278.315 61.985 ;
        RECT 283.605 61.925 283.925 61.985 ;
        RECT 289.125 61.925 289.445 61.985 ;
        RECT 295.580 61.940 295.870 62.170 ;
        RECT 297.860 62.125 298.510 62.170 ;
        RECT 301.460 62.125 301.750 62.170 ;
        RECT 297.860 61.985 301.750 62.125 ;
        RECT 297.860 61.940 298.510 61.985 ;
        RECT 301.160 61.940 301.750 61.985 ;
        RECT 258.320 61.645 261.845 61.785 ;
        RECT 258.320 61.600 258.610 61.645 ;
        RECT 261.525 61.585 261.845 61.645 ;
        RECT 269.665 61.645 278.315 61.785 ;
        RECT 269.665 61.445 269.805 61.645 ;
        RECT 274.420 61.600 274.710 61.645 ;
        RECT 278.545 61.585 278.865 61.845 ;
        RECT 279.465 61.785 279.785 61.845 ;
        RECT 279.940 61.785 280.230 61.830 ;
        RECT 279.465 61.645 280.230 61.785 ;
        RECT 279.465 61.585 279.785 61.645 ;
        RECT 279.940 61.600 280.230 61.645 ;
        RECT 283.145 61.785 283.465 61.845 ;
        RECT 287.760 61.785 288.050 61.830 ;
        RECT 288.205 61.785 288.525 61.845 ;
        RECT 283.145 61.585 283.605 61.785 ;
        RECT 287.760 61.645 288.525 61.785 ;
        RECT 287.760 61.600 288.050 61.645 ;
        RECT 288.205 61.585 288.525 61.645 ;
        RECT 292.820 61.785 293.110 61.830 ;
        RECT 293.725 61.785 294.045 61.845 ;
        RECT 292.820 61.645 294.045 61.785 ;
        RECT 292.820 61.600 293.110 61.645 ;
        RECT 293.725 61.585 294.045 61.645 ;
        RECT 294.665 61.785 294.955 61.830 ;
        RECT 296.500 61.785 296.790 61.830 ;
        RECT 300.080 61.785 300.370 61.830 ;
        RECT 294.665 61.645 300.370 61.785 ;
        RECT 294.665 61.600 294.955 61.645 ;
        RECT 296.500 61.600 296.790 61.645 ;
        RECT 300.080 61.600 300.370 61.645 ;
        RECT 301.160 61.785 301.450 61.940 ;
        RECT 305.225 61.785 305.545 61.845 ;
        RECT 301.160 61.645 305.545 61.785 ;
        RECT 301.160 61.625 301.450 61.645 ;
        RECT 305.225 61.585 305.545 61.645 ;
        RECT 254.255 61.305 269.805 61.445 ;
        RECT 250.025 61.245 250.345 61.305 ;
        RECT 252.340 61.260 252.630 61.305 ;
        RECT 270.725 61.245 271.045 61.505 ;
        RECT 275.325 61.245 275.645 61.505 ;
        RECT 283.465 61.445 283.605 61.585 ;
        RECT 284.065 61.445 284.385 61.505 ;
        RECT 283.465 61.305 284.385 61.445 ;
        RECT 284.065 61.245 284.385 61.305 ;
        RECT 284.525 61.245 284.845 61.505 ;
        RECT 285.460 61.445 285.750 61.490 ;
        RECT 287.300 61.445 287.590 61.490 ;
        RECT 285.075 61.305 290.735 61.445 ;
        RECT 233.465 61.105 233.785 61.165 ;
        RECT 226.565 60.965 233.785 61.105 ;
        RECT 214.605 60.905 214.925 60.965 ;
        RECT 217.455 60.765 217.595 60.965 ;
        RECT 226.565 60.905 226.885 60.965 ;
        RECT 233.465 60.905 233.785 60.965 ;
        RECT 233.925 60.905 234.245 61.165 ;
        RECT 234.400 61.105 234.690 61.150 ;
        RECT 235.305 61.105 235.625 61.165 ;
        RECT 257.845 61.105 258.165 61.165 ;
        RECT 266.585 61.105 266.905 61.165 ;
        RECT 280.860 61.105 281.150 61.150 ;
        RECT 285.075 61.105 285.215 61.305 ;
        RECT 285.460 61.260 285.750 61.305 ;
        RECT 287.300 61.260 287.590 61.305 ;
        RECT 234.400 60.965 235.625 61.105 ;
        RECT 234.400 60.920 234.690 60.965 ;
        RECT 235.305 60.905 235.625 60.965 ;
        RECT 255.865 60.965 266.905 61.105 ;
        RECT 211.935 60.625 217.595 60.765 ;
        RECT 221.505 60.765 221.825 60.825 ;
        RECT 234.015 60.765 234.155 60.905 ;
        RECT 221.505 60.625 234.155 60.765 ;
        RECT 234.860 60.765 235.150 60.810 ;
        RECT 238.065 60.765 238.385 60.825 ;
        RECT 234.860 60.625 238.385 60.765 ;
        RECT 210.925 60.565 211.245 60.625 ;
        RECT 211.400 60.580 211.690 60.625 ;
        RECT 221.505 60.565 221.825 60.625 ;
        RECT 234.860 60.580 235.150 60.625 ;
        RECT 238.065 60.565 238.385 60.625 ;
        RECT 240.365 60.765 240.685 60.825 ;
        RECT 252.800 60.765 253.090 60.810 ;
        RECT 255.865 60.765 256.005 60.965 ;
        RECT 257.845 60.905 258.165 60.965 ;
        RECT 266.585 60.905 266.905 60.965 ;
        RECT 269.665 60.965 279.235 61.105 ;
        RECT 240.365 60.625 256.005 60.765 ;
        RECT 258.320 60.765 258.610 60.810 ;
        RECT 260.605 60.765 260.925 60.825 ;
        RECT 258.320 60.625 260.925 60.765 ;
        RECT 240.365 60.565 240.685 60.625 ;
        RECT 252.800 60.580 253.090 60.625 ;
        RECT 258.320 60.580 258.610 60.625 ;
        RECT 260.605 60.565 260.925 60.625 ;
        RECT 264.285 60.765 264.605 60.825 ;
        RECT 267.520 60.765 267.810 60.810 ;
        RECT 264.285 60.625 267.810 60.765 ;
        RECT 264.285 60.565 264.605 60.625 ;
        RECT 267.520 60.580 267.810 60.625 ;
        RECT 268.425 60.765 268.745 60.825 ;
        RECT 269.665 60.765 269.805 60.965 ;
        RECT 279.095 60.810 279.235 60.965 ;
        RECT 280.860 60.965 285.215 61.105 ;
        RECT 280.860 60.920 281.150 60.965 ;
        RECT 268.425 60.625 269.805 60.765 ;
        RECT 268.425 60.565 268.745 60.625 ;
        RECT 279.020 60.580 279.310 60.810 ;
        RECT 282.225 60.565 282.545 60.825 ;
        RECT 290.045 60.565 290.365 60.825 ;
        RECT 290.595 60.765 290.735 61.305 ;
        RECT 294.185 61.245 294.505 61.505 ;
        RECT 295.070 61.105 295.360 61.150 ;
        RECT 296.960 61.105 297.250 61.150 ;
        RECT 300.080 61.105 300.370 61.150 ;
        RECT 295.070 60.965 300.370 61.105 ;
        RECT 295.070 60.920 295.360 60.965 ;
        RECT 296.960 60.920 297.250 60.965 ;
        RECT 300.080 60.920 300.370 60.965 ;
        RECT 296.485 60.765 296.805 60.825 ;
        RECT 290.595 60.625 296.805 60.765 ;
        RECT 296.485 60.565 296.805 60.625 ;
        RECT 162.095 59.945 311.135 60.425 ;
        RECT 192.525 59.745 192.845 59.805 ;
        RECT 187.095 59.605 192.845 59.745 ;
        RECT 166.270 59.405 166.560 59.450 ;
        RECT 168.160 59.405 168.450 59.450 ;
        RECT 171.280 59.405 171.570 59.450 ;
        RECT 166.270 59.265 171.570 59.405 ;
        RECT 166.270 59.220 166.560 59.265 ;
        RECT 168.160 59.220 168.450 59.265 ;
        RECT 171.280 59.220 171.570 59.265 ;
        RECT 166.780 59.065 167.070 59.110 ;
        RECT 168.605 59.065 168.925 59.125 ;
        RECT 166.780 58.925 168.925 59.065 ;
        RECT 166.780 58.880 167.070 58.925 ;
        RECT 168.605 58.865 168.925 58.925 ;
        RECT 174.585 59.065 174.905 59.125 ;
        RECT 176.425 59.065 176.745 59.125 ;
        RECT 178.280 59.065 178.570 59.110 ;
        RECT 174.585 58.925 178.570 59.065 ;
        RECT 174.585 58.865 174.905 58.925 ;
        RECT 176.425 58.865 176.745 58.925 ;
        RECT 165.385 58.525 165.705 58.785 ;
        RECT 165.865 58.725 166.155 58.770 ;
        RECT 167.700 58.725 167.990 58.770 ;
        RECT 171.280 58.725 171.570 58.770 ;
        RECT 165.865 58.585 171.570 58.725 ;
        RECT 165.865 58.540 166.155 58.585 ;
        RECT 167.700 58.540 167.990 58.585 ;
        RECT 171.280 58.540 171.570 58.585 ;
        RECT 172.360 58.430 172.650 58.745 ;
        RECT 169.060 58.385 169.710 58.430 ;
        RECT 172.360 58.385 172.950 58.430 ;
        RECT 169.060 58.245 174.815 58.385 ;
        RECT 169.060 58.200 169.710 58.245 ;
        RECT 172.660 58.200 172.950 58.245 ;
        RECT 174.675 58.105 174.815 58.245 ;
        RECT 174.125 57.845 174.445 58.105 ;
        RECT 174.585 57.845 174.905 58.105 ;
        RECT 175.965 57.845 176.285 58.105 ;
        RECT 176.975 58.045 177.115 58.925 ;
        RECT 178.280 58.880 178.570 58.925 ;
        RECT 179.185 59.065 179.505 59.125 ;
        RECT 183.340 59.065 183.630 59.110 ;
        RECT 187.095 59.065 187.235 59.605 ;
        RECT 192.525 59.545 192.845 59.605 ;
        RECT 198.045 59.545 198.365 59.805 ;
        RECT 214.605 59.745 214.925 59.805 ;
        RECT 206.875 59.605 214.925 59.745 ;
        RECT 188.810 59.405 189.100 59.450 ;
        RECT 190.700 59.405 190.990 59.450 ;
        RECT 193.820 59.405 194.110 59.450 ;
        RECT 188.810 59.265 194.110 59.405 ;
        RECT 198.135 59.405 198.275 59.545 ;
        RECT 203.120 59.405 203.410 59.450 ;
        RECT 206.875 59.405 207.015 59.605 ;
        RECT 214.605 59.545 214.925 59.605 ;
        RECT 231.625 59.745 231.945 59.805 ;
        RECT 251.405 59.745 251.725 59.805 ;
        RECT 231.625 59.605 251.725 59.745 ;
        RECT 231.625 59.545 231.945 59.605 ;
        RECT 251.405 59.545 251.725 59.605 ;
        RECT 253.705 59.545 254.025 59.805 ;
        RECT 282.225 59.745 282.545 59.805 ;
        RECT 279.095 59.605 282.545 59.745 ;
        RECT 198.135 59.265 203.410 59.405 ;
        RECT 188.810 59.220 189.100 59.265 ;
        RECT 190.700 59.220 190.990 59.265 ;
        RECT 193.820 59.220 194.110 59.265 ;
        RECT 203.120 59.220 203.410 59.265 ;
        RECT 205.495 59.265 207.015 59.405 ;
        RECT 207.245 59.405 207.565 59.465 ;
        RECT 209.100 59.405 209.390 59.450 ;
        RECT 213.685 59.405 214.005 59.465 ;
        RECT 207.245 59.265 214.005 59.405 ;
        RECT 179.185 58.925 187.235 59.065 ;
        RECT 189.320 59.065 189.610 59.110 ;
        RECT 192.065 59.065 192.385 59.125 ;
        RECT 198.060 59.065 198.350 59.110 ;
        RECT 203.565 59.065 203.885 59.125 ;
        RECT 189.320 58.925 192.385 59.065 ;
        RECT 179.185 58.865 179.505 58.925 ;
        RECT 183.340 58.880 183.630 58.925 ;
        RECT 189.320 58.880 189.610 58.925 ;
        RECT 192.065 58.865 192.385 58.925 ;
        RECT 194.455 58.925 197.815 59.065 ;
        RECT 194.455 58.785 194.595 58.925 ;
        RECT 177.345 58.725 177.665 58.785 ;
        RECT 187.925 58.725 188.245 58.785 ;
        RECT 177.345 58.585 188.245 58.725 ;
        RECT 177.345 58.525 177.665 58.585 ;
        RECT 187.925 58.525 188.245 58.585 ;
        RECT 188.405 58.725 188.695 58.770 ;
        RECT 190.240 58.725 190.530 58.770 ;
        RECT 193.820 58.725 194.110 58.770 ;
        RECT 188.405 58.585 194.110 58.725 ;
        RECT 188.405 58.540 188.695 58.585 ;
        RECT 190.240 58.540 190.530 58.585 ;
        RECT 193.820 58.540 194.110 58.585 ;
        RECT 194.365 58.525 194.685 58.785 ;
        RECT 177.805 58.185 178.125 58.445 ;
        RECT 194.900 58.430 195.190 58.745 ;
        RECT 197.675 58.725 197.815 58.925 ;
        RECT 198.060 58.925 203.885 59.065 ;
        RECT 198.060 58.880 198.350 58.925 ;
        RECT 203.565 58.865 203.885 58.925 ;
        RECT 199.440 58.725 199.730 58.770 ;
        RECT 202.645 58.725 202.965 58.785 ;
        RECT 197.675 58.585 199.195 58.725 ;
        RECT 191.600 58.385 192.250 58.430 ;
        RECT 194.900 58.385 195.490 58.430 ;
        RECT 198.045 58.385 198.365 58.445 ;
        RECT 179.735 58.245 191.375 58.385 ;
        RECT 179.735 58.045 179.875 58.245 ;
        RECT 176.975 57.905 179.875 58.045 ;
        RECT 180.120 58.045 180.410 58.090 ;
        RECT 181.485 58.045 181.805 58.105 ;
        RECT 180.120 57.905 181.805 58.045 ;
        RECT 180.120 57.860 180.410 57.905 ;
        RECT 181.485 57.845 181.805 57.905 ;
        RECT 181.945 57.845 182.265 58.105 ;
        RECT 182.420 58.045 182.710 58.090 ;
        RECT 186.085 58.045 186.405 58.105 ;
        RECT 182.420 57.905 186.405 58.045 ;
        RECT 191.235 58.045 191.375 58.245 ;
        RECT 191.600 58.245 198.365 58.385 ;
        RECT 199.055 58.385 199.195 58.585 ;
        RECT 199.440 58.585 202.965 58.725 ;
        RECT 199.440 58.540 199.730 58.585 ;
        RECT 202.645 58.525 202.965 58.585 ;
        RECT 204.945 58.525 205.265 58.785 ;
        RECT 205.495 58.770 205.635 59.265 ;
        RECT 207.245 59.205 207.565 59.265 ;
        RECT 209.100 59.220 209.390 59.265 ;
        RECT 213.685 59.205 214.005 59.265 ;
        RECT 215.065 59.405 215.385 59.465 ;
        RECT 217.840 59.405 218.130 59.450 ;
        RECT 215.065 59.265 218.130 59.405 ;
        RECT 215.065 59.205 215.385 59.265 ;
        RECT 217.840 59.220 218.130 59.265 ;
        RECT 224.280 59.405 224.570 59.450 ;
        RECT 250.485 59.405 250.805 59.465 ;
        RECT 252.785 59.405 253.105 59.465 ;
        RECT 224.280 59.265 235.995 59.405 ;
        RECT 224.280 59.220 224.570 59.265 ;
        RECT 206.340 59.065 206.630 59.110 ;
        RECT 206.785 59.065 207.105 59.125 ;
        RECT 230.245 59.065 230.565 59.125 ;
        RECT 231.625 59.065 231.945 59.125 ;
        RECT 206.340 58.925 207.105 59.065 ;
        RECT 206.340 58.880 206.630 58.925 ;
        RECT 206.785 58.865 207.105 58.925 ;
        RECT 207.340 58.925 229.095 59.065 ;
        RECT 205.420 58.540 205.710 58.770 ;
        RECT 207.340 58.385 207.480 58.925 ;
        RECT 225.275 58.770 225.415 58.925 ;
        RECT 218.760 58.725 219.050 58.770 ;
        RECT 215.615 58.585 219.050 58.725 ;
        RECT 215.615 58.445 215.755 58.585 ;
        RECT 218.760 58.540 219.050 58.585 ;
        RECT 219.680 58.540 219.970 58.770 ;
        RECT 225.200 58.540 225.490 58.770 ;
        RECT 199.055 58.245 207.480 58.385 ;
        RECT 207.720 58.385 208.010 58.430 ;
        RECT 208.625 58.385 208.945 58.445 ;
        RECT 207.720 58.245 208.945 58.385 ;
        RECT 191.600 58.200 192.250 58.245 ;
        RECT 195.200 58.200 195.490 58.245 ;
        RECT 198.045 58.185 198.365 58.245 ;
        RECT 207.720 58.200 208.010 58.245 ;
        RECT 208.625 58.185 208.945 58.245 ;
        RECT 215.525 58.185 215.845 58.445 ;
        RECT 216.445 58.385 216.765 58.445 ;
        RECT 219.755 58.385 219.895 58.540 ;
        RECT 226.105 58.525 226.425 58.785 ;
        RECT 227.040 58.725 227.330 58.770 ;
        RECT 227.485 58.725 227.805 58.785 ;
        RECT 228.955 58.770 229.095 58.925 ;
        RECT 230.245 58.925 231.945 59.065 ;
        RECT 230.245 58.865 230.565 58.925 ;
        RECT 227.040 58.585 227.805 58.725 ;
        RECT 227.040 58.540 227.330 58.585 ;
        RECT 227.485 58.525 227.805 58.585 ;
        RECT 227.960 58.540 228.250 58.770 ;
        RECT 228.420 58.540 228.710 58.770 ;
        RECT 228.880 58.725 229.170 58.770 ;
        RECT 229.325 58.725 229.645 58.785 ;
        RECT 230.795 58.770 230.935 58.925 ;
        RECT 231.625 58.865 231.945 58.925 ;
        RECT 233.465 59.065 233.785 59.125 ;
        RECT 235.855 59.110 235.995 59.265 ;
        RECT 241.835 59.265 243.355 59.405 ;
        RECT 241.835 59.125 241.975 59.265 ;
        RECT 234.860 59.065 235.150 59.110 ;
        RECT 233.465 58.925 235.150 59.065 ;
        RECT 233.465 58.865 233.785 58.925 ;
        RECT 234.860 58.880 235.150 58.925 ;
        RECT 235.780 58.880 236.070 59.110 ;
        RECT 236.240 59.065 236.530 59.110 ;
        RECT 237.605 59.065 237.925 59.125 ;
        RECT 236.240 58.925 237.925 59.065 ;
        RECT 236.240 58.880 236.530 58.925 ;
        RECT 237.605 58.865 237.925 58.925 ;
        RECT 241.745 58.865 242.065 59.125 ;
        RECT 242.680 58.880 242.970 59.110 ;
        RECT 243.215 59.065 243.355 59.265 ;
        RECT 245.055 59.265 253.105 59.405 ;
        RECT 253.795 59.405 253.935 59.545 ;
        RECT 263.380 59.405 263.670 59.450 ;
        RECT 253.795 59.265 256.005 59.405 ;
        RECT 245.055 59.125 245.195 59.265 ;
        RECT 250.485 59.205 250.805 59.265 ;
        RECT 252.785 59.205 253.105 59.265 ;
        RECT 243.600 59.065 243.890 59.110 ;
        RECT 243.215 58.925 243.890 59.065 ;
        RECT 243.600 58.880 243.890 58.925 ;
        RECT 228.880 58.585 229.645 58.725 ;
        RECT 228.880 58.540 229.170 58.585 ;
        RECT 216.445 58.245 219.895 58.385 ;
        RECT 216.445 58.185 216.765 58.245 ;
        RECT 194.365 58.045 194.685 58.105 ;
        RECT 191.235 57.905 194.685 58.045 ;
        RECT 182.420 57.860 182.710 57.905 ;
        RECT 186.085 57.845 186.405 57.905 ;
        RECT 194.365 57.845 194.685 57.905 ;
        RECT 195.745 58.045 196.065 58.105 ;
        RECT 198.520 58.045 198.810 58.090 ;
        RECT 195.745 57.905 198.810 58.045 ;
        RECT 195.745 57.845 196.065 57.905 ;
        RECT 198.520 57.860 198.810 57.905 ;
        RECT 204.945 58.045 205.265 58.105 ;
        RECT 216.535 58.045 216.675 58.185 ;
        RECT 204.945 57.905 216.675 58.045 ;
        RECT 219.755 58.045 219.895 58.245 ;
        RECT 221.505 58.045 221.825 58.105 ;
        RECT 219.755 57.905 221.825 58.045 ;
        RECT 204.945 57.845 205.265 57.905 ;
        RECT 221.505 57.845 221.825 57.905 ;
        RECT 224.725 58.045 225.045 58.105 ;
        RECT 228.035 58.045 228.175 58.540 ;
        RECT 228.495 58.385 228.635 58.540 ;
        RECT 229.325 58.525 229.645 58.585 ;
        RECT 230.720 58.540 231.010 58.770 ;
        RECT 231.165 58.525 231.485 58.785 ;
        RECT 232.085 58.525 232.405 58.785 ;
        RECT 236.685 58.725 237.005 58.785 ;
        RECT 234.935 58.585 237.005 58.725 ;
        RECT 234.935 58.445 235.075 58.585 ;
        RECT 236.685 58.525 237.005 58.585 ;
        RECT 237.160 58.540 237.450 58.770 ;
        RECT 239.000 58.725 239.290 58.770 ;
        RECT 240.365 58.725 240.685 58.785 ;
        RECT 239.000 58.585 240.685 58.725 ;
        RECT 239.000 58.540 239.290 58.585 ;
        RECT 232.545 58.385 232.865 58.445 ;
        RECT 228.495 58.245 232.865 58.385 ;
        RECT 228.955 58.105 229.095 58.245 ;
        RECT 232.545 58.185 232.865 58.245 ;
        RECT 234.385 58.185 234.705 58.445 ;
        RECT 234.845 58.185 235.165 58.445 ;
        RECT 237.235 58.385 237.375 58.540 ;
        RECT 237.605 58.385 237.925 58.445 ;
        RECT 237.235 58.245 237.925 58.385 ;
        RECT 237.605 58.185 237.925 58.245 ;
        RECT 224.725 57.905 228.175 58.045 ;
        RECT 224.725 57.845 225.045 57.905 ;
        RECT 228.865 57.845 229.185 58.105 ;
        RECT 230.245 57.845 230.565 58.105 ;
        RECT 234.475 58.045 234.615 58.185 ;
        RECT 239.075 58.045 239.215 58.540 ;
        RECT 240.365 58.525 240.685 58.585 ;
        RECT 240.840 58.725 241.130 58.770 ;
        RECT 242.220 58.725 242.510 58.770 ;
        RECT 240.840 58.585 242.510 58.725 ;
        RECT 240.840 58.540 241.130 58.585 ;
        RECT 242.220 58.540 242.510 58.585 ;
        RECT 239.920 58.385 240.210 58.430 ;
        RECT 239.920 58.245 241.975 58.385 ;
        RECT 239.920 58.200 240.210 58.245 ;
        RECT 240.915 58.105 241.055 58.245 ;
        RECT 241.835 58.105 241.975 58.245 ;
        RECT 234.475 57.905 239.215 58.045 ;
        RECT 240.825 57.845 241.145 58.105 ;
        RECT 241.285 57.845 241.605 58.105 ;
        RECT 241.745 57.845 242.065 58.105 ;
        RECT 242.755 58.045 242.895 58.880 ;
        RECT 244.965 58.865 245.285 59.125 ;
        RECT 249.105 59.065 249.425 59.125 ;
        RECT 255.865 59.065 256.005 59.265 ;
        RECT 263.380 59.265 265.435 59.405 ;
        RECT 263.380 59.220 263.670 59.265 ;
        RECT 259.700 59.065 259.990 59.110 ;
        RECT 262.460 59.065 262.750 59.110 ;
        RECT 264.300 59.065 264.590 59.110 ;
        RECT 246.895 58.925 249.425 59.065 ;
        RECT 243.140 58.725 243.430 58.770 ;
        RECT 246.895 58.725 247.035 58.925 ;
        RECT 249.105 58.865 249.425 58.925 ;
        RECT 250.575 58.925 255.315 59.065 ;
        RECT 255.865 58.925 259.455 59.065 ;
        RECT 243.140 58.585 247.035 58.725 ;
        RECT 247.265 58.725 247.585 58.785 ;
        RECT 249.580 58.725 249.870 58.770 ;
        RECT 247.265 58.585 249.870 58.725 ;
        RECT 243.140 58.540 243.430 58.585 ;
        RECT 247.265 58.525 247.585 58.585 ;
        RECT 249.580 58.540 249.870 58.585 ;
        RECT 245.440 58.385 245.730 58.430 ;
        RECT 247.725 58.385 248.045 58.445 ;
        RECT 248.200 58.385 248.490 58.430 ;
        RECT 250.025 58.385 250.345 58.445 ;
        RECT 245.440 58.245 250.345 58.385 ;
        RECT 245.440 58.200 245.730 58.245 ;
        RECT 247.725 58.185 248.045 58.245 ;
        RECT 248.200 58.200 248.490 58.245 ;
        RECT 250.025 58.185 250.345 58.245 ;
        RECT 245.885 58.045 246.205 58.105 ;
        RECT 242.755 57.905 246.205 58.045 ;
        RECT 245.885 57.845 246.205 57.905 ;
        RECT 249.105 57.845 249.425 58.105 ;
        RECT 249.565 58.045 249.885 58.105 ;
        RECT 250.575 58.045 250.715 58.925 ;
        RECT 251.865 58.725 252.185 58.785 ;
        RECT 253.245 58.725 253.565 58.785 ;
        RECT 255.175 58.770 255.315 58.925 ;
        RECT 254.180 58.725 254.470 58.770 ;
        RECT 251.865 58.585 254.470 58.725 ;
        RECT 251.865 58.525 252.185 58.585 ;
        RECT 253.245 58.525 253.565 58.585 ;
        RECT 254.180 58.540 254.470 58.585 ;
        RECT 255.100 58.540 255.390 58.770 ;
        RECT 255.545 58.525 255.865 58.785 ;
        RECT 256.020 58.725 256.310 58.770 ;
        RECT 258.780 58.725 259.070 58.770 ;
        RECT 256.020 58.585 259.070 58.725 ;
        RECT 256.020 58.540 256.310 58.585 ;
        RECT 258.780 58.540 259.070 58.585 ;
        RECT 250.945 58.385 251.265 58.445 ;
        RECT 256.095 58.385 256.235 58.540 ;
        RECT 250.945 58.245 256.235 58.385 ;
        RECT 250.945 58.185 251.265 58.245 ;
        RECT 257.845 58.185 258.165 58.445 ;
        RECT 259.315 58.385 259.455 58.925 ;
        RECT 259.700 58.925 262.750 59.065 ;
        RECT 259.700 58.880 259.990 58.925 ;
        RECT 262.460 58.880 262.750 58.925 ;
        RECT 263.455 58.925 264.590 59.065 ;
        RECT 263.455 58.785 263.595 58.925 ;
        RECT 264.300 58.880 264.590 58.925 ;
        RECT 261.065 58.525 261.385 58.785 ;
        RECT 261.540 58.540 261.830 58.770 ;
        RECT 262.000 58.725 262.290 58.770 ;
        RECT 262.905 58.725 263.225 58.785 ;
        RECT 262.000 58.585 263.225 58.725 ;
        RECT 262.000 58.540 262.290 58.585 ;
        RECT 261.615 58.385 261.755 58.540 ;
        RECT 262.905 58.525 263.225 58.585 ;
        RECT 263.365 58.525 263.685 58.785 ;
        RECT 265.295 58.770 265.435 59.265 ;
        RECT 263.840 58.540 264.130 58.770 ;
        RECT 265.220 58.540 265.510 58.770 ;
        RECT 259.315 58.245 261.755 58.385 ;
        RECT 263.915 58.385 264.055 58.540 ;
        RECT 265.665 58.525 265.985 58.785 ;
        RECT 279.095 58.770 279.235 59.605 ;
        RECT 282.225 59.545 282.545 59.605 ;
        RECT 289.125 59.545 289.445 59.805 ;
        RECT 293.725 59.745 294.045 59.805 ;
        RECT 294.660 59.745 294.950 59.790 ;
        RECT 293.725 59.605 294.950 59.745 ;
        RECT 293.725 59.545 294.045 59.605 ;
        RECT 294.660 59.560 294.950 59.605 ;
        RECT 281.270 59.405 281.560 59.450 ;
        RECT 283.160 59.405 283.450 59.450 ;
        RECT 286.280 59.405 286.570 59.450 ;
        RECT 281.270 59.265 286.570 59.405 ;
        RECT 281.270 59.220 281.560 59.265 ;
        RECT 283.160 59.220 283.450 59.265 ;
        RECT 286.280 59.220 286.570 59.265 ;
        RECT 296.485 59.065 296.805 59.125 ;
        RECT 297.420 59.065 297.710 59.110 ;
        RECT 296.485 58.925 297.710 59.065 ;
        RECT 296.485 58.865 296.805 58.925 ;
        RECT 297.420 58.880 297.710 58.925 ;
        RECT 271.660 58.725 271.950 58.770 ;
        RECT 271.660 58.585 272.335 58.725 ;
        RECT 271.660 58.540 271.950 58.585 ;
        RECT 268.440 58.385 268.730 58.430 ;
        RECT 263.915 58.245 268.730 58.385 ;
        RECT 268.440 58.200 268.730 58.245 ;
        RECT 272.195 58.105 272.335 58.585 ;
        RECT 279.020 58.540 279.310 58.770 ;
        RECT 280.385 58.525 280.705 58.785 ;
        RECT 280.865 58.725 281.155 58.770 ;
        RECT 282.700 58.725 282.990 58.770 ;
        RECT 286.280 58.725 286.570 58.770 ;
        RECT 280.865 58.585 286.570 58.725 ;
        RECT 280.865 58.540 281.155 58.585 ;
        RECT 282.700 58.540 282.990 58.585 ;
        RECT 286.280 58.540 286.570 58.585 ;
        RECT 287.360 58.430 287.650 58.745 ;
        RECT 290.045 58.725 290.365 58.785 ;
        RECT 290.520 58.725 290.810 58.770 ;
        RECT 290.045 58.585 290.810 58.725 ;
        RECT 290.045 58.525 290.365 58.585 ;
        RECT 290.520 58.540 290.810 58.585 ;
        RECT 296.025 58.525 296.345 58.785 ;
        RECT 299.245 58.725 299.565 58.785 ;
        RECT 299.720 58.725 300.010 58.770 ;
        RECT 299.245 58.585 300.010 58.725 ;
        RECT 299.245 58.525 299.565 58.585 ;
        RECT 299.720 58.540 300.010 58.585 ;
        RECT 281.780 58.385 282.070 58.430 ;
        RECT 280.015 58.245 282.070 58.385 ;
        RECT 249.565 57.905 250.715 58.045 ;
        RECT 249.565 57.845 249.885 57.905 ;
        RECT 257.385 57.845 257.705 58.105 ;
        RECT 262.445 58.045 262.765 58.105 ;
        RECT 266.125 58.045 266.445 58.105 ;
        RECT 262.445 57.905 266.445 58.045 ;
        RECT 262.445 57.845 262.765 57.905 ;
        RECT 266.125 57.845 266.445 57.905 ;
        RECT 266.585 57.845 266.905 58.105 ;
        RECT 272.105 57.845 272.425 58.105 ;
        RECT 280.015 58.090 280.155 58.245 ;
        RECT 281.780 58.200 282.070 58.245 ;
        RECT 284.060 58.385 284.710 58.430 ;
        RECT 287.360 58.385 287.950 58.430 ;
        RECT 288.665 58.385 288.985 58.445 ;
        RECT 296.115 58.385 296.255 58.525 ;
        RECT 296.500 58.385 296.790 58.430 ;
        RECT 284.060 58.245 295.795 58.385 ;
        RECT 296.115 58.245 296.790 58.385 ;
        RECT 284.060 58.200 284.710 58.245 ;
        RECT 287.660 58.200 287.950 58.245 ;
        RECT 288.665 58.185 288.985 58.245 ;
        RECT 279.940 57.860 280.230 58.090 ;
        RECT 289.585 57.845 289.905 58.105 ;
        RECT 295.655 58.045 295.795 58.245 ;
        RECT 296.500 58.200 296.790 58.245 ;
        RECT 296.960 58.385 297.250 58.430 ;
        RECT 297.405 58.385 297.725 58.445 ;
        RECT 305.225 58.385 305.545 58.445 ;
        RECT 296.960 58.245 297.725 58.385 ;
        RECT 296.960 58.200 297.250 58.245 ;
        RECT 297.405 58.185 297.725 58.245 ;
        RECT 297.955 58.245 305.545 58.385 ;
        RECT 297.955 58.045 298.095 58.245 ;
        RECT 305.225 58.185 305.545 58.245 ;
        RECT 295.655 57.905 298.095 58.045 ;
        RECT 298.785 57.845 299.105 58.105 ;
        RECT 162.095 57.225 311.935 57.705 ;
        RECT 165.385 56.825 165.705 57.085 ;
        RECT 195.745 57.025 196.065 57.085 ;
        RECT 167.775 56.885 177.575 57.025 ;
        RECT 165.475 56.685 165.615 56.825 ;
        RECT 167.775 56.685 167.915 56.885 ;
        RECT 165.475 56.545 167.915 56.685 ;
        RECT 167.775 56.390 167.915 56.545 ;
        RECT 171.360 56.685 172.010 56.730 ;
        RECT 174.960 56.685 175.250 56.730 ;
        RECT 171.360 56.545 175.250 56.685 ;
        RECT 171.360 56.500 172.010 56.545 ;
        RECT 174.660 56.500 175.250 56.545 ;
        RECT 174.660 56.405 174.950 56.500 ;
        RECT 177.435 56.405 177.575 56.885 ;
        RECT 192.615 56.885 196.065 57.025 ;
        RECT 192.615 56.730 192.755 56.885 ;
        RECT 195.745 56.825 196.065 56.885 ;
        RECT 197.585 57.025 197.905 57.085 ;
        RECT 199.900 57.025 200.190 57.070 ;
        RECT 197.585 56.885 200.190 57.025 ;
        RECT 197.585 56.825 197.905 56.885 ;
        RECT 199.900 56.840 200.190 56.885 ;
        RECT 202.645 56.825 202.965 57.085 ;
        RECT 204.500 57.025 204.790 57.070 ;
        RECT 211.385 57.025 211.705 57.085 ;
        RECT 204.500 56.885 211.705 57.025 ;
        RECT 204.500 56.840 204.790 56.885 ;
        RECT 211.385 56.825 211.705 56.885 ;
        RECT 214.145 57.025 214.465 57.085 ;
        RECT 227.500 57.025 227.790 57.070 ;
        RECT 228.405 57.025 228.725 57.085 ;
        RECT 214.145 56.885 227.285 57.025 ;
        RECT 214.145 56.825 214.465 56.885 ;
        RECT 181.020 56.685 181.670 56.730 ;
        RECT 184.620 56.685 184.910 56.730 ;
        RECT 181.020 56.545 184.910 56.685 ;
        RECT 181.020 56.500 181.670 56.545 ;
        RECT 184.320 56.500 184.910 56.545 ;
        RECT 192.540 56.500 192.830 56.730 ;
        RECT 194.820 56.685 195.470 56.730 ;
        RECT 198.420 56.685 198.710 56.730 ;
        RECT 194.820 56.545 198.710 56.685 ;
        RECT 194.820 56.500 195.470 56.545 ;
        RECT 198.120 56.500 198.710 56.545 ;
        RECT 167.240 56.160 167.530 56.390 ;
        RECT 167.700 56.160 167.990 56.390 ;
        RECT 168.165 56.345 168.455 56.390 ;
        RECT 170.000 56.345 170.290 56.390 ;
        RECT 173.580 56.345 173.870 56.390 ;
        RECT 168.165 56.205 173.870 56.345 ;
        RECT 168.165 56.160 168.455 56.205 ;
        RECT 170.000 56.160 170.290 56.205 ;
        RECT 173.580 56.160 173.870 56.205 ;
        RECT 174.585 56.345 174.950 56.405 ;
        RECT 174.585 56.205 177.115 56.345 ;
        RECT 174.585 56.185 174.950 56.205 ;
        RECT 166.320 55.325 166.610 55.370 ;
        RECT 166.765 55.325 167.085 55.385 ;
        RECT 166.320 55.185 167.085 55.325 ;
        RECT 167.315 55.325 167.455 56.160 ;
        RECT 174.585 56.145 174.905 56.185 ;
        RECT 169.065 55.805 169.385 56.065 ;
        RECT 176.425 55.805 176.745 56.065 ;
        RECT 168.570 55.665 168.860 55.710 ;
        RECT 170.460 55.665 170.750 55.710 ;
        RECT 173.580 55.665 173.870 55.710 ;
        RECT 168.570 55.525 173.870 55.665 ;
        RECT 168.570 55.480 168.860 55.525 ;
        RECT 170.460 55.480 170.750 55.525 ;
        RECT 173.580 55.480 173.870 55.525 ;
        RECT 175.045 55.325 175.365 55.385 ;
        RECT 167.315 55.185 175.365 55.325 ;
        RECT 176.975 55.325 177.115 56.205 ;
        RECT 177.345 56.145 177.665 56.405 ;
        RECT 177.825 56.345 178.115 56.390 ;
        RECT 179.660 56.345 179.950 56.390 ;
        RECT 183.240 56.345 183.530 56.390 ;
        RECT 177.825 56.205 183.530 56.345 ;
        RECT 177.825 56.160 178.115 56.205 ;
        RECT 179.660 56.160 179.950 56.205 ;
        RECT 183.240 56.160 183.530 56.205 ;
        RECT 184.320 56.185 184.610 56.500 ;
        RECT 198.120 56.405 198.410 56.500 ;
        RECT 204.945 56.485 205.265 56.745 ;
        RECT 208.640 56.685 208.930 56.730 ;
        RECT 206.415 56.545 208.930 56.685 ;
        RECT 206.415 56.405 206.555 56.545 ;
        RECT 208.640 56.500 208.930 56.545 ;
        RECT 210.925 56.485 211.245 56.745 ;
        RECT 214.605 56.685 214.925 56.745 ;
        RECT 227.145 56.730 227.285 56.885 ;
        RECT 227.500 56.885 228.725 57.025 ;
        RECT 227.500 56.840 227.790 56.885 ;
        RECT 228.405 56.825 228.725 56.885 ;
        RECT 233.925 56.825 234.245 57.085 ;
        RECT 246.820 57.025 247.110 57.070 ;
        RECT 247.265 57.025 247.585 57.085 ;
        RECT 252.340 57.025 252.630 57.070 ;
        RECT 240.455 56.885 245.655 57.025 ;
        RECT 227.070 56.685 227.360 56.730 ;
        RECT 211.935 56.545 215.755 56.685 ;
        RECT 191.625 56.345 191.915 56.390 ;
        RECT 193.460 56.345 193.750 56.390 ;
        RECT 197.040 56.345 197.330 56.390 ;
        RECT 191.625 56.205 197.330 56.345 ;
        RECT 178.725 55.805 179.045 56.065 ;
        RECT 178.230 55.665 178.520 55.710 ;
        RECT 180.120 55.665 180.410 55.710 ;
        RECT 183.240 55.665 183.530 55.710 ;
        RECT 178.230 55.525 183.530 55.665 ;
        RECT 178.230 55.480 178.520 55.525 ;
        RECT 180.120 55.480 180.410 55.525 ;
        RECT 183.240 55.480 183.530 55.525 ;
        RECT 184.335 55.665 184.475 56.185 ;
        RECT 191.625 56.160 191.915 56.205 ;
        RECT 193.460 56.160 193.750 56.205 ;
        RECT 197.040 56.160 197.330 56.205 ;
        RECT 198.045 56.345 198.410 56.405 ;
        RECT 200.345 56.345 200.665 56.405 ;
        RECT 198.045 56.205 200.665 56.345 ;
        RECT 198.045 56.185 198.410 56.205 ;
        RECT 198.045 56.145 198.365 56.185 ;
        RECT 200.345 56.145 200.665 56.205 ;
        RECT 206.325 56.145 206.645 56.405 ;
        RECT 211.935 56.390 212.075 56.545 ;
        RECT 214.605 56.485 214.925 56.545 ;
        RECT 208.180 56.345 208.470 56.390 ;
        RECT 211.860 56.345 212.150 56.390 ;
        RECT 208.180 56.205 212.150 56.345 ;
        RECT 208.180 56.160 208.470 56.205 ;
        RECT 211.860 56.160 212.150 56.205 ;
        RECT 212.305 56.345 212.625 56.405 ;
        RECT 215.615 56.390 215.755 56.545 ;
        RECT 227.070 56.545 230.475 56.685 ;
        RECT 227.070 56.500 227.360 56.545 ;
        RECT 213.240 56.345 213.530 56.390 ;
        RECT 212.305 56.205 213.530 56.345 ;
        RECT 212.305 56.145 212.625 56.205 ;
        RECT 213.240 56.160 213.530 56.205 ;
        RECT 214.160 56.345 214.450 56.390 ;
        RECT 215.540 56.345 215.830 56.390 ;
        RECT 221.045 56.345 221.365 56.405 ;
        RECT 214.160 56.205 215.295 56.345 ;
        RECT 214.160 56.160 214.450 56.205 ;
        RECT 186.545 56.005 186.865 56.065 ;
        RECT 187.480 56.005 187.770 56.050 ;
        RECT 186.545 55.865 187.770 56.005 ;
        RECT 186.545 55.805 186.865 55.865 ;
        RECT 187.480 55.820 187.770 55.865 ;
        RECT 187.925 56.005 188.245 56.065 ;
        RECT 191.160 56.005 191.450 56.050 ;
        RECT 198.135 56.005 198.275 56.145 ;
        RECT 207.705 56.050 208.025 56.065 ;
        RECT 187.925 55.865 191.450 56.005 ;
        RECT 187.925 55.805 188.245 55.865 ;
        RECT 191.160 55.820 191.450 55.865 ;
        RECT 191.695 55.865 198.275 56.005 ;
        RECT 205.880 56.005 206.170 56.050 ;
        RECT 205.880 55.865 207.015 56.005 ;
        RECT 191.695 55.665 191.835 55.865 ;
        RECT 205.880 55.820 206.170 55.865 ;
        RECT 184.335 55.525 191.835 55.665 ;
        RECT 192.030 55.665 192.320 55.710 ;
        RECT 193.920 55.665 194.210 55.710 ;
        RECT 197.040 55.665 197.330 55.710 ;
        RECT 192.030 55.525 197.330 55.665 ;
        RECT 184.335 55.325 184.475 55.525 ;
        RECT 192.030 55.480 192.320 55.525 ;
        RECT 193.920 55.480 194.210 55.525 ;
        RECT 197.040 55.480 197.330 55.525 ;
        RECT 206.875 55.385 207.015 55.865 ;
        RECT 207.595 55.820 208.025 56.050 ;
        RECT 210.020 55.820 210.310 56.050 ;
        RECT 213.315 56.005 213.455 56.160 ;
        RECT 214.620 56.005 214.910 56.050 ;
        RECT 213.315 55.865 214.910 56.005 ;
        RECT 215.155 56.005 215.295 56.205 ;
        RECT 215.540 56.205 221.365 56.345 ;
        RECT 215.540 56.160 215.830 56.205 ;
        RECT 221.045 56.145 221.365 56.205 ;
        RECT 223.805 56.145 224.125 56.405 ;
        RECT 225.645 56.145 225.965 56.405 ;
        RECT 227.960 56.345 228.250 56.390 ;
        RECT 229.800 56.345 230.090 56.390 ;
        RECT 227.575 56.205 230.090 56.345 ;
        RECT 230.335 56.345 230.475 56.545 ;
        RECT 233.940 56.345 234.230 56.390 ;
        RECT 239.445 56.345 239.765 56.405 ;
        RECT 230.335 56.205 239.765 56.345 ;
        RECT 216.460 56.005 216.750 56.050 ;
        RECT 219.205 56.005 219.525 56.065 ;
        RECT 215.155 55.865 215.755 56.005 ;
        RECT 214.620 55.820 214.910 55.865 ;
        RECT 207.705 55.805 208.025 55.820 ;
        RECT 176.975 55.185 184.475 55.325 ;
        RECT 166.320 55.140 166.610 55.185 ;
        RECT 166.765 55.125 167.085 55.185 ;
        RECT 175.045 55.125 175.365 55.185 ;
        RECT 206.785 55.125 207.105 55.385 ;
        RECT 210.095 55.325 210.235 55.820 ;
        RECT 215.615 55.725 215.755 55.865 ;
        RECT 216.460 55.865 219.525 56.005 ;
        RECT 216.460 55.820 216.750 55.865 ;
        RECT 219.205 55.805 219.525 55.865 ;
        RECT 210.465 55.665 210.785 55.725 ;
        RECT 212.780 55.665 213.070 55.710 ;
        RECT 213.225 55.665 213.545 55.725 ;
        RECT 210.465 55.525 213.545 55.665 ;
        RECT 210.465 55.465 210.785 55.525 ;
        RECT 212.780 55.480 213.070 55.525 ;
        RECT 213.225 55.465 213.545 55.525 ;
        RECT 214.145 55.465 214.465 55.725 ;
        RECT 215.525 55.465 215.845 55.725 ;
        RECT 227.575 55.665 227.715 56.205 ;
        RECT 227.960 56.160 228.250 56.205 ;
        RECT 229.800 56.160 230.090 56.205 ;
        RECT 233.940 56.160 234.230 56.205 ;
        RECT 228.865 55.805 229.185 56.065 ;
        RECT 229.325 55.805 229.645 56.065 ;
        RECT 229.875 56.005 230.015 56.160 ;
        RECT 239.445 56.145 239.765 56.205 ;
        RECT 240.455 56.065 240.595 56.885 ;
        RECT 240.825 56.485 241.145 56.745 ;
        RECT 240.915 56.295 241.055 56.485 ;
        RECT 241.300 56.295 241.590 56.390 ;
        RECT 240.915 56.160 241.590 56.295 ;
        RECT 241.760 56.160 242.050 56.390 ;
        RECT 242.220 56.345 242.510 56.390 ;
        RECT 242.665 56.345 242.985 56.405 ;
        RECT 242.220 56.205 242.985 56.345 ;
        RECT 242.220 56.160 242.510 56.205 ;
        RECT 240.915 56.155 241.515 56.160 ;
        RECT 240.365 56.005 240.685 56.065 ;
        RECT 229.875 55.865 240.685 56.005 ;
        RECT 240.365 55.805 240.685 55.865 ;
        RECT 216.535 55.525 227.715 55.665 ;
        RECT 228.955 55.665 229.095 55.805 ;
        RECT 240.825 55.665 241.145 55.725 ;
        RECT 241.835 55.665 241.975 56.160 ;
        RECT 242.665 56.145 242.985 56.205 ;
        RECT 243.140 56.345 243.430 56.390 ;
        RECT 244.045 56.345 244.365 56.405 ;
        RECT 243.140 56.205 244.365 56.345 ;
        RECT 243.140 56.160 243.430 56.205 ;
        RECT 244.045 56.145 244.365 56.205 ;
        RECT 244.505 56.345 244.825 56.405 ;
        RECT 244.980 56.345 245.270 56.390 ;
        RECT 244.505 56.205 245.270 56.345 ;
        RECT 245.515 56.345 245.655 56.885 ;
        RECT 246.820 56.885 247.585 57.025 ;
        RECT 246.820 56.840 247.110 56.885 ;
        RECT 247.265 56.825 247.585 56.885 ;
        RECT 248.735 56.885 252.630 57.025 ;
        RECT 248.185 56.345 248.505 56.405 ;
        RECT 248.735 56.390 248.875 56.885 ;
        RECT 252.340 56.840 252.630 56.885 ;
        RECT 252.800 57.025 253.090 57.070 ;
        RECT 253.245 57.025 253.565 57.085 ;
        RECT 252.800 56.885 253.565 57.025 ;
        RECT 252.800 56.840 253.090 56.885 ;
        RECT 253.245 56.825 253.565 56.885 ;
        RECT 257.385 56.825 257.705 57.085 ;
        RECT 263.365 56.825 263.685 57.085 ;
        RECT 266.585 57.025 266.905 57.085 ;
        RECT 280.385 57.025 280.705 57.085 ;
        RECT 288.205 57.025 288.525 57.085 ;
        RECT 298.325 57.025 298.645 57.085 ;
        RECT 306.160 57.025 306.450 57.070 ;
        RECT 266.585 56.885 279.695 57.025 ;
        RECT 266.585 56.825 266.905 56.885 ;
        RECT 249.195 56.545 255.315 56.685 ;
        RECT 249.195 56.405 249.335 56.545 ;
        RECT 248.660 56.345 248.950 56.390 ;
        RECT 245.515 56.205 248.950 56.345 ;
        RECT 244.505 56.145 244.825 56.205 ;
        RECT 244.980 56.160 245.270 56.205 ;
        RECT 248.185 56.145 248.505 56.205 ;
        RECT 248.660 56.160 248.950 56.205 ;
        RECT 249.105 56.145 249.425 56.405 ;
        RECT 250.500 56.345 250.790 56.390 ;
        RECT 251.955 56.345 253.015 56.360 ;
        RECT 250.500 56.220 253.015 56.345 ;
        RECT 250.500 56.205 252.095 56.220 ;
        RECT 250.500 56.160 250.790 56.205 ;
        RECT 228.955 55.525 241.975 55.665 ;
        RECT 242.755 55.665 242.895 56.145 ;
        RECT 243.585 56.005 243.905 56.065 ;
        RECT 245.440 56.005 245.730 56.050 ;
        RECT 243.585 55.865 245.730 56.005 ;
        RECT 243.585 55.805 243.905 55.865 ;
        RECT 245.440 55.820 245.730 55.865 ;
        RECT 247.740 55.820 248.030 56.050 ;
        RECT 250.025 56.005 250.345 56.065 ;
        RECT 250.945 56.005 251.265 56.065 ;
        RECT 250.025 55.865 251.265 56.005 ;
        RECT 247.815 55.665 247.955 55.820 ;
        RECT 250.025 55.805 250.345 55.865 ;
        RECT 250.945 55.805 251.265 55.865 ;
        RECT 251.420 55.820 251.710 56.050 ;
        RECT 252.875 56.005 253.015 56.220 ;
        RECT 253.245 56.145 253.565 56.405 ;
        RECT 255.175 56.390 255.315 56.545 ;
        RECT 255.100 56.160 255.390 56.390 ;
        RECT 257.475 56.345 257.615 56.825 ;
        RECT 263.455 56.685 263.595 56.825 ;
        RECT 279.555 56.730 279.695 56.885 ;
        RECT 280.385 56.885 290.735 57.025 ;
        RECT 280.385 56.825 280.705 56.885 ;
        RECT 288.205 56.825 288.525 56.885 ;
        RECT 273.600 56.685 273.890 56.730 ;
        RECT 276.840 56.685 277.490 56.730 ;
        RECT 263.455 56.545 264.975 56.685 ;
        RECT 262.460 56.345 262.750 56.390 ;
        RECT 257.475 56.205 262.750 56.345 ;
        RECT 262.460 56.160 262.750 56.205 ;
        RECT 263.365 56.145 263.685 56.405 ;
        RECT 263.840 56.345 264.130 56.390 ;
        RECT 264.285 56.345 264.605 56.405 ;
        RECT 264.835 56.390 264.975 56.545 ;
        RECT 273.600 56.545 277.490 56.685 ;
        RECT 273.600 56.500 274.190 56.545 ;
        RECT 276.840 56.500 277.490 56.545 ;
        RECT 279.480 56.500 279.770 56.730 ;
        RECT 280.475 56.685 280.615 56.825 ;
        RECT 283.260 56.685 283.550 56.730 ;
        RECT 286.500 56.685 287.150 56.730 ;
        RECT 288.665 56.685 288.985 56.745 ;
        RECT 280.475 56.545 281.075 56.685 ;
        RECT 263.840 56.205 264.605 56.345 ;
        RECT 263.840 56.160 264.130 56.205 ;
        RECT 264.285 56.145 264.605 56.205 ;
        RECT 264.760 56.160 265.050 56.390 ;
        RECT 265.680 56.345 265.970 56.390 ;
        RECT 266.125 56.345 266.445 56.405 ;
        RECT 265.680 56.205 266.445 56.345 ;
        RECT 265.680 56.160 265.970 56.205 ;
        RECT 266.125 56.145 266.445 56.205 ;
        RECT 266.585 56.145 266.905 56.405 ;
        RECT 267.060 56.345 267.350 56.390 ;
        RECT 267.505 56.345 267.825 56.405 ;
        RECT 267.060 56.205 267.825 56.345 ;
        RECT 267.060 56.160 267.350 56.205 ;
        RECT 267.505 56.145 267.825 56.205 ;
        RECT 267.980 56.160 268.270 56.390 ;
        RECT 272.565 56.345 272.885 56.405 ;
        RECT 273.900 56.345 274.190 56.500 ;
        RECT 280.935 56.390 281.075 56.545 ;
        RECT 283.260 56.545 288.985 56.685 ;
        RECT 283.260 56.500 283.850 56.545 ;
        RECT 286.500 56.500 287.150 56.545 ;
        RECT 272.565 56.205 274.190 56.345 ;
        RECT 256.465 56.005 256.785 56.065 ;
        RECT 252.875 55.865 256.785 56.005 ;
        RECT 249.565 55.665 249.885 55.725 ;
        RECT 242.755 55.525 249.885 55.665 ;
        RECT 214.235 55.325 214.375 55.465 ;
        RECT 216.535 55.385 216.675 55.525 ;
        RECT 240.825 55.465 241.145 55.525 ;
        RECT 210.095 55.185 214.375 55.325 ;
        RECT 216.445 55.125 216.765 55.385 ;
        RECT 224.740 55.325 225.030 55.370 ;
        RECT 229.325 55.325 229.645 55.385 ;
        RECT 224.740 55.185 229.645 55.325 ;
        RECT 224.740 55.140 225.030 55.185 ;
        RECT 229.325 55.125 229.645 55.185 ;
        RECT 237.145 55.325 237.465 55.385 ;
        RECT 239.920 55.325 240.210 55.370 ;
        RECT 237.145 55.185 240.210 55.325 ;
        RECT 241.835 55.325 241.975 55.525 ;
        RECT 249.565 55.465 249.885 55.525 ;
        RECT 250.485 55.665 250.805 55.725 ;
        RECT 251.495 55.665 251.635 55.820 ;
        RECT 256.465 55.805 256.785 55.865 ;
        RECT 261.065 56.005 261.385 56.065 ;
        RECT 268.055 56.005 268.195 56.160 ;
        RECT 272.565 56.145 272.885 56.205 ;
        RECT 273.900 56.185 274.190 56.205 ;
        RECT 274.980 56.345 275.270 56.390 ;
        RECT 278.560 56.345 278.850 56.390 ;
        RECT 280.395 56.345 280.685 56.390 ;
        RECT 274.980 56.205 280.685 56.345 ;
        RECT 261.065 55.865 268.195 56.005 ;
        RECT 274.035 56.005 274.175 56.185 ;
        RECT 274.980 56.160 275.270 56.205 ;
        RECT 278.560 56.160 278.850 56.205 ;
        RECT 280.395 56.160 280.685 56.205 ;
        RECT 280.860 56.160 281.150 56.390 ;
        RECT 283.560 56.345 283.850 56.500 ;
        RECT 288.665 56.485 288.985 56.545 ;
        RECT 289.140 56.685 289.430 56.730 ;
        RECT 289.585 56.685 289.905 56.745 ;
        RECT 289.140 56.545 289.905 56.685 ;
        RECT 289.140 56.500 289.430 56.545 ;
        RECT 289.585 56.485 289.905 56.545 ;
        RECT 290.595 56.390 290.735 56.885 ;
        RECT 298.325 56.885 306.450 57.025 ;
        RECT 298.325 56.825 298.645 56.885 ;
        RECT 306.160 56.840 306.450 56.885 ;
        RECT 298.785 56.485 299.105 56.745 ;
        RECT 301.080 56.685 301.730 56.730 ;
        RECT 304.680 56.685 304.970 56.730 ;
        RECT 301.080 56.545 304.970 56.685 ;
        RECT 301.080 56.500 301.730 56.545 ;
        RECT 304.380 56.500 304.970 56.545 ;
        RECT 284.640 56.345 284.930 56.390 ;
        RECT 288.220 56.345 288.510 56.390 ;
        RECT 290.055 56.345 290.345 56.390 ;
        RECT 281.395 56.205 284.295 56.345 ;
        RECT 281.395 56.005 281.535 56.205 ;
        RECT 283.560 56.185 283.850 56.205 ;
        RECT 274.035 55.865 281.535 56.005 ;
        RECT 261.065 55.805 261.385 55.865 ;
        RECT 283.145 55.805 283.465 56.065 ;
        RECT 284.155 56.005 284.295 56.205 ;
        RECT 284.640 56.205 290.345 56.345 ;
        RECT 284.640 56.160 284.930 56.205 ;
        RECT 288.220 56.160 288.510 56.205 ;
        RECT 290.055 56.160 290.345 56.205 ;
        RECT 290.520 56.160 290.810 56.390 ;
        RECT 293.280 56.345 293.570 56.390 ;
        RECT 295.565 56.345 295.885 56.405 ;
        RECT 293.280 56.205 295.885 56.345 ;
        RECT 293.280 56.160 293.570 56.205 ;
        RECT 288.665 56.005 288.985 56.065 ;
        RECT 284.155 55.865 288.985 56.005 ;
        RECT 290.595 56.005 290.735 56.160 ;
        RECT 295.565 56.145 295.885 56.205 ;
        RECT 297.885 56.345 298.175 56.390 ;
        RECT 299.720 56.345 300.010 56.390 ;
        RECT 303.300 56.345 303.590 56.390 ;
        RECT 297.885 56.205 303.590 56.345 ;
        RECT 297.885 56.160 298.175 56.205 ;
        RECT 299.720 56.160 300.010 56.205 ;
        RECT 303.300 56.160 303.590 56.205 ;
        RECT 304.380 56.345 304.670 56.500 ;
        RECT 305.225 56.345 305.545 56.405 ;
        RECT 304.380 56.205 305.545 56.345 ;
        RECT 304.380 56.185 304.670 56.205 ;
        RECT 305.225 56.145 305.545 56.205 ;
        RECT 309.380 56.345 309.670 56.390 ;
        RECT 310.745 56.345 311.065 56.405 ;
        RECT 309.380 56.205 311.065 56.345 ;
        RECT 309.380 56.160 309.670 56.205 ;
        RECT 310.745 56.145 311.065 56.205 ;
        RECT 294.185 56.005 294.505 56.065 ;
        RECT 297.420 56.005 297.710 56.050 ;
        RECT 290.595 55.865 297.710 56.005 ;
        RECT 288.665 55.805 288.985 55.865 ;
        RECT 294.185 55.805 294.505 55.865 ;
        RECT 297.420 55.820 297.710 55.865 ;
        RECT 250.485 55.525 251.635 55.665 ;
        RECT 254.640 55.665 254.930 55.710 ;
        RECT 262.920 55.665 263.210 55.710 ;
        RECT 263.825 55.665 264.145 55.725 ;
        RECT 254.640 55.525 262.215 55.665 ;
        RECT 250.485 55.465 250.805 55.525 ;
        RECT 254.640 55.480 254.930 55.525 ;
        RECT 244.965 55.325 245.285 55.385 ;
        RECT 241.835 55.185 245.285 55.325 ;
        RECT 237.145 55.125 237.465 55.185 ;
        RECT 239.920 55.140 240.210 55.185 ;
        RECT 244.965 55.125 245.285 55.185 ;
        RECT 245.900 55.325 246.190 55.370 ;
        RECT 246.345 55.325 246.665 55.385 ;
        RECT 245.900 55.185 246.665 55.325 ;
        RECT 245.900 55.140 246.190 55.185 ;
        RECT 246.345 55.125 246.665 55.185 ;
        RECT 250.040 55.325 250.330 55.370 ;
        RECT 250.945 55.325 251.265 55.385 ;
        RECT 250.040 55.185 251.265 55.325 ;
        RECT 250.040 55.140 250.330 55.185 ;
        RECT 250.945 55.125 251.265 55.185 ;
        RECT 256.925 55.125 257.245 55.385 ;
        RECT 257.845 55.125 258.165 55.385 ;
        RECT 261.525 55.125 261.845 55.385 ;
        RECT 262.075 55.325 262.215 55.525 ;
        RECT 262.920 55.525 264.145 55.665 ;
        RECT 262.920 55.480 263.210 55.525 ;
        RECT 263.825 55.465 264.145 55.525 ;
        RECT 265.665 55.465 265.985 55.725 ;
        RECT 267.520 55.665 267.810 55.710 ;
        RECT 267.965 55.665 268.285 55.725 ;
        RECT 267.520 55.525 268.285 55.665 ;
        RECT 267.520 55.480 267.810 55.525 ;
        RECT 267.965 55.465 268.285 55.525 ;
        RECT 274.980 55.665 275.270 55.710 ;
        RECT 278.100 55.665 278.390 55.710 ;
        RECT 279.990 55.665 280.280 55.710 ;
        RECT 274.980 55.525 280.280 55.665 ;
        RECT 274.980 55.480 275.270 55.525 ;
        RECT 278.100 55.480 278.390 55.525 ;
        RECT 279.990 55.480 280.280 55.525 ;
        RECT 281.780 55.665 282.070 55.710 ;
        RECT 283.235 55.665 283.375 55.805 ;
        RECT 281.780 55.525 283.375 55.665 ;
        RECT 284.640 55.665 284.930 55.710 ;
        RECT 287.760 55.665 288.050 55.710 ;
        RECT 289.650 55.665 289.940 55.710 ;
        RECT 284.640 55.525 289.940 55.665 ;
        RECT 281.780 55.480 282.070 55.525 ;
        RECT 284.640 55.480 284.930 55.525 ;
        RECT 287.760 55.480 288.050 55.525 ;
        RECT 289.650 55.480 289.940 55.525 ;
        RECT 298.290 55.665 298.580 55.710 ;
        RECT 300.180 55.665 300.470 55.710 ;
        RECT 303.300 55.665 303.590 55.710 ;
        RECT 298.290 55.525 303.590 55.665 ;
        RECT 298.290 55.480 298.580 55.525 ;
        RECT 300.180 55.480 300.470 55.525 ;
        RECT 303.300 55.480 303.590 55.525 ;
        RECT 265.755 55.325 265.895 55.465 ;
        RECT 262.075 55.185 265.895 55.325 ;
        RECT 268.425 55.325 268.745 55.385 ;
        RECT 269.360 55.325 269.650 55.370 ;
        RECT 268.425 55.185 269.650 55.325 ;
        RECT 268.425 55.125 268.745 55.185 ;
        RECT 269.360 55.140 269.650 55.185 ;
        RECT 272.105 55.125 272.425 55.385 ;
        RECT 294.185 55.125 294.505 55.385 ;
        RECT 308.445 55.125 308.765 55.385 ;
        RECT 162.095 54.505 311.135 54.985 ;
        RECT 165.385 54.105 165.705 54.365 ;
        RECT 169.065 54.305 169.385 54.365 ;
        RECT 175.520 54.305 175.810 54.350 ;
        RECT 169.065 54.165 175.810 54.305 ;
        RECT 169.065 54.105 169.385 54.165 ;
        RECT 175.520 54.120 175.810 54.165 ;
        RECT 175.965 54.105 176.285 54.365 ;
        RECT 178.725 54.305 179.045 54.365 ;
        RECT 180.580 54.305 180.870 54.350 ;
        RECT 178.725 54.165 180.870 54.305 ;
        RECT 178.725 54.105 179.045 54.165 ;
        RECT 180.580 54.120 180.870 54.165 ;
        RECT 181.945 54.105 182.265 54.365 ;
        RECT 216.920 54.305 217.210 54.350 ;
        RECT 224.725 54.305 225.045 54.365 ;
        RECT 204.575 54.165 207.705 54.305 ;
        RECT 165.475 53.670 165.615 54.105 ;
        RECT 166.270 53.965 166.560 54.010 ;
        RECT 168.160 53.965 168.450 54.010 ;
        RECT 171.280 53.965 171.570 54.010 ;
        RECT 174.585 53.965 174.905 54.025 ;
        RECT 166.270 53.825 171.570 53.965 ;
        RECT 166.270 53.780 166.560 53.825 ;
        RECT 168.160 53.780 168.450 53.825 ;
        RECT 171.280 53.780 171.570 53.825 ;
        RECT 173.065 53.825 174.905 53.965 ;
        RECT 165.400 53.440 165.690 53.670 ;
        RECT 166.765 53.425 167.085 53.685 ;
        RECT 165.865 53.285 166.155 53.330 ;
        RECT 167.700 53.285 167.990 53.330 ;
        RECT 171.280 53.285 171.570 53.330 ;
        RECT 165.865 53.145 171.570 53.285 ;
        RECT 165.865 53.100 166.155 53.145 ;
        RECT 167.700 53.100 167.990 53.145 ;
        RECT 171.280 53.100 171.570 53.145 ;
        RECT 172.360 53.285 172.650 53.305 ;
        RECT 173.065 53.285 173.205 53.825 ;
        RECT 174.585 53.765 174.905 53.825 ;
        RECT 172.360 53.145 173.205 53.285 ;
        RECT 172.360 52.990 172.650 53.145 ;
        RECT 174.125 53.085 174.445 53.345 ;
        RECT 176.055 53.285 176.195 54.105 ;
        RECT 176.440 53.285 176.730 53.330 ;
        RECT 176.055 53.145 176.730 53.285 ;
        RECT 176.440 53.100 176.730 53.145 ;
        RECT 181.500 53.285 181.790 53.330 ;
        RECT 182.035 53.285 182.175 54.105 ;
        RECT 202.185 53.965 202.505 54.025 ;
        RECT 204.040 53.965 204.330 54.010 ;
        RECT 202.185 53.825 204.330 53.965 ;
        RECT 202.185 53.765 202.505 53.825 ;
        RECT 204.040 53.780 204.330 53.825 ;
        RECT 204.575 53.685 204.715 54.165 ;
        RECT 207.565 53.965 207.705 54.165 ;
        RECT 216.920 54.165 225.045 54.305 ;
        RECT 216.920 54.120 217.210 54.165 ;
        RECT 224.725 54.105 225.045 54.165 ;
        RECT 225.645 54.105 225.965 54.365 ;
        RECT 229.325 54.305 229.645 54.365 ;
        RECT 240.825 54.305 241.145 54.365 ;
        RECT 241.300 54.305 241.590 54.350 ;
        RECT 229.325 54.165 237.835 54.305 ;
        RECT 229.325 54.105 229.645 54.165 ;
        RECT 214.145 53.965 214.465 54.025 ;
        RECT 207.565 53.825 214.465 53.965 ;
        RECT 214.145 53.765 214.465 53.825 ;
        RECT 204.485 53.425 204.805 53.685 ;
        RECT 205.420 53.440 205.710 53.670 ;
        RECT 219.220 53.625 219.510 53.670 ;
        RECT 216.075 53.485 219.510 53.625 ;
        RECT 181.500 53.145 182.175 53.285 ;
        RECT 201.265 53.285 201.585 53.345 ;
        RECT 201.740 53.285 202.030 53.330 ;
        RECT 201.265 53.145 202.030 53.285 ;
        RECT 181.500 53.100 181.790 53.145 ;
        RECT 201.265 53.085 201.585 53.145 ;
        RECT 201.740 53.100 202.030 53.145 ;
        RECT 202.200 53.100 202.490 53.330 ;
        RECT 204.025 53.285 204.345 53.345 ;
        RECT 205.495 53.285 205.635 53.440 ;
        RECT 216.075 53.345 216.215 53.485 ;
        RECT 219.220 53.440 219.510 53.485 ;
        RECT 220.675 53.485 223.575 53.625 ;
        RECT 204.025 53.145 205.635 53.285 ;
        RECT 169.060 52.945 169.710 52.990 ;
        RECT 172.360 52.945 172.950 52.990 ;
        RECT 169.060 52.805 172.950 52.945 ;
        RECT 169.060 52.760 169.710 52.805 ;
        RECT 172.660 52.760 172.950 52.805 ;
        RECT 174.215 52.650 174.355 53.085 ;
        RECT 190.225 52.945 190.545 53.005 ;
        RECT 190.700 52.945 190.990 52.990 ;
        RECT 190.225 52.805 190.990 52.945 ;
        RECT 190.225 52.745 190.545 52.805 ;
        RECT 190.700 52.760 190.990 52.805 ;
        RECT 194.825 52.745 195.145 53.005 ;
        RECT 202.275 52.945 202.415 53.100 ;
        RECT 204.025 53.085 204.345 53.145 ;
        RECT 209.545 53.085 209.865 53.345 ;
        RECT 210.465 53.085 210.785 53.345 ;
        RECT 212.320 53.285 212.610 53.330 ;
        RECT 215.540 53.285 215.830 53.330 ;
        RECT 215.985 53.285 216.305 53.345 ;
        RECT 212.320 53.145 216.305 53.285 ;
        RECT 212.320 53.100 212.610 53.145 ;
        RECT 215.540 53.100 215.830 53.145 ;
        RECT 215.985 53.085 216.305 53.145 ;
        RECT 216.445 53.285 216.765 53.345 ;
        RECT 218.300 53.285 218.590 53.330 ;
        RECT 216.445 53.145 218.590 53.285 ;
        RECT 216.445 53.085 216.765 53.145 ;
        RECT 218.300 53.100 218.590 53.145 ;
        RECT 218.760 53.100 219.050 53.330 ;
        RECT 219.680 53.285 219.970 53.330 ;
        RECT 219.295 53.145 219.970 53.285 ;
        RECT 206.325 52.945 206.645 53.005 ;
        RECT 210.005 52.945 210.325 53.005 ;
        RECT 213.240 52.945 213.530 52.990 ;
        RECT 215.080 52.945 215.370 52.990 ;
        RECT 218.835 52.945 218.975 53.100 ;
        RECT 202.275 52.805 215.370 52.945 ;
        RECT 174.140 52.420 174.430 52.650 ;
        RECT 200.805 52.605 201.125 52.665 ;
        RECT 202.275 52.605 202.415 52.805 ;
        RECT 206.325 52.745 206.645 52.805 ;
        RECT 210.005 52.745 210.325 52.805 ;
        RECT 213.240 52.760 213.530 52.805 ;
        RECT 215.080 52.760 215.370 52.805 ;
        RECT 215.615 52.805 218.975 52.945 ;
        RECT 200.805 52.465 202.415 52.605 ;
        RECT 202.645 52.605 202.965 52.665 ;
        RECT 210.925 52.605 211.245 52.665 ;
        RECT 202.645 52.465 211.245 52.605 ;
        RECT 200.805 52.405 201.125 52.465 ;
        RECT 202.645 52.405 202.965 52.465 ;
        RECT 210.925 52.405 211.245 52.465 ;
        RECT 211.385 52.605 211.705 52.665 ;
        RECT 212.780 52.605 213.070 52.650 ;
        RECT 211.385 52.465 213.070 52.605 ;
        RECT 211.385 52.405 211.705 52.465 ;
        RECT 212.780 52.420 213.070 52.465 ;
        RECT 214.145 52.605 214.465 52.665 ;
        RECT 215.615 52.605 215.755 52.805 ;
        RECT 214.145 52.465 215.755 52.605 ;
        RECT 216.000 52.605 216.290 52.650 ;
        RECT 216.905 52.605 217.225 52.665 ;
        RECT 219.295 52.605 219.435 53.145 ;
        RECT 219.680 53.100 219.970 53.145 ;
        RECT 216.000 52.465 219.435 52.605 ;
        RECT 219.665 52.605 219.985 52.665 ;
        RECT 220.675 52.650 220.815 53.485 ;
        RECT 221.045 53.085 221.365 53.345 ;
        RECT 223.435 53.330 223.575 53.485 ;
        RECT 222.900 53.100 223.190 53.330 ;
        RECT 223.360 53.100 223.650 53.330 ;
        RECT 225.735 53.285 225.875 54.105 ;
        RECT 235.305 53.965 235.625 54.025 ;
        RECT 235.780 53.965 236.070 54.010 ;
        RECT 235.305 53.825 236.070 53.965 ;
        RECT 235.305 53.765 235.625 53.825 ;
        RECT 235.780 53.780 236.070 53.825 ;
        RECT 237.145 53.765 237.465 54.025 ;
        RECT 228.495 53.485 233.695 53.625 ;
        RECT 228.495 53.330 228.635 53.485 ;
        RECT 233.555 53.345 233.695 53.485 ;
        RECT 233.925 53.425 234.245 53.685 ;
        RECT 237.235 53.625 237.375 53.765 ;
        RECT 235.395 53.485 237.375 53.625 ;
        RECT 237.695 53.625 237.835 54.165 ;
        RECT 240.825 54.165 241.590 54.305 ;
        RECT 240.825 54.105 241.145 54.165 ;
        RECT 241.300 54.120 241.590 54.165 ;
        RECT 248.185 54.305 248.505 54.365 ;
        RECT 248.185 54.165 249.335 54.305 ;
        RECT 248.185 54.105 248.505 54.165 ;
        RECT 248.660 53.965 248.950 54.010 ;
        RECT 245.975 53.825 248.950 53.965 ;
        RECT 238.525 53.625 238.845 53.685 ;
        RECT 237.695 53.485 244.735 53.625 ;
        RECT 227.960 53.285 228.250 53.330 ;
        RECT 225.735 53.145 228.250 53.285 ;
        RECT 227.960 53.100 228.250 53.145 ;
        RECT 228.420 53.100 228.710 53.330 ;
        RECT 229.800 53.285 230.090 53.330 ;
        RECT 230.720 53.285 231.010 53.330 ;
        RECT 229.800 53.145 231.010 53.285 ;
        RECT 229.800 53.100 230.090 53.145 ;
        RECT 230.720 53.100 231.010 53.145 ;
        RECT 222.975 52.945 223.115 53.100 ;
        RECT 233.465 53.085 233.785 53.345 ;
        RECT 235.395 53.330 235.535 53.485 ;
        RECT 235.320 53.100 235.610 53.330 ;
        RECT 235.765 53.085 236.085 53.345 ;
        RECT 236.240 53.100 236.530 53.330 ;
        RECT 236.700 53.285 236.990 53.330 ;
        RECT 237.145 53.285 237.465 53.345 ;
        RECT 237.695 53.330 237.835 53.485 ;
        RECT 238.525 53.425 238.845 53.485 ;
        RECT 236.700 53.145 237.465 53.285 ;
        RECT 236.700 53.100 236.990 53.145 ;
        RECT 235.855 52.945 235.995 53.085 ;
        RECT 222.975 52.805 235.995 52.945 ;
        RECT 236.315 52.945 236.455 53.100 ;
        RECT 237.145 53.085 237.465 53.145 ;
        RECT 237.620 53.100 237.910 53.330 ;
        RECT 238.065 53.085 238.385 53.345 ;
        RECT 239.445 53.085 239.765 53.345 ;
        RECT 240.365 53.085 240.685 53.345 ;
        RECT 240.825 53.285 241.145 53.345 ;
        RECT 241.745 53.285 242.065 53.345 ;
        RECT 240.825 53.145 242.065 53.285 ;
        RECT 240.825 53.085 241.145 53.145 ;
        RECT 241.745 53.085 242.065 53.145 ;
        RECT 244.045 53.085 244.365 53.345 ;
        RECT 238.155 52.945 238.295 53.085 ;
        RECT 236.315 52.805 238.295 52.945 ;
        RECT 220.600 52.605 220.890 52.650 ;
        RECT 219.665 52.465 220.890 52.605 ;
        RECT 214.145 52.405 214.465 52.465 ;
        RECT 216.000 52.420 216.290 52.465 ;
        RECT 216.905 52.405 217.225 52.465 ;
        RECT 219.665 52.405 219.985 52.465 ;
        RECT 220.600 52.420 220.890 52.465 ;
        RECT 226.565 52.605 226.885 52.665 ;
        RECT 227.040 52.605 227.330 52.650 ;
        RECT 226.565 52.465 227.330 52.605 ;
        RECT 226.565 52.405 226.885 52.465 ;
        RECT 227.040 52.420 227.330 52.465 ;
        RECT 234.385 52.405 234.705 52.665 ;
        RECT 238.065 52.405 238.385 52.665 ;
        RECT 239.535 52.605 239.675 53.085 ;
        RECT 239.920 52.945 240.210 52.990 ;
        RECT 244.135 52.945 244.275 53.085 ;
        RECT 239.920 52.805 244.275 52.945 ;
        RECT 244.595 52.945 244.735 53.485 ;
        RECT 244.965 53.425 245.285 53.685 ;
        RECT 245.975 53.330 246.115 53.825 ;
        RECT 248.660 53.780 248.950 53.825 ;
        RECT 246.345 53.425 246.665 53.685 ;
        RECT 246.805 53.425 247.125 53.685 ;
        RECT 249.195 53.625 249.335 54.165 ;
        RECT 249.565 54.105 249.885 54.365 ;
        RECT 253.260 54.305 253.550 54.350 ;
        RECT 256.465 54.305 256.785 54.365 ;
        RECT 271.200 54.305 271.490 54.350 ;
        RECT 253.260 54.165 256.785 54.305 ;
        RECT 253.260 54.120 253.550 54.165 ;
        RECT 256.465 54.105 256.785 54.165 ;
        RECT 260.695 54.165 271.490 54.305 ;
        RECT 251.420 53.965 251.710 54.010 ;
        RECT 256.925 53.965 257.245 54.025 ;
        RECT 251.420 53.825 257.245 53.965 ;
        RECT 251.420 53.780 251.710 53.825 ;
        RECT 256.925 53.765 257.245 53.825 ;
        RECT 249.195 53.485 253.015 53.625 ;
        RECT 245.900 53.100 246.190 53.330 ;
        RECT 247.265 53.085 247.585 53.345 ;
        RECT 252.875 53.330 253.015 53.485 ;
        RECT 253.245 53.425 253.565 53.685 ;
        RECT 248.200 53.285 248.490 53.330 ;
        RECT 248.200 53.145 252.555 53.285 ;
        RECT 248.200 53.100 248.490 53.145 ;
        RECT 248.275 52.945 248.415 53.100 ;
        RECT 244.595 52.805 248.415 52.945 ;
        RECT 249.105 52.945 249.425 53.005 ;
        RECT 249.580 52.945 249.870 52.990 ;
        RECT 249.105 52.805 249.870 52.945 ;
        RECT 239.920 52.760 240.210 52.805 ;
        RECT 249.105 52.745 249.425 52.805 ;
        RECT 249.580 52.760 249.870 52.805 ;
        RECT 251.865 52.745 252.185 53.005 ;
        RECT 252.415 52.945 252.555 53.145 ;
        RECT 252.830 53.100 253.120 53.330 ;
        RECT 253.335 53.285 253.475 53.425 ;
        RECT 260.695 53.330 260.835 54.165 ;
        RECT 271.200 54.120 271.490 54.165 ;
        RECT 302.925 54.305 303.245 54.365 ;
        RECT 303.400 54.305 303.690 54.350 ;
        RECT 307.065 54.305 307.385 54.365 ;
        RECT 302.925 54.165 307.385 54.305 ;
        RECT 302.925 54.105 303.245 54.165 ;
        RECT 303.400 54.120 303.690 54.165 ;
        RECT 307.065 54.105 307.385 54.165 ;
        RECT 261.065 53.765 261.385 54.025 ;
        RECT 261.525 53.765 261.845 54.025 ;
        RECT 262.870 53.965 263.160 54.010 ;
        RECT 264.760 53.965 265.050 54.010 ;
        RECT 267.880 53.965 268.170 54.010 ;
        RECT 262.870 53.825 268.170 53.965 ;
        RECT 262.870 53.780 263.160 53.825 ;
        RECT 264.760 53.780 265.050 53.825 ;
        RECT 267.880 53.780 268.170 53.825 ;
        RECT 270.725 53.765 271.045 54.025 ;
        RECT 295.530 53.965 295.820 54.010 ;
        RECT 297.420 53.965 297.710 54.010 ;
        RECT 300.540 53.965 300.830 54.010 ;
        RECT 295.530 53.825 300.830 53.965 ;
        RECT 295.530 53.780 295.820 53.825 ;
        RECT 297.420 53.780 297.710 53.825 ;
        RECT 300.540 53.780 300.830 53.825 ;
        RECT 253.720 53.285 254.010 53.330 ;
        RECT 253.335 53.145 254.010 53.285 ;
        RECT 253.720 53.100 254.010 53.145 ;
        RECT 260.620 53.100 260.910 53.330 ;
        RECT 261.155 53.285 261.295 53.765 ;
        RECT 261.615 53.625 261.755 53.765 ;
        RECT 263.380 53.625 263.670 53.670 ;
        RECT 261.615 53.485 263.670 53.625 ;
        RECT 263.380 53.440 263.670 53.485 ;
        RECT 272.105 53.625 272.425 53.685 ;
        RECT 294.660 53.625 294.950 53.670 ;
        RECT 272.105 53.485 282.915 53.625 ;
        RECT 272.105 53.425 272.425 53.485 ;
        RECT 261.540 53.285 261.830 53.330 ;
        RECT 261.155 53.145 261.830 53.285 ;
        RECT 261.540 53.100 261.830 53.145 ;
        RECT 262.000 53.100 262.290 53.330 ;
        RECT 262.465 53.285 262.755 53.330 ;
        RECT 264.300 53.285 264.590 53.330 ;
        RECT 267.880 53.285 268.170 53.330 ;
        RECT 262.465 53.145 268.170 53.285 ;
        RECT 262.465 53.100 262.755 53.145 ;
        RECT 264.300 53.100 264.590 53.145 ;
        RECT 267.880 53.100 268.170 53.145 ;
        RECT 259.700 52.945 259.990 52.990 ;
        RECT 252.415 52.805 259.990 52.945 ;
        RECT 262.075 52.945 262.215 53.100 ;
        RECT 265.665 52.990 265.985 53.005 ;
        RECT 268.960 52.990 269.250 53.305 ;
        RECT 274.420 53.285 274.710 53.330 ;
        RECT 274.865 53.285 275.185 53.345 ;
        RECT 274.420 53.145 275.185 53.285 ;
        RECT 274.420 53.100 274.710 53.145 ;
        RECT 274.865 53.085 275.185 53.145 ;
        RECT 278.085 53.085 278.405 53.345 ;
        RECT 281.305 53.085 281.625 53.345 ;
        RECT 281.780 53.100 282.070 53.330 ;
        RECT 282.775 53.285 282.915 53.485 ;
        RECT 288.295 53.485 294.950 53.625 ;
        RECT 288.295 53.345 288.435 53.485 ;
        RECT 294.660 53.440 294.950 53.485 ;
        RECT 284.540 53.285 284.830 53.330 ;
        RECT 285.905 53.285 286.225 53.345 ;
        RECT 282.775 53.145 283.605 53.285 ;
        RECT 265.660 52.945 266.310 52.990 ;
        RECT 268.960 52.945 269.550 52.990 ;
        RECT 262.075 52.805 262.675 52.945 ;
        RECT 259.700 52.760 259.990 52.805 ;
        RECT 251.955 52.605 252.095 52.745 ;
        RECT 239.535 52.465 252.095 52.605 ;
        RECT 259.775 52.605 259.915 52.760 ;
        RECT 261.985 52.605 262.305 52.665 ;
        RECT 259.775 52.465 262.305 52.605 ;
        RECT 262.535 52.605 262.675 52.805 ;
        RECT 265.660 52.805 269.550 52.945 ;
        RECT 278.175 52.945 278.315 53.085 ;
        RECT 281.855 52.945 281.995 53.100 ;
        RECT 278.175 52.805 281.995 52.945 ;
        RECT 265.660 52.760 266.310 52.805 ;
        RECT 269.260 52.760 269.550 52.805 ;
        RECT 265.665 52.745 265.985 52.760 ;
        RECT 265.205 52.605 265.525 52.665 ;
        RECT 262.535 52.465 265.525 52.605 ;
        RECT 261.985 52.405 262.305 52.465 ;
        RECT 265.205 52.405 265.525 52.465 ;
        RECT 280.385 52.405 280.705 52.665 ;
        RECT 283.465 52.605 283.605 53.145 ;
        RECT 284.540 53.145 286.225 53.285 ;
        RECT 284.540 53.100 284.830 53.145 ;
        RECT 285.905 53.085 286.225 53.145 ;
        RECT 288.205 53.085 288.525 53.345 ;
        RECT 292.360 53.100 292.650 53.330 ;
        RECT 293.280 53.285 293.570 53.330 ;
        RECT 293.725 53.285 294.045 53.345 ;
        RECT 293.280 53.145 294.045 53.285 ;
        RECT 293.280 53.100 293.570 53.145 ;
        RECT 288.665 52.745 288.985 53.005 ;
        RECT 292.435 52.945 292.575 53.100 ;
        RECT 293.725 53.085 294.045 53.145 ;
        RECT 294.185 53.085 294.505 53.345 ;
        RECT 295.125 53.285 295.415 53.330 ;
        RECT 296.960 53.285 297.250 53.330 ;
        RECT 300.540 53.285 300.830 53.330 ;
        RECT 295.125 53.145 300.830 53.285 ;
        RECT 295.125 53.100 295.415 53.145 ;
        RECT 296.960 53.100 297.250 53.145 ;
        RECT 300.540 53.100 300.830 53.145 ;
        RECT 289.215 52.805 292.575 52.945 ;
        RECT 294.275 52.945 294.415 53.085 ;
        RECT 298.325 52.990 298.645 53.005 ;
        RECT 301.620 52.990 301.910 53.305 ;
        RECT 308.905 53.085 309.225 53.345 ;
        RECT 296.040 52.945 296.330 52.990 ;
        RECT 294.275 52.805 296.330 52.945 ;
        RECT 289.215 52.605 289.355 52.805 ;
        RECT 296.040 52.760 296.330 52.805 ;
        RECT 298.320 52.945 298.970 52.990 ;
        RECT 301.620 52.945 302.210 52.990 ;
        RECT 298.320 52.805 302.210 52.945 ;
        RECT 298.320 52.760 298.970 52.805 ;
        RECT 301.920 52.760 302.210 52.805 ;
        RECT 298.325 52.745 298.645 52.760 ;
        RECT 283.465 52.465 289.355 52.605 ;
        RECT 290.965 52.605 291.285 52.665 ;
        RECT 291.440 52.605 291.730 52.650 ;
        RECT 290.965 52.465 291.730 52.605 ;
        RECT 290.965 52.405 291.285 52.465 ;
        RECT 291.440 52.420 291.730 52.465 ;
        RECT 306.160 52.605 306.450 52.650 ;
        RECT 307.065 52.605 307.385 52.665 ;
        RECT 306.160 52.465 307.385 52.605 ;
        RECT 306.160 52.420 306.450 52.465 ;
        RECT 307.065 52.405 307.385 52.465 ;
        RECT 162.095 51.785 311.935 52.265 ;
        RECT 203.105 51.585 203.425 51.645 ;
        RECT 204.500 51.585 204.790 51.630 ;
        RECT 203.105 51.445 204.790 51.585 ;
        RECT 203.105 51.385 203.425 51.445 ;
        RECT 204.500 51.400 204.790 51.445 ;
        RECT 207.245 51.385 207.565 51.645 ;
        RECT 208.165 51.585 208.485 51.645 ;
        RECT 211.385 51.585 211.705 51.645 ;
        RECT 208.165 51.445 211.705 51.585 ;
        RECT 208.165 51.385 208.485 51.445 ;
        RECT 211.385 51.385 211.705 51.445 ;
        RECT 212.305 51.385 212.625 51.645 ;
        RECT 215.525 51.585 215.845 51.645 ;
        RECT 217.380 51.585 217.670 51.630 ;
        RECT 242.205 51.585 242.525 51.645 ;
        RECT 215.525 51.445 217.670 51.585 ;
        RECT 215.525 51.385 215.845 51.445 ;
        RECT 217.380 51.400 217.670 51.445 ;
        RECT 222.515 51.445 256.005 51.585 ;
        RECT 187.925 51.245 188.245 51.305 ;
        RECT 190.240 51.245 190.530 51.290 ;
        RECT 190.685 51.245 191.005 51.305 ;
        RECT 187.925 51.105 191.005 51.245 ;
        RECT 187.925 51.045 188.245 51.105 ;
        RECT 190.240 51.060 190.530 51.105 ;
        RECT 190.685 51.045 191.005 51.105 ;
        RECT 194.380 51.245 194.670 51.290 ;
        RECT 194.825 51.245 195.145 51.305 ;
        RECT 194.380 51.105 220.355 51.245 ;
        RECT 194.380 51.060 194.670 51.105 ;
        RECT 194.825 51.045 195.145 51.105 ;
        RECT 220.215 50.965 220.355 51.105 ;
        RECT 198.980 50.905 199.270 50.950 ;
        RECT 207.720 50.905 208.010 50.950 ;
        RECT 210.005 50.905 210.325 50.965 ;
        RECT 210.480 50.905 210.770 50.950 ;
        RECT 198.980 50.765 205.635 50.905 ;
        RECT 198.980 50.720 199.270 50.765 ;
        RECT 201.265 50.565 201.585 50.625 ;
        RECT 200.435 50.425 201.585 50.565 ;
        RECT 192.985 50.225 193.305 50.285 ;
        RECT 200.435 50.270 200.575 50.425 ;
        RECT 201.265 50.365 201.585 50.425 ;
        RECT 203.105 50.565 203.425 50.625 ;
        RECT 204.485 50.565 204.805 50.625 ;
        RECT 203.105 50.425 204.805 50.565 ;
        RECT 203.105 50.365 203.425 50.425 ;
        RECT 204.485 50.365 204.805 50.425 ;
        RECT 200.360 50.225 200.650 50.270 ;
        RECT 192.985 50.085 200.650 50.225 ;
        RECT 192.985 50.025 193.305 50.085 ;
        RECT 200.360 50.040 200.650 50.085 ;
        RECT 200.805 50.225 201.125 50.285 ;
        RECT 205.495 50.270 205.635 50.765 ;
        RECT 207.720 50.765 209.340 50.905 ;
        RECT 207.720 50.720 208.010 50.765 ;
        RECT 208.180 50.380 208.470 50.610 ;
        RECT 202.660 50.225 202.950 50.270 ;
        RECT 200.805 50.085 202.950 50.225 ;
        RECT 200.805 50.025 201.125 50.085 ;
        RECT 202.660 50.040 202.950 50.085 ;
        RECT 205.420 50.040 205.710 50.270 ;
        RECT 206.785 50.225 207.105 50.285 ;
        RECT 208.255 50.225 208.395 50.380 ;
        RECT 206.785 50.085 208.395 50.225 ;
        RECT 209.200 50.225 209.340 50.765 ;
        RECT 210.005 50.765 210.770 50.905 ;
        RECT 210.005 50.705 210.325 50.765 ;
        RECT 210.480 50.720 210.770 50.765 ;
        RECT 210.925 50.705 211.245 50.965 ;
        RECT 214.145 50.705 214.465 50.965 ;
        RECT 216.585 50.905 216.875 50.950 ;
        RECT 216.535 50.720 216.875 50.905 ;
        RECT 220.125 50.905 220.445 50.965 ;
        RECT 222.515 50.950 222.655 51.445 ;
        RECT 242.205 51.385 242.525 51.445 ;
        RECT 226.120 51.245 226.410 51.290 ;
        RECT 226.565 51.245 226.885 51.305 ;
        RECT 226.120 51.105 226.885 51.245 ;
        RECT 226.120 51.060 226.410 51.105 ;
        RECT 226.565 51.045 226.885 51.105 ;
        RECT 227.485 51.245 227.805 51.305 ;
        RECT 228.400 51.245 229.050 51.290 ;
        RECT 232.000 51.245 232.290 51.290 ;
        RECT 245.440 51.245 245.730 51.290 ;
        RECT 227.485 51.105 232.290 51.245 ;
        RECT 227.485 51.045 227.805 51.105 ;
        RECT 228.400 51.060 229.050 51.105 ;
        RECT 231.700 51.060 232.290 51.105 ;
        RECT 236.315 51.105 245.730 51.245 ;
        RECT 255.865 51.245 256.005 51.445 ;
        RECT 260.605 51.385 260.925 51.645 ;
        RECT 268.885 51.585 269.205 51.645 ;
        RECT 262.535 51.445 284.755 51.585 ;
        RECT 259.240 51.245 259.530 51.290 ;
        RECT 262.535 51.245 262.675 51.445 ;
        RECT 268.885 51.385 269.205 51.445 ;
        RECT 255.865 51.105 262.675 51.245 ;
        RECT 222.440 50.905 222.730 50.950 ;
        RECT 220.125 50.765 222.730 50.905 ;
        RECT 209.545 50.565 209.865 50.625 ;
        RECT 214.235 50.565 214.375 50.705 ;
        RECT 215.540 50.565 215.830 50.610 ;
        RECT 209.545 50.425 214.375 50.565 ;
        RECT 214.695 50.425 215.830 50.565 ;
        RECT 209.545 50.365 209.865 50.425 ;
        RECT 210.005 50.225 210.325 50.285 ;
        RECT 214.695 50.225 214.835 50.425 ;
        RECT 215.540 50.380 215.830 50.425 ;
        RECT 215.985 50.365 216.305 50.625 ;
        RECT 209.200 50.085 209.775 50.225 ;
        RECT 206.785 50.025 207.105 50.085 ;
        RECT 199.900 49.885 200.190 49.930 ;
        RECT 201.265 49.885 201.585 49.945 ;
        RECT 199.900 49.745 201.585 49.885 ;
        RECT 199.900 49.700 200.190 49.745 ;
        RECT 201.265 49.685 201.585 49.745 ;
        RECT 202.185 49.685 202.505 49.945 ;
        RECT 209.635 49.885 209.775 50.085 ;
        RECT 210.005 50.085 214.835 50.225 ;
        RECT 215.065 50.225 215.385 50.285 ;
        RECT 216.535 50.225 216.675 50.720 ;
        RECT 220.125 50.705 220.445 50.765 ;
        RECT 222.440 50.720 222.730 50.765 ;
        RECT 225.205 50.905 225.495 50.950 ;
        RECT 227.040 50.905 227.330 50.950 ;
        RECT 230.620 50.905 230.910 50.950 ;
        RECT 225.205 50.765 230.910 50.905 ;
        RECT 225.205 50.720 225.495 50.765 ;
        RECT 227.040 50.720 227.330 50.765 ;
        RECT 230.620 50.720 230.910 50.765 ;
        RECT 231.700 50.745 231.990 51.060 ;
        RECT 236.315 50.950 236.455 51.105 ;
        RECT 245.440 51.060 245.730 51.105 ;
        RECT 259.240 51.060 259.530 51.105 ;
        RECT 262.905 51.045 263.225 51.305 ;
        RECT 267.060 51.245 267.350 51.290 ;
        RECT 268.425 51.245 268.745 51.305 ;
        RECT 269.345 51.290 269.665 51.305 ;
        RECT 284.615 51.290 284.755 51.445 ;
        RECT 295.565 51.385 295.885 51.645 ;
        RECT 297.420 51.585 297.710 51.630 ;
        RECT 302.925 51.585 303.245 51.645 ;
        RECT 308.905 51.630 309.225 51.645 ;
        RECT 297.420 51.445 303.245 51.585 ;
        RECT 297.420 51.400 297.710 51.445 ;
        RECT 302.925 51.385 303.245 51.445 ;
        RECT 308.690 51.400 309.225 51.630 ;
        RECT 308.905 51.385 309.225 51.400 ;
        RECT 267.060 51.105 268.745 51.245 ;
        RECT 267.060 51.060 267.350 51.105 ;
        RECT 268.425 51.045 268.745 51.105 ;
        RECT 269.340 51.245 269.990 51.290 ;
        RECT 272.940 51.245 273.230 51.290 ;
        RECT 282.240 51.245 282.530 51.290 ;
        RECT 269.340 51.105 273.230 51.245 ;
        RECT 269.340 51.060 269.990 51.105 ;
        RECT 272.640 51.060 273.230 51.105 ;
        RECT 279.555 51.105 282.530 51.245 ;
        RECT 269.345 51.045 269.665 51.060 ;
        RECT 236.240 50.720 236.530 50.950 ;
        RECT 237.620 50.720 237.910 50.950 ;
        RECT 218.760 50.565 219.050 50.610 ;
        RECT 219.665 50.565 219.985 50.625 ;
        RECT 224.740 50.565 225.030 50.610 ;
        RECT 218.760 50.425 225.030 50.565 ;
        RECT 237.695 50.565 237.835 50.720 ;
        RECT 238.065 50.705 238.385 50.965 ;
        RECT 241.285 50.705 241.605 50.965 ;
        RECT 243.125 50.905 243.445 50.965 ;
        RECT 257.845 50.905 258.165 50.965 ;
        RECT 260.325 50.905 260.615 50.950 ;
        RECT 243.125 50.765 253.935 50.905 ;
        RECT 243.125 50.705 243.445 50.765 ;
        RECT 241.375 50.565 241.515 50.705 ;
        RECT 253.795 50.625 253.935 50.765 ;
        RECT 257.845 50.765 260.615 50.905 ;
        RECT 257.845 50.705 258.165 50.765 ;
        RECT 260.325 50.720 260.615 50.765 ;
        RECT 262.460 50.905 262.750 50.950 ;
        RECT 262.995 50.905 263.135 51.045 ;
        RECT 262.460 50.765 263.135 50.905 ;
        RECT 266.145 50.905 266.435 50.950 ;
        RECT 267.980 50.905 268.270 50.950 ;
        RECT 271.560 50.905 271.850 50.950 ;
        RECT 266.145 50.765 271.850 50.905 ;
        RECT 262.460 50.720 262.750 50.765 ;
        RECT 266.145 50.720 266.435 50.765 ;
        RECT 267.980 50.720 268.270 50.765 ;
        RECT 271.560 50.720 271.850 50.765 ;
        RECT 272.640 50.745 272.930 51.060 ;
        RECT 279.555 50.965 279.695 51.105 ;
        RECT 282.240 51.060 282.530 51.105 ;
        RECT 284.540 51.245 284.830 51.290 ;
        RECT 285.905 51.245 286.225 51.305 ;
        RECT 284.540 51.105 286.225 51.245 ;
        RECT 284.540 51.060 284.830 51.105 ;
        RECT 285.905 51.045 286.225 51.105 ;
        RECT 288.205 51.245 288.525 51.305 ;
        RECT 294.185 51.245 294.505 51.305 ;
        RECT 300.645 51.245 300.935 51.290 ;
        RECT 302.505 51.245 302.795 51.290 ;
        RECT 288.205 51.105 299.935 51.245 ;
        RECT 288.205 51.045 288.525 51.105 ;
        RECT 294.185 51.045 294.505 51.105 ;
        RECT 275.800 50.905 276.090 50.950 ;
        RECT 273.115 50.765 276.090 50.905 ;
        RECT 237.695 50.425 241.515 50.565 ;
        RECT 218.760 50.380 219.050 50.425 ;
        RECT 219.665 50.365 219.985 50.425 ;
        RECT 224.740 50.380 225.030 50.425 ;
        RECT 248.660 50.380 248.950 50.610 ;
        RECT 216.905 50.225 217.225 50.285 ;
        RECT 215.065 50.085 217.225 50.225 ;
        RECT 210.005 50.025 210.325 50.085 ;
        RECT 215.065 50.025 215.385 50.085 ;
        RECT 216.905 50.025 217.225 50.085 ;
        RECT 220.585 50.025 220.905 50.285 ;
        RECT 225.610 50.225 225.900 50.270 ;
        RECT 227.500 50.225 227.790 50.270 ;
        RECT 230.620 50.225 230.910 50.270 ;
        RECT 225.610 50.085 230.910 50.225 ;
        RECT 225.610 50.040 225.900 50.085 ;
        RECT 227.500 50.040 227.790 50.085 ;
        RECT 230.620 50.040 230.910 50.085 ;
        RECT 233.480 50.225 233.770 50.270 ;
        RECT 233.925 50.225 234.245 50.285 ;
        RECT 233.480 50.085 234.245 50.225 ;
        RECT 233.480 50.040 233.770 50.085 ;
        RECT 233.925 50.025 234.245 50.085 ;
        RECT 237.605 50.225 237.925 50.285 ;
        RECT 239.920 50.225 240.210 50.270 ;
        RECT 237.605 50.085 240.210 50.225 ;
        RECT 237.605 50.025 237.925 50.085 ;
        RECT 239.920 50.040 240.210 50.085 ;
        RECT 247.725 50.225 248.045 50.285 ;
        RECT 248.735 50.225 248.875 50.380 ;
        RECT 253.705 50.365 254.025 50.625 ;
        RECT 255.560 50.565 255.850 50.610 ;
        RECT 256.925 50.565 257.245 50.625 ;
        RECT 255.560 50.425 257.245 50.565 ;
        RECT 255.560 50.380 255.850 50.425 ;
        RECT 256.925 50.365 257.245 50.425 ;
        RECT 262.905 50.365 263.225 50.625 ;
        RECT 265.205 50.565 265.525 50.625 ;
        RECT 265.680 50.565 265.970 50.610 ;
        RECT 265.205 50.425 265.970 50.565 ;
        RECT 265.205 50.365 265.525 50.425 ;
        RECT 265.680 50.380 265.970 50.425 ;
        RECT 270.725 50.565 271.045 50.625 ;
        RECT 273.115 50.565 273.255 50.765 ;
        RECT 275.800 50.720 276.090 50.765 ;
        RECT 277.255 50.765 278.315 50.905 ;
        RECT 270.725 50.425 273.255 50.565 ;
        RECT 274.880 50.565 275.170 50.610 ;
        RECT 277.255 50.565 277.395 50.765 ;
        RECT 278.175 50.625 278.315 50.765 ;
        RECT 279.465 50.705 279.785 50.965 ;
        RECT 280.385 50.905 280.705 50.965 ;
        RECT 299.795 50.950 299.935 51.105 ;
        RECT 300.645 51.105 302.795 51.245 ;
        RECT 300.645 51.060 300.935 51.105 ;
        RECT 302.505 51.060 302.795 51.105 ;
        RECT 303.425 51.245 303.715 51.290 ;
        RECT 305.225 51.245 305.545 51.305 ;
        RECT 306.685 51.245 306.975 51.290 ;
        RECT 303.425 51.105 306.975 51.245 ;
        RECT 303.425 51.060 303.715 51.105 ;
        RECT 280.860 50.905 281.150 50.950 ;
        RECT 280.385 50.765 281.150 50.905 ;
        RECT 280.385 50.705 280.705 50.765 ;
        RECT 280.860 50.720 281.150 50.765 ;
        RECT 281.325 50.720 281.615 50.950 ;
        RECT 282.700 50.720 282.990 50.950 ;
        RECT 283.185 50.720 283.475 50.950 ;
        RECT 299.720 50.720 300.010 50.950 ;
        RECT 301.560 50.720 301.850 50.950 ;
        RECT 302.580 50.905 302.795 51.060 ;
        RECT 305.225 51.045 305.545 51.105 ;
        RECT 306.685 51.060 306.975 51.105 ;
        RECT 304.825 50.905 305.115 50.950 ;
        RECT 302.580 50.765 305.115 50.905 ;
        RECT 304.825 50.720 305.115 50.765 ;
        RECT 274.880 50.425 277.395 50.565 ;
        RECT 270.725 50.365 271.045 50.425 ;
        RECT 274.880 50.380 275.170 50.425 ;
        RECT 277.625 50.365 277.945 50.625 ;
        RECT 278.085 50.365 278.405 50.625 ;
        RECT 281.395 50.565 281.535 50.720 ;
        RECT 280.475 50.425 281.535 50.565 ;
        RECT 266.550 50.225 266.840 50.270 ;
        RECT 268.440 50.225 268.730 50.270 ;
        RECT 271.560 50.225 271.850 50.270 ;
        RECT 247.725 50.085 266.355 50.225 ;
        RECT 247.725 50.025 248.045 50.085 ;
        RECT 220.675 49.885 220.815 50.025 ;
        RECT 209.635 49.745 220.815 49.885 ;
        RECT 221.505 49.885 221.825 49.945 ;
        RECT 227.945 49.885 228.265 49.945 ;
        RECT 221.505 49.745 228.265 49.885 ;
        RECT 221.505 49.685 221.825 49.745 ;
        RECT 227.945 49.685 228.265 49.745 ;
        RECT 236.700 49.885 236.990 49.930 ;
        RECT 238.525 49.885 238.845 49.945 ;
        RECT 236.700 49.745 238.845 49.885 ;
        RECT 236.700 49.700 236.990 49.745 ;
        RECT 238.525 49.685 238.845 49.745 ;
        RECT 239.000 49.885 239.290 49.930 ;
        RECT 240.365 49.885 240.685 49.945 ;
        RECT 239.000 49.745 240.685 49.885 ;
        RECT 239.000 49.700 239.290 49.745 ;
        RECT 240.365 49.685 240.685 49.745 ;
        RECT 259.685 49.685 260.005 49.945 ;
        RECT 266.215 49.885 266.355 50.085 ;
        RECT 266.550 50.085 271.850 50.225 ;
        RECT 266.550 50.040 266.840 50.085 ;
        RECT 268.440 50.040 268.730 50.085 ;
        RECT 271.560 50.040 271.850 50.085 ;
        RECT 273.485 50.225 273.805 50.285 ;
        RECT 280.475 50.270 280.615 50.425 ;
        RECT 273.485 50.085 280.155 50.225 ;
        RECT 273.485 50.025 273.805 50.085 ;
        RECT 269.805 49.885 270.125 49.945 ;
        RECT 266.215 49.745 270.125 49.885 ;
        RECT 269.805 49.685 270.125 49.745 ;
        RECT 270.265 49.885 270.585 49.945 ;
        RECT 274.420 49.885 274.710 49.930 ;
        RECT 274.865 49.885 275.185 49.945 ;
        RECT 270.265 49.745 275.185 49.885 ;
        RECT 270.265 49.685 270.585 49.745 ;
        RECT 274.420 49.700 274.710 49.745 ;
        RECT 274.865 49.685 275.185 49.745 ;
        RECT 276.705 49.685 277.025 49.945 ;
        RECT 280.015 49.885 280.155 50.085 ;
        RECT 280.400 50.040 280.690 50.270 ;
        RECT 282.225 49.885 282.545 49.945 ;
        RECT 280.015 49.745 282.545 49.885 ;
        RECT 282.775 49.885 282.915 50.720 ;
        RECT 283.235 50.285 283.375 50.720 ;
        RECT 291.440 50.380 291.730 50.610 ;
        RECT 283.145 50.025 283.465 50.285 ;
        RECT 284.080 50.225 284.370 50.270 ;
        RECT 291.515 50.225 291.655 50.380 ;
        RECT 297.865 50.365 298.185 50.625 ;
        RECT 298.340 50.380 298.630 50.610 ;
        RECT 301.635 50.565 301.775 50.720 ;
        RECT 305.685 50.565 306.005 50.625 ;
        RECT 301.635 50.425 306.005 50.565 ;
        RECT 284.080 50.085 291.655 50.225 ;
        RECT 295.105 50.225 295.425 50.285 ;
        RECT 298.415 50.225 298.555 50.380 ;
        RECT 305.685 50.365 306.005 50.425 ;
        RECT 295.105 50.085 298.555 50.225 ;
        RECT 300.185 50.225 300.475 50.270 ;
        RECT 302.045 50.225 302.335 50.270 ;
        RECT 304.825 50.225 305.115 50.270 ;
        RECT 300.185 50.085 305.115 50.225 ;
        RECT 284.080 50.040 284.370 50.085 ;
        RECT 295.105 50.025 295.425 50.085 ;
        RECT 300.185 50.040 300.475 50.085 ;
        RECT 302.045 50.040 302.335 50.085 ;
        RECT 304.825 50.040 305.115 50.085 ;
        RECT 285.445 49.885 285.765 49.945 ;
        RECT 282.775 49.745 285.765 49.885 ;
        RECT 282.225 49.685 282.545 49.745 ;
        RECT 285.445 49.685 285.765 49.745 ;
        RECT 294.645 49.685 294.965 49.945 ;
        RECT 162.095 49.065 311.135 49.545 ;
        RECT 201.725 48.865 202.045 48.925 ;
        RECT 204.945 48.865 205.265 48.925 ;
        RECT 189.855 48.725 201.495 48.865 ;
        RECT 177.820 48.525 178.110 48.570 ;
        RECT 180.530 48.525 180.820 48.570 ;
        RECT 182.420 48.525 182.710 48.570 ;
        RECT 185.540 48.525 185.830 48.570 ;
        RECT 177.820 48.385 180.335 48.525 ;
        RECT 177.820 48.340 178.110 48.385 ;
        RECT 177.345 48.185 177.665 48.245 ;
        RECT 179.660 48.185 179.950 48.230 ;
        RECT 177.345 48.045 179.950 48.185 ;
        RECT 180.195 48.185 180.335 48.385 ;
        RECT 180.530 48.385 185.830 48.525 ;
        RECT 180.530 48.340 180.820 48.385 ;
        RECT 182.420 48.340 182.710 48.385 ;
        RECT 185.540 48.340 185.830 48.385 ;
        RECT 181.040 48.185 181.330 48.230 ;
        RECT 180.195 48.045 181.330 48.185 ;
        RECT 177.345 47.985 177.665 48.045 ;
        RECT 179.660 48.000 179.950 48.045 ;
        RECT 181.040 48.000 181.330 48.045 ;
        RECT 176.900 47.845 177.190 47.890 ;
        RECT 180.125 47.845 180.415 47.890 ;
        RECT 181.960 47.845 182.250 47.890 ;
        RECT 185.540 47.845 185.830 47.890 ;
        RECT 176.900 47.705 179.875 47.845 ;
        RECT 176.900 47.660 177.190 47.705 ;
        RECT 179.735 47.165 179.875 47.705 ;
        RECT 180.125 47.705 185.830 47.845 ;
        RECT 180.125 47.660 180.415 47.705 ;
        RECT 181.960 47.660 182.250 47.705 ;
        RECT 185.540 47.660 185.830 47.705 ;
        RECT 183.320 47.505 183.970 47.550 ;
        RECT 186.085 47.505 186.405 47.565 ;
        RECT 186.620 47.550 186.910 47.865 ;
        RECT 189.855 47.565 189.995 48.725 ;
        RECT 192.490 48.525 192.780 48.570 ;
        RECT 194.380 48.525 194.670 48.570 ;
        RECT 197.500 48.525 197.790 48.570 ;
        RECT 192.490 48.385 197.790 48.525 ;
        RECT 201.355 48.525 201.495 48.725 ;
        RECT 201.725 48.725 205.265 48.865 ;
        RECT 201.725 48.665 202.045 48.725 ;
        RECT 204.945 48.665 205.265 48.725 ;
        RECT 205.420 48.865 205.710 48.910 ;
        RECT 207.705 48.865 208.025 48.925 ;
        RECT 205.420 48.725 208.025 48.865 ;
        RECT 205.420 48.680 205.710 48.725 ;
        RECT 207.705 48.665 208.025 48.725 ;
        RECT 210.005 48.665 210.325 48.925 ;
        RECT 210.925 48.865 211.245 48.925 ;
        RECT 215.525 48.865 215.845 48.925 ;
        RECT 210.925 48.725 215.845 48.865 ;
        RECT 210.925 48.665 211.245 48.725 ;
        RECT 215.525 48.665 215.845 48.725 ;
        RECT 219.680 48.865 219.970 48.910 ;
        RECT 223.805 48.865 224.125 48.925 ;
        RECT 219.680 48.725 224.125 48.865 ;
        RECT 219.680 48.680 219.970 48.725 ;
        RECT 223.805 48.665 224.125 48.725 ;
        RECT 230.245 48.665 230.565 48.925 ;
        RECT 243.125 48.865 243.445 48.925 ;
        RECT 239.535 48.725 243.445 48.865 ;
        RECT 202.185 48.525 202.505 48.585 ;
        RECT 201.355 48.385 202.505 48.525 ;
        RECT 210.095 48.525 210.235 48.665 ;
        RECT 213.700 48.525 213.990 48.570 ;
        RECT 210.095 48.385 213.990 48.525 ;
        RECT 192.490 48.340 192.780 48.385 ;
        RECT 194.380 48.340 194.670 48.385 ;
        RECT 197.500 48.340 197.790 48.385 ;
        RECT 202.185 48.325 202.505 48.385 ;
        RECT 213.700 48.340 213.990 48.385 ;
        RECT 220.585 48.525 220.905 48.585 ;
        RECT 223.360 48.525 223.650 48.570 ;
        RECT 230.335 48.525 230.475 48.665 ;
        RECT 220.585 48.385 230.475 48.525 ;
        RECT 230.670 48.525 230.960 48.570 ;
        RECT 232.560 48.525 232.850 48.570 ;
        RECT 235.680 48.525 235.970 48.570 ;
        RECT 230.670 48.385 235.970 48.525 ;
        RECT 220.585 48.325 220.905 48.385 ;
        RECT 223.360 48.340 223.650 48.385 ;
        RECT 230.670 48.340 230.960 48.385 ;
        RECT 232.560 48.340 232.850 48.385 ;
        RECT 235.680 48.340 235.970 48.385 ;
        RECT 238.540 48.525 238.830 48.570 ;
        RECT 239.535 48.525 239.675 48.725 ;
        RECT 243.125 48.665 243.445 48.725 ;
        RECT 247.725 48.665 248.045 48.925 ;
        RECT 256.875 48.865 257.165 48.910 ;
        RECT 259.685 48.865 260.005 48.925 ;
        RECT 256.875 48.725 260.005 48.865 ;
        RECT 256.875 48.680 257.165 48.725 ;
        RECT 259.685 48.665 260.005 48.725 ;
        RECT 262.905 48.865 263.225 48.925 ;
        RECT 267.980 48.865 268.270 48.910 ;
        RECT 271.645 48.865 271.965 48.925 ;
        RECT 262.905 48.725 271.965 48.865 ;
        RECT 262.905 48.665 263.225 48.725 ;
        RECT 267.980 48.680 268.270 48.725 ;
        RECT 271.645 48.665 271.965 48.725 ;
        RECT 272.105 48.665 272.425 48.925 ;
        RECT 293.725 48.665 294.045 48.925 ;
        RECT 238.540 48.385 239.675 48.525 ;
        RECT 239.870 48.525 240.160 48.570 ;
        RECT 241.760 48.525 242.050 48.570 ;
        RECT 244.880 48.525 245.170 48.570 ;
        RECT 239.870 48.385 245.170 48.525 ;
        RECT 238.540 48.340 238.830 48.385 ;
        RECT 239.870 48.340 240.160 48.385 ;
        RECT 241.760 48.340 242.050 48.385 ;
        RECT 244.880 48.340 245.170 48.385 ;
        RECT 256.430 48.525 256.720 48.570 ;
        RECT 258.320 48.525 258.610 48.570 ;
        RECT 261.440 48.525 261.730 48.570 ;
        RECT 256.430 48.385 261.730 48.525 ;
        RECT 256.430 48.340 256.720 48.385 ;
        RECT 258.320 48.340 258.610 48.385 ;
        RECT 261.440 48.340 261.730 48.385 ;
        RECT 266.125 48.525 266.445 48.585 ;
        RECT 269.345 48.525 269.665 48.585 ;
        RECT 266.125 48.385 269.665 48.525 ;
        RECT 266.125 48.325 266.445 48.385 ;
        RECT 269.345 48.325 269.665 48.385 ;
        RECT 273.025 48.325 273.345 48.585 ;
        RECT 288.320 48.525 288.610 48.570 ;
        RECT 291.440 48.525 291.730 48.570 ;
        RECT 293.330 48.525 293.620 48.570 ;
        RECT 288.320 48.385 293.620 48.525 ;
        RECT 288.320 48.340 288.610 48.385 ;
        RECT 291.440 48.340 291.730 48.385 ;
        RECT 293.330 48.340 293.620 48.385 ;
        RECT 193.445 48.185 193.765 48.245 ;
        RECT 190.315 48.045 193.765 48.185 ;
        RECT 190.315 47.890 190.455 48.045 ;
        RECT 193.445 47.985 193.765 48.045 ;
        RECT 200.360 48.185 200.650 48.230 ;
        RECT 214.605 48.185 214.925 48.245 ;
        RECT 217.840 48.185 218.130 48.230 ;
        RECT 200.360 48.045 209.775 48.185 ;
        RECT 200.360 48.000 200.650 48.045 ;
        RECT 190.240 47.660 190.530 47.890 ;
        RECT 190.685 47.845 191.005 47.905 ;
        RECT 191.620 47.845 191.910 47.890 ;
        RECT 190.685 47.705 191.910 47.845 ;
        RECT 190.685 47.645 191.005 47.705 ;
        RECT 191.620 47.660 191.910 47.705 ;
        RECT 192.085 47.845 192.375 47.890 ;
        RECT 193.920 47.845 194.210 47.890 ;
        RECT 197.500 47.845 197.790 47.890 ;
        RECT 192.085 47.705 197.790 47.845 ;
        RECT 192.085 47.660 192.375 47.705 ;
        RECT 193.920 47.660 194.210 47.705 ;
        RECT 197.500 47.660 197.790 47.705 ;
        RECT 186.620 47.505 187.210 47.550 ;
        RECT 183.320 47.365 187.210 47.505 ;
        RECT 183.320 47.320 183.970 47.365 ;
        RECT 186.085 47.305 186.405 47.365 ;
        RECT 186.920 47.320 187.210 47.365 ;
        RECT 189.765 47.305 190.085 47.565 ;
        RECT 198.580 47.550 198.870 47.865 ;
        RECT 202.185 47.645 202.505 47.905 ;
        RECT 203.195 47.890 203.335 48.045 ;
        RECT 209.635 47.905 209.775 48.045 ;
        RECT 214.605 48.045 218.130 48.185 ;
        RECT 214.605 47.985 214.925 48.045 ;
        RECT 217.840 48.000 218.130 48.045 ;
        RECT 219.665 48.185 219.985 48.245 ;
        RECT 229.800 48.185 230.090 48.230 ;
        RECT 219.665 48.045 230.090 48.185 ;
        RECT 219.665 47.985 219.985 48.045 ;
        RECT 229.800 48.000 230.090 48.045 ;
        RECT 231.180 48.185 231.470 48.230 ;
        RECT 234.385 48.185 234.705 48.245 ;
        RECT 231.180 48.045 234.705 48.185 ;
        RECT 231.180 48.000 231.470 48.045 ;
        RECT 234.385 47.985 234.705 48.045 ;
        RECT 240.365 47.985 240.685 48.245 ;
        RECT 255.560 48.185 255.850 48.230 ;
        RECT 256.925 48.185 257.245 48.245 ;
        RECT 259.225 48.185 259.545 48.245 ;
        RECT 255.560 48.045 259.545 48.185 ;
        RECT 255.560 48.000 255.850 48.045 ;
        RECT 256.925 47.985 257.245 48.045 ;
        RECT 259.225 47.985 259.545 48.045 ;
        RECT 264.300 48.185 264.590 48.230 ;
        RECT 264.760 48.185 265.050 48.230 ;
        RECT 273.115 48.185 273.255 48.325 ;
        RECT 278.560 48.185 278.850 48.230 ;
        RECT 284.080 48.185 284.370 48.230 ;
        RECT 293.815 48.185 293.955 48.665 ;
        RECT 295.530 48.525 295.820 48.570 ;
        RECT 297.420 48.525 297.710 48.570 ;
        RECT 300.540 48.525 300.830 48.570 ;
        RECT 295.530 48.385 300.830 48.525 ;
        RECT 295.530 48.340 295.820 48.385 ;
        RECT 297.420 48.340 297.710 48.385 ;
        RECT 300.540 48.340 300.830 48.385 ;
        RECT 264.300 48.045 265.050 48.185 ;
        RECT 264.300 48.000 264.590 48.045 ;
        RECT 264.760 48.000 265.050 48.045 ;
        RECT 269.410 48.045 272.885 48.185 ;
        RECT 273.115 48.045 274.175 48.185 ;
        RECT 203.120 47.660 203.410 47.890 ;
        RECT 204.500 47.845 204.790 47.890 ;
        RECT 203.655 47.705 204.790 47.845 ;
        RECT 193.000 47.505 193.290 47.550 ;
        RECT 191.235 47.365 193.290 47.505 ;
        RECT 181.945 47.165 182.265 47.225 ;
        RECT 191.235 47.210 191.375 47.365 ;
        RECT 193.000 47.320 193.290 47.365 ;
        RECT 195.280 47.505 195.930 47.550 ;
        RECT 198.580 47.505 199.170 47.550 ;
        RECT 200.345 47.505 200.665 47.565 ;
        RECT 195.280 47.365 200.665 47.505 ;
        RECT 202.275 47.505 202.415 47.645 ;
        RECT 203.655 47.505 203.795 47.705 ;
        RECT 204.500 47.660 204.790 47.705 ;
        RECT 204.945 47.845 205.265 47.905 ;
        RECT 205.420 47.845 205.710 47.890 ;
        RECT 208.165 47.845 208.485 47.905 ;
        RECT 204.945 47.705 208.485 47.845 ;
        RECT 204.945 47.645 205.265 47.705 ;
        RECT 205.420 47.660 205.710 47.705 ;
        RECT 208.165 47.645 208.485 47.705 ;
        RECT 209.545 47.645 209.865 47.905 ;
        RECT 218.760 47.845 219.050 47.890 ;
        RECT 219.205 47.845 219.525 47.905 ;
        RECT 218.760 47.705 219.525 47.845 ;
        RECT 218.760 47.660 219.050 47.705 ;
        RECT 219.205 47.645 219.525 47.705 ;
        RECT 220.125 47.645 220.445 47.905 ;
        RECT 222.425 47.845 222.745 47.905 ;
        RECT 222.425 47.705 225.415 47.845 ;
        RECT 222.425 47.645 222.745 47.705 ;
        RECT 209.100 47.505 209.390 47.550 ;
        RECT 202.275 47.365 203.795 47.505 ;
        RECT 204.575 47.365 209.390 47.505 ;
        RECT 195.280 47.320 195.930 47.365 ;
        RECT 198.880 47.320 199.170 47.365 ;
        RECT 200.345 47.305 200.665 47.365 ;
        RECT 204.575 47.225 204.715 47.365 ;
        RECT 209.100 47.320 209.390 47.365 ;
        RECT 213.240 47.505 213.530 47.550 ;
        RECT 220.215 47.505 220.355 47.645 ;
        RECT 213.240 47.365 220.355 47.505 ;
        RECT 213.240 47.320 213.530 47.365 ;
        RECT 179.735 47.025 182.265 47.165 ;
        RECT 181.945 46.965 182.265 47.025 ;
        RECT 191.160 46.980 191.450 47.210 ;
        RECT 202.660 47.165 202.950 47.210 ;
        RECT 203.105 47.165 203.425 47.225 ;
        RECT 202.660 47.025 203.425 47.165 ;
        RECT 202.660 46.980 202.950 47.025 ;
        RECT 203.105 46.965 203.425 47.025 ;
        RECT 204.485 46.965 204.805 47.225 ;
        RECT 208.165 47.165 208.485 47.225 ;
        RECT 215.065 47.165 215.385 47.225 ;
        RECT 215.540 47.165 215.830 47.210 ;
        RECT 208.165 47.025 215.830 47.165 ;
        RECT 208.165 46.965 208.485 47.025 ;
        RECT 215.065 46.965 215.385 47.025 ;
        RECT 215.540 46.980 215.830 47.025 ;
        RECT 216.445 46.965 216.765 47.225 ;
        RECT 224.725 46.965 225.045 47.225 ;
        RECT 225.275 47.165 225.415 47.705 ;
        RECT 225.660 47.660 225.950 47.890 ;
        RECT 225.735 47.505 225.875 47.660 ;
        RECT 227.025 47.645 227.345 47.905 ;
        RECT 230.265 47.845 230.555 47.890 ;
        RECT 232.100 47.845 232.390 47.890 ;
        RECT 235.680 47.845 235.970 47.890 ;
        RECT 230.265 47.705 235.970 47.845 ;
        RECT 230.265 47.660 230.555 47.705 ;
        RECT 232.100 47.660 232.390 47.705 ;
        RECT 235.680 47.660 235.970 47.705 ;
        RECT 228.405 47.505 228.725 47.565 ;
        RECT 236.760 47.550 237.050 47.865 ;
        RECT 238.985 47.645 239.305 47.905 ;
        RECT 269.410 47.890 269.550 48.045 ;
        RECT 272.745 47.905 272.885 48.045 ;
        RECT 239.465 47.845 239.755 47.890 ;
        RECT 241.300 47.845 241.590 47.890 ;
        RECT 244.880 47.845 245.170 47.890 ;
        RECT 239.465 47.705 245.170 47.845 ;
        RECT 239.465 47.660 239.755 47.705 ;
        RECT 241.300 47.660 241.590 47.705 ;
        RECT 244.880 47.660 245.170 47.705 ;
        RECT 242.665 47.550 242.985 47.565 ;
        RECT 245.960 47.550 246.250 47.865 ;
        RECT 256.025 47.845 256.315 47.890 ;
        RECT 257.860 47.845 258.150 47.890 ;
        RECT 261.440 47.845 261.730 47.890 ;
        RECT 256.025 47.705 261.730 47.845 ;
        RECT 256.025 47.660 256.315 47.705 ;
        RECT 257.860 47.660 258.150 47.705 ;
        RECT 261.440 47.660 261.730 47.705 ;
        RECT 262.520 47.550 262.810 47.865 ;
        RECT 269.335 47.660 269.625 47.890 ;
        RECT 225.735 47.365 228.725 47.505 ;
        RECT 228.405 47.305 228.725 47.365 ;
        RECT 233.460 47.505 234.110 47.550 ;
        RECT 236.760 47.505 237.350 47.550 ;
        RECT 242.660 47.505 243.310 47.550 ;
        RECT 245.960 47.505 246.550 47.550 ;
        RECT 233.460 47.365 246.550 47.505 ;
        RECT 233.460 47.320 234.110 47.365 ;
        RECT 237.060 47.320 237.350 47.365 ;
        RECT 242.660 47.320 243.310 47.365 ;
        RECT 246.260 47.320 246.550 47.365 ;
        RECT 259.220 47.505 259.870 47.550 ;
        RECT 262.520 47.505 263.110 47.550 ;
        RECT 265.665 47.505 265.985 47.565 ;
        RECT 266.585 47.505 266.905 47.565 ;
        RECT 269.410 47.505 269.550 47.660 ;
        RECT 269.805 47.645 270.125 47.905 ;
        RECT 271.185 47.645 271.505 47.905 ;
        RECT 271.645 47.645 271.965 47.905 ;
        RECT 272.565 47.890 272.885 47.905 ;
        RECT 272.565 47.660 273.100 47.890 ;
        RECT 272.565 47.645 272.885 47.660 ;
        RECT 273.485 47.645 273.805 47.905 ;
        RECT 274.035 47.845 274.175 48.045 ;
        RECT 274.955 48.045 278.850 48.185 ;
        RECT 274.955 47.890 275.095 48.045 ;
        RECT 278.560 48.000 278.850 48.045 ;
        RECT 279.095 48.045 293.955 48.185 ;
        RECT 294.185 48.185 294.505 48.245 ;
        RECT 294.660 48.185 294.950 48.230 ;
        RECT 294.185 48.045 294.950 48.185 ;
        RECT 274.035 47.705 274.635 47.845 ;
        RECT 270.280 47.505 270.570 47.550 ;
        RECT 259.220 47.365 266.905 47.505 ;
        RECT 259.220 47.320 259.870 47.365 ;
        RECT 262.820 47.320 263.110 47.365 ;
        RECT 242.665 47.305 242.985 47.320 ;
        RECT 265.665 47.305 265.985 47.365 ;
        RECT 266.585 47.305 266.905 47.365 ;
        RECT 268.055 47.365 269.550 47.505 ;
        RECT 269.895 47.365 270.570 47.505 ;
        RECT 226.105 47.165 226.425 47.225 ;
        RECT 225.275 47.025 226.425 47.165 ;
        RECT 226.105 46.965 226.425 47.025 ;
        RECT 227.945 47.165 228.265 47.225 ;
        RECT 234.385 47.165 234.705 47.225 ;
        RECT 227.945 47.025 234.705 47.165 ;
        RECT 227.945 46.965 228.265 47.025 ;
        RECT 234.385 46.965 234.705 47.025 ;
        RECT 260.605 47.165 260.925 47.225 ;
        RECT 268.055 47.165 268.195 47.365 ;
        RECT 269.895 47.225 270.035 47.365 ;
        RECT 270.280 47.320 270.570 47.365 ;
        RECT 273.960 47.320 274.250 47.550 ;
        RECT 274.495 47.505 274.635 47.705 ;
        RECT 274.875 47.660 275.165 47.890 ;
        RECT 275.340 47.845 275.630 47.890 ;
        RECT 275.800 47.845 276.090 47.890 ;
        RECT 275.340 47.705 276.090 47.845 ;
        RECT 275.340 47.660 275.630 47.705 ;
        RECT 275.800 47.660 276.090 47.705 ;
        RECT 276.720 47.660 277.010 47.890 ;
        RECT 277.640 47.845 277.930 47.890 ;
        RECT 278.085 47.845 278.405 47.905 ;
        RECT 279.095 47.845 279.235 48.045 ;
        RECT 284.080 48.000 284.370 48.045 ;
        RECT 294.185 47.985 294.505 48.045 ;
        RECT 294.660 48.000 294.950 48.045 ;
        RECT 303.400 48.185 303.690 48.230 ;
        RECT 307.080 48.185 307.370 48.230 ;
        RECT 303.400 48.045 307.370 48.185 ;
        RECT 303.400 48.000 303.690 48.045 ;
        RECT 307.080 48.000 307.370 48.045 ;
        RECT 277.640 47.705 279.235 47.845 ;
        RECT 280.845 47.845 281.165 47.905 ;
        RECT 281.320 47.845 281.610 47.890 ;
        RECT 280.845 47.705 281.610 47.845 ;
        RECT 277.640 47.660 277.930 47.705 ;
        RECT 276.795 47.505 276.935 47.660 ;
        RECT 278.085 47.645 278.405 47.705 ;
        RECT 280.845 47.645 281.165 47.705 ;
        RECT 281.320 47.660 281.610 47.705 ;
        RECT 281.765 47.845 282.085 47.905 ;
        RECT 283.160 47.845 283.450 47.890 ;
        RECT 281.765 47.705 283.450 47.845 ;
        RECT 281.765 47.645 282.085 47.705 ;
        RECT 283.160 47.660 283.450 47.705 ;
        RECT 279.465 47.505 279.785 47.565 ;
        RECT 287.240 47.550 287.530 47.865 ;
        RECT 288.320 47.845 288.610 47.890 ;
        RECT 291.900 47.845 292.190 47.890 ;
        RECT 293.735 47.845 294.025 47.890 ;
        RECT 288.320 47.705 294.025 47.845 ;
        RECT 288.320 47.660 288.610 47.705 ;
        RECT 291.900 47.660 292.190 47.705 ;
        RECT 293.735 47.660 294.025 47.705 ;
        RECT 295.125 47.845 295.415 47.890 ;
        RECT 296.960 47.845 297.250 47.890 ;
        RECT 300.540 47.845 300.830 47.890 ;
        RECT 295.125 47.705 300.830 47.845 ;
        RECT 295.125 47.660 295.415 47.705 ;
        RECT 296.960 47.660 297.250 47.705 ;
        RECT 300.540 47.660 300.830 47.705 ;
        RECT 290.505 47.550 290.825 47.565 ;
        RECT 274.495 47.365 276.935 47.505 ;
        RECT 278.175 47.365 279.785 47.505 ;
        RECT 260.605 47.025 268.195 47.165 ;
        RECT 260.605 46.965 260.925 47.025 ;
        RECT 268.425 46.965 268.745 47.225 ;
        RECT 269.805 46.965 270.125 47.225 ;
        RECT 274.035 47.165 274.175 47.320 ;
        RECT 274.865 47.165 275.185 47.225 ;
        RECT 278.175 47.165 278.315 47.365 ;
        RECT 279.465 47.305 279.785 47.365 ;
        RECT 286.940 47.505 287.530 47.550 ;
        RECT 290.180 47.505 290.830 47.550 ;
        RECT 292.820 47.505 293.110 47.550 ;
        RECT 294.645 47.505 294.965 47.565 ;
        RECT 286.940 47.365 292.575 47.505 ;
        RECT 286.940 47.320 287.230 47.365 ;
        RECT 290.180 47.320 290.830 47.365 ;
        RECT 290.505 47.305 290.825 47.320 ;
        RECT 274.035 47.025 278.315 47.165 ;
        RECT 278.545 47.165 278.865 47.225 ;
        RECT 282.240 47.165 282.530 47.210 ;
        RECT 278.545 47.025 282.530 47.165 ;
        RECT 274.865 46.965 275.185 47.025 ;
        RECT 278.545 46.965 278.865 47.025 ;
        RECT 282.240 46.980 282.530 47.025 ;
        RECT 285.445 47.165 285.765 47.225 ;
        RECT 291.885 47.165 292.205 47.225 ;
        RECT 285.445 47.025 292.205 47.165 ;
        RECT 292.435 47.165 292.575 47.365 ;
        RECT 292.820 47.365 294.965 47.505 ;
        RECT 292.820 47.320 293.110 47.365 ;
        RECT 294.645 47.305 294.965 47.365 ;
        RECT 295.565 47.305 295.885 47.565 ;
        RECT 296.025 47.305 296.345 47.565 ;
        RECT 301.620 47.550 301.910 47.865 ;
        RECT 298.320 47.505 298.970 47.550 ;
        RECT 301.620 47.505 302.210 47.550 ;
        RECT 305.225 47.505 305.545 47.565 ;
        RECT 298.320 47.365 305.545 47.505 ;
        RECT 298.320 47.320 298.970 47.365 ;
        RECT 301.920 47.320 302.210 47.365 ;
        RECT 305.225 47.305 305.545 47.365 ;
        RECT 295.655 47.165 295.795 47.305 ;
        RECT 292.435 47.025 295.795 47.165 ;
        RECT 297.865 47.165 298.185 47.225 ;
        RECT 304.320 47.165 304.610 47.210 ;
        RECT 297.865 47.025 304.610 47.165 ;
        RECT 285.445 46.965 285.765 47.025 ;
        RECT 291.885 46.965 292.205 47.025 ;
        RECT 297.865 46.965 298.185 47.025 ;
        RECT 304.320 46.980 304.610 47.025 ;
        RECT 162.095 46.345 311.935 46.825 ;
        RECT 193.445 45.945 193.765 46.205 ;
        RECT 195.300 46.145 195.590 46.190 ;
        RECT 203.105 46.145 203.425 46.205 ;
        RECT 195.300 46.005 203.425 46.145 ;
        RECT 195.300 45.960 195.590 46.005 ;
        RECT 203.105 45.945 203.425 46.005 ;
        RECT 215.985 46.145 216.305 46.205 ;
        RECT 217.380 46.145 217.670 46.190 ;
        RECT 215.985 46.005 217.670 46.145 ;
        RECT 215.985 45.945 216.305 46.005 ;
        RECT 217.380 45.960 217.670 46.005 ;
        RECT 242.665 45.945 242.985 46.205 ;
        RECT 249.105 46.145 249.425 46.205 ;
        RECT 246.895 46.005 249.425 46.145 ;
        RECT 181.020 45.805 181.670 45.850 ;
        RECT 184.620 45.805 184.910 45.850 ;
        RECT 181.020 45.665 184.910 45.805 ;
        RECT 181.020 45.620 181.670 45.665 ;
        RECT 184.320 45.620 184.910 45.665 ;
        RECT 187.480 45.805 187.770 45.850 ;
        RECT 190.240 45.805 190.530 45.850 ;
        RECT 192.985 45.805 193.305 45.865 ;
        RECT 187.480 45.665 193.305 45.805 ;
        RECT 187.480 45.620 187.770 45.665 ;
        RECT 190.240 45.620 190.530 45.665 ;
        RECT 177.825 45.465 178.115 45.510 ;
        RECT 179.660 45.465 179.950 45.510 ;
        RECT 183.240 45.465 183.530 45.510 ;
        RECT 177.825 45.325 183.530 45.465 ;
        RECT 177.825 45.280 178.115 45.325 ;
        RECT 179.660 45.280 179.950 45.325 ;
        RECT 183.240 45.280 183.530 45.325 ;
        RECT 184.320 45.465 184.610 45.620 ;
        RECT 192.985 45.605 193.305 45.665 ;
        RECT 203.560 45.805 204.210 45.850 ;
        RECT 207.160 45.805 207.450 45.850 ;
        RECT 203.560 45.665 207.450 45.805 ;
        RECT 203.560 45.620 204.210 45.665 ;
        RECT 206.860 45.620 207.450 45.665 ;
        RECT 215.540 45.805 215.830 45.850 ;
        RECT 216.445 45.805 216.765 45.865 ;
        RECT 215.540 45.665 216.765 45.805 ;
        RECT 215.540 45.620 215.830 45.665 ;
        RECT 186.085 45.465 186.405 45.525 ;
        RECT 195.285 45.465 195.605 45.525 ;
        RECT 184.320 45.325 195.605 45.465 ;
        RECT 184.320 45.305 184.610 45.325 ;
        RECT 176.425 44.925 176.745 45.185 ;
        RECT 177.360 44.940 177.650 45.170 ;
        RECT 177.435 44.505 177.575 44.940 ;
        RECT 178.725 44.925 179.045 45.185 ;
        RECT 179.185 45.125 179.505 45.185 ;
        RECT 184.335 45.125 184.475 45.305 ;
        RECT 186.085 45.265 186.405 45.325 ;
        RECT 195.285 45.265 195.605 45.325 ;
        RECT 195.760 45.465 196.050 45.510 ;
        RECT 200.365 45.465 200.655 45.510 ;
        RECT 202.200 45.465 202.490 45.510 ;
        RECT 205.780 45.465 206.070 45.510 ;
        RECT 195.760 45.325 198.275 45.465 ;
        RECT 195.760 45.280 196.050 45.325 ;
        RECT 198.135 45.185 198.275 45.325 ;
        RECT 200.365 45.325 206.070 45.465 ;
        RECT 200.365 45.280 200.655 45.325 ;
        RECT 202.200 45.280 202.490 45.325 ;
        RECT 205.780 45.280 206.070 45.325 ;
        RECT 206.860 45.465 207.150 45.620 ;
        RECT 216.445 45.605 216.765 45.665 ;
        RECT 223.340 45.805 223.990 45.850 ;
        RECT 226.940 45.805 227.230 45.850 ;
        RECT 223.340 45.665 227.230 45.805 ;
        RECT 242.755 45.805 242.895 45.945 ;
        RECT 246.895 45.805 247.035 46.005 ;
        RECT 249.105 45.945 249.425 46.005 ;
        RECT 257.845 46.145 258.165 46.205 ;
        RECT 269.805 46.145 270.125 46.205 ;
        RECT 274.865 46.145 275.185 46.205 ;
        RECT 257.845 46.005 275.185 46.145 ;
        RECT 257.845 45.945 258.165 46.005 ;
        RECT 269.805 45.945 270.125 46.005 ;
        RECT 274.865 45.945 275.185 46.005 ;
        RECT 277.625 46.145 277.945 46.205 ;
        RECT 281.780 46.145 282.070 46.190 ;
        RECT 290.505 46.145 290.825 46.205 ;
        RECT 295.105 46.145 295.425 46.205 ;
        RECT 277.625 46.005 282.070 46.145 ;
        RECT 277.625 45.945 277.945 46.005 ;
        RECT 281.780 45.960 282.070 46.005 ;
        RECT 283.465 46.005 290.825 46.145 ;
        RECT 247.260 45.805 247.910 45.850 ;
        RECT 250.860 45.805 251.150 45.850 ;
        RECT 242.755 45.665 251.150 45.805 ;
        RECT 223.340 45.620 223.990 45.665 ;
        RECT 226.640 45.620 227.230 45.665 ;
        RECT 247.260 45.620 247.910 45.665 ;
        RECT 250.560 45.620 251.150 45.665 ;
        RECT 264.760 45.805 265.050 45.850 ;
        RECT 268.885 45.805 269.205 45.865 ;
        RECT 264.760 45.665 269.205 45.805 ;
        RECT 264.760 45.620 265.050 45.665 ;
        RECT 226.640 45.525 226.930 45.620 ;
        RECT 209.085 45.465 209.405 45.525 ;
        RECT 216.920 45.465 217.210 45.510 ;
        RECT 206.860 45.325 209.405 45.465 ;
        RECT 206.860 45.305 207.150 45.325 ;
        RECT 209.085 45.265 209.405 45.325 ;
        RECT 215.615 45.325 217.210 45.465 ;
        RECT 215.615 45.185 215.755 45.325 ;
        RECT 216.920 45.280 217.210 45.325 ;
        RECT 220.145 45.465 220.435 45.510 ;
        RECT 221.980 45.465 222.270 45.510 ;
        RECT 225.560 45.465 225.850 45.510 ;
        RECT 220.145 45.325 225.850 45.465 ;
        RECT 220.145 45.280 220.435 45.325 ;
        RECT 221.980 45.280 222.270 45.325 ;
        RECT 225.560 45.280 225.850 45.325 ;
        RECT 226.565 45.305 226.930 45.525 ;
        RECT 230.705 45.465 231.025 45.525 ;
        RECT 233.005 45.465 233.325 45.525 ;
        RECT 230.705 45.325 233.325 45.465 ;
        RECT 226.565 45.265 226.885 45.305 ;
        RECT 230.705 45.265 231.025 45.325 ;
        RECT 233.005 45.265 233.325 45.325 ;
        RECT 244.065 45.465 244.355 45.510 ;
        RECT 245.900 45.465 246.190 45.510 ;
        RECT 249.480 45.465 249.770 45.510 ;
        RECT 244.065 45.325 249.770 45.465 ;
        RECT 244.065 45.280 244.355 45.325 ;
        RECT 245.900 45.280 246.190 45.325 ;
        RECT 249.480 45.280 249.770 45.325 ;
        RECT 250.560 45.305 250.850 45.620 ;
        RECT 268.885 45.605 269.205 45.665 ;
        RECT 271.200 45.805 271.490 45.850 ;
        RECT 271.645 45.805 271.965 45.865 ;
        RECT 271.200 45.665 271.965 45.805 ;
        RECT 271.200 45.620 271.490 45.665 ;
        RECT 271.645 45.605 271.965 45.665 ;
        RECT 272.105 45.805 272.425 45.865 ;
        RECT 283.465 45.850 283.605 46.005 ;
        RECT 273.960 45.805 274.250 45.850 ;
        RECT 272.105 45.665 274.250 45.805 ;
        RECT 272.105 45.605 272.425 45.665 ;
        RECT 273.960 45.620 274.250 45.665 ;
        RECT 276.240 45.805 276.890 45.850 ;
        RECT 279.840 45.805 280.130 45.850 ;
        RECT 276.240 45.665 280.130 45.805 ;
        RECT 276.240 45.620 276.890 45.665 ;
        RECT 279.540 45.620 280.130 45.665 ;
        RECT 283.260 45.805 283.605 45.850 ;
        RECT 286.500 45.805 287.150 45.850 ;
        RECT 287.745 45.805 288.065 45.865 ;
        RECT 288.295 45.805 288.435 46.005 ;
        RECT 290.505 45.945 290.825 46.005 ;
        RECT 292.895 46.005 295.425 46.145 ;
        RECT 283.260 45.665 288.435 45.805 ;
        RECT 288.665 45.805 288.985 45.865 ;
        RECT 292.895 45.850 293.035 46.005 ;
        RECT 295.105 45.945 295.425 46.005 ;
        RECT 296.025 46.145 296.345 46.205 ;
        RECT 298.800 46.145 299.090 46.190 ;
        RECT 296.025 46.005 299.090 46.145 ;
        RECT 296.025 45.945 296.345 46.005 ;
        RECT 298.800 45.960 299.090 46.005 ;
        RECT 288.665 45.665 290.735 45.805 ;
        RECT 283.260 45.620 283.850 45.665 ;
        RECT 286.500 45.620 287.150 45.665 ;
        RECT 253.260 45.465 253.550 45.510 ;
        RECT 251.495 45.325 253.550 45.465 ;
        RECT 179.185 44.985 184.475 45.125 ;
        RECT 179.185 44.925 179.505 44.985 ;
        RECT 190.685 44.925 191.005 45.185 ;
        RECT 191.620 45.125 191.910 45.170 ;
        RECT 196.680 45.125 196.970 45.170 ;
        RECT 191.620 44.985 197.355 45.125 ;
        RECT 191.620 44.940 191.910 44.985 ;
        RECT 196.680 44.940 196.970 44.985 ;
        RECT 197.215 44.845 197.355 44.985 ;
        RECT 198.045 44.925 198.365 45.185 ;
        RECT 199.900 44.940 200.190 45.170 ;
        RECT 178.230 44.785 178.520 44.830 ;
        RECT 180.120 44.785 180.410 44.830 ;
        RECT 183.240 44.785 183.530 44.830 ;
        RECT 178.230 44.645 183.530 44.785 ;
        RECT 178.230 44.600 178.520 44.645 ;
        RECT 180.120 44.600 180.410 44.645 ;
        RECT 183.240 44.600 183.530 44.645 ;
        RECT 183.875 44.645 190.455 44.785 ;
        RECT 173.665 44.245 173.985 44.505 ;
        RECT 177.345 44.445 177.665 44.505 ;
        RECT 183.875 44.445 184.015 44.645 ;
        RECT 190.315 44.505 190.455 44.645 ;
        RECT 197.125 44.585 197.445 44.845 ;
        RECT 199.975 44.785 200.115 44.940 ;
        RECT 201.265 44.925 201.585 45.185 ;
        RECT 207.705 45.125 208.025 45.185 ;
        RECT 208.625 45.125 208.945 45.185 ;
        RECT 210.020 45.125 210.310 45.170 ;
        RECT 207.705 44.985 210.310 45.125 ;
        RECT 207.705 44.925 208.025 44.985 ;
        RECT 208.625 44.925 208.945 44.985 ;
        RECT 210.020 44.940 210.310 44.985 ;
        RECT 215.525 44.925 215.845 45.185 ;
        RECT 216.445 45.125 216.765 45.185 ;
        RECT 219.665 45.125 219.985 45.185 ;
        RECT 216.445 44.985 219.985 45.125 ;
        RECT 216.445 44.925 216.765 44.985 ;
        RECT 219.665 44.925 219.985 44.985 ;
        RECT 221.060 45.125 221.350 45.170 ;
        RECT 224.725 45.125 225.045 45.185 ;
        RECT 221.060 44.985 225.045 45.125 ;
        RECT 221.060 44.940 221.350 44.985 ;
        RECT 224.725 44.925 225.045 44.985 ;
        RECT 226.105 45.125 226.425 45.185 ;
        RECT 229.800 45.125 230.090 45.170 ;
        RECT 226.105 44.985 230.090 45.125 ;
        RECT 226.105 44.925 226.425 44.985 ;
        RECT 229.800 44.940 230.090 44.985 ;
        RECT 231.625 45.125 231.945 45.185 ;
        RECT 232.100 45.125 232.390 45.170 ;
        RECT 231.625 44.985 232.390 45.125 ;
        RECT 231.625 44.925 231.945 44.985 ;
        RECT 232.100 44.940 232.390 44.985 ;
        RECT 238.985 45.125 239.305 45.185 ;
        RECT 241.745 45.125 242.065 45.185 ;
        RECT 243.600 45.125 243.890 45.170 ;
        RECT 238.985 44.985 243.890 45.125 ;
        RECT 238.985 44.925 239.305 44.985 ;
        RECT 241.745 44.925 242.065 44.985 ;
        RECT 243.600 44.940 243.890 44.985 ;
        RECT 244.965 44.925 245.285 45.185 ;
        RECT 247.265 45.125 247.585 45.185 ;
        RECT 251.495 45.125 251.635 45.325 ;
        RECT 253.260 45.280 253.550 45.325 ;
        RECT 253.705 45.465 254.025 45.525 ;
        RECT 257.860 45.465 258.150 45.510 ;
        RECT 253.705 45.325 258.150 45.465 ;
        RECT 253.705 45.265 254.025 45.325 ;
        RECT 257.860 45.280 258.150 45.325 ;
        RECT 258.855 45.325 268.195 45.465 ;
        RECT 247.265 44.985 251.635 45.125 ;
        RECT 252.340 45.125 252.630 45.170 ;
        RECT 256.020 45.125 256.310 45.170 ;
        RECT 252.340 44.985 256.310 45.125 ;
        RECT 247.265 44.925 247.585 44.985 ;
        RECT 252.340 44.940 252.630 44.985 ;
        RECT 256.020 44.940 256.310 44.985 ;
        RECT 258.305 45.125 258.625 45.185 ;
        RECT 258.855 45.170 258.995 45.325 ;
        RECT 258.780 45.125 259.070 45.170 ;
        RECT 258.305 44.985 259.070 45.125 ;
        RECT 258.305 44.925 258.625 44.985 ;
        RECT 258.780 44.940 259.070 44.985 ;
        RECT 261.065 44.925 261.385 45.185 ;
        RECT 268.055 45.125 268.195 45.325 ;
        RECT 268.425 45.265 268.745 45.525 ;
        RECT 270.265 45.265 270.585 45.525 ;
        RECT 273.045 45.465 273.335 45.510 ;
        RECT 274.880 45.465 275.170 45.510 ;
        RECT 278.460 45.465 278.750 45.510 ;
        RECT 279.540 45.465 279.830 45.620 ;
        RECT 283.465 45.465 283.850 45.620 ;
        RECT 287.745 45.605 288.065 45.665 ;
        RECT 288.665 45.605 288.985 45.665 ;
        RECT 290.595 45.510 290.735 45.665 ;
        RECT 292.820 45.620 293.110 45.850 ;
        RECT 293.280 45.805 293.570 45.850 ;
        RECT 297.865 45.805 298.185 45.865 ;
        RECT 305.225 45.850 305.545 45.865 ;
        RECT 293.280 45.665 298.185 45.805 ;
        RECT 293.280 45.620 293.570 45.665 ;
        RECT 297.865 45.605 298.185 45.665 ;
        RECT 301.955 45.805 302.245 45.850 ;
        RECT 305.215 45.805 305.545 45.850 ;
        RECT 301.955 45.665 305.545 45.805 ;
        RECT 301.955 45.620 302.245 45.665 ;
        RECT 305.215 45.620 305.545 45.665 ;
        RECT 305.225 45.605 305.545 45.620 ;
        RECT 306.135 45.805 306.425 45.850 ;
        RECT 307.995 45.805 308.285 45.850 ;
        RECT 306.135 45.665 308.285 45.805 ;
        RECT 306.135 45.620 306.425 45.665 ;
        RECT 307.995 45.620 308.285 45.665 ;
        RECT 273.045 45.325 278.750 45.465 ;
        RECT 273.045 45.280 273.335 45.325 ;
        RECT 274.880 45.280 275.170 45.325 ;
        RECT 278.460 45.280 278.750 45.325 ;
        RECT 279.095 45.325 283.850 45.465 ;
        RECT 269.345 45.125 269.665 45.185 ;
        RECT 268.055 44.985 269.665 45.125 ;
        RECT 269.345 44.925 269.665 44.985 ;
        RECT 272.580 44.940 272.870 45.170 ;
        RECT 198.135 44.645 200.115 44.785 ;
        RECT 200.770 44.785 201.060 44.830 ;
        RECT 202.660 44.785 202.950 44.830 ;
        RECT 205.780 44.785 206.070 44.830 ;
        RECT 200.770 44.645 206.070 44.785 ;
        RECT 177.345 44.305 184.015 44.445 ;
        RECT 184.245 44.445 184.565 44.505 ;
        RECT 188.400 44.445 188.690 44.490 ;
        RECT 184.245 44.305 188.690 44.445 ;
        RECT 177.345 44.245 177.665 44.305 ;
        RECT 184.245 44.245 184.565 44.305 ;
        RECT 188.400 44.260 188.690 44.305 ;
        RECT 190.225 44.445 190.545 44.505 ;
        RECT 198.135 44.445 198.275 44.645 ;
        RECT 200.770 44.600 201.060 44.645 ;
        RECT 202.660 44.600 202.950 44.645 ;
        RECT 205.780 44.600 206.070 44.645 ;
        RECT 220.550 44.785 220.840 44.830 ;
        RECT 222.440 44.785 222.730 44.830 ;
        RECT 225.560 44.785 225.850 44.830 ;
        RECT 220.550 44.645 225.850 44.785 ;
        RECT 220.550 44.600 220.840 44.645 ;
        RECT 222.440 44.600 222.730 44.645 ;
        RECT 225.560 44.600 225.850 44.645 ;
        RECT 190.225 44.305 198.275 44.445 ;
        RECT 216.000 44.445 216.290 44.490 ;
        RECT 216.905 44.445 217.225 44.505 ;
        RECT 216.000 44.305 217.225 44.445 ;
        RECT 190.225 44.245 190.545 44.305 ;
        RECT 216.000 44.260 216.290 44.305 ;
        RECT 216.905 44.245 217.225 44.305 ;
        RECT 224.265 44.445 224.585 44.505 ;
        RECT 231.715 44.445 231.855 44.925 ;
        RECT 244.470 44.785 244.760 44.830 ;
        RECT 246.360 44.785 246.650 44.830 ;
        RECT 249.480 44.785 249.770 44.830 ;
        RECT 244.470 44.645 249.770 44.785 ;
        RECT 261.155 44.785 261.295 44.925 ;
        RECT 265.205 44.785 265.525 44.845 ;
        RECT 272.655 44.785 272.795 44.940 ;
        RECT 261.155 44.645 272.795 44.785 ;
        RECT 273.450 44.785 273.740 44.830 ;
        RECT 275.340 44.785 275.630 44.830 ;
        RECT 278.460 44.785 278.750 44.830 ;
        RECT 273.450 44.645 278.750 44.785 ;
        RECT 244.470 44.600 244.760 44.645 ;
        RECT 246.360 44.600 246.650 44.645 ;
        RECT 249.480 44.600 249.770 44.645 ;
        RECT 265.205 44.585 265.525 44.645 ;
        RECT 273.450 44.600 273.740 44.645 ;
        RECT 275.340 44.600 275.630 44.645 ;
        RECT 278.460 44.600 278.750 44.645 ;
        RECT 224.265 44.305 231.855 44.445 ;
        RECT 224.265 44.245 224.585 44.305 ;
        RECT 256.925 44.245 257.245 44.505 ;
        RECT 265.665 44.245 265.985 44.505 ;
        RECT 272.105 44.445 272.425 44.505 ;
        RECT 279.095 44.445 279.235 45.325 ;
        RECT 279.540 45.305 279.830 45.325 ;
        RECT 283.560 45.305 283.850 45.325 ;
        RECT 284.640 45.465 284.930 45.510 ;
        RECT 288.220 45.465 288.510 45.510 ;
        RECT 290.055 45.465 290.345 45.510 ;
        RECT 284.640 45.325 290.345 45.465 ;
        RECT 284.640 45.280 284.930 45.325 ;
        RECT 288.220 45.280 288.510 45.325 ;
        RECT 290.055 45.280 290.345 45.325 ;
        RECT 290.520 45.280 290.810 45.510 ;
        RECT 290.965 45.465 291.285 45.525 ;
        RECT 291.440 45.465 291.730 45.510 ;
        RECT 290.965 45.325 291.730 45.465 ;
        RECT 290.965 45.265 291.285 45.325 ;
        RECT 291.440 45.280 291.730 45.325 ;
        RECT 291.885 45.265 292.205 45.525 ;
        RECT 293.725 45.510 294.045 45.525 ;
        RECT 293.725 45.280 294.055 45.510 ;
        RECT 303.815 45.465 304.105 45.510 ;
        RECT 306.135 45.465 306.350 45.620 ;
        RECT 303.815 45.325 306.350 45.465 ;
        RECT 303.815 45.280 304.105 45.325 ;
        RECT 293.725 45.265 294.045 45.280 ;
        RECT 307.065 45.265 307.385 45.525 ;
        RECT 289.125 44.925 289.445 45.185 ;
        RECT 295.580 44.940 295.870 45.170 ;
        RECT 299.950 45.125 300.240 45.170 ;
        RECT 299.950 44.985 300.855 45.125 ;
        RECT 299.950 44.940 300.240 44.985 ;
        RECT 284.065 44.785 284.385 44.845 ;
        RECT 281.395 44.645 284.385 44.785 ;
        RECT 281.395 44.490 281.535 44.645 ;
        RECT 284.065 44.585 284.385 44.645 ;
        RECT 284.640 44.785 284.930 44.830 ;
        RECT 287.760 44.785 288.050 44.830 ;
        RECT 289.650 44.785 289.940 44.830 ;
        RECT 284.640 44.645 289.940 44.785 ;
        RECT 284.640 44.600 284.930 44.645 ;
        RECT 287.760 44.600 288.050 44.645 ;
        RECT 289.650 44.600 289.940 44.645 ;
        RECT 294.660 44.785 294.950 44.830 ;
        RECT 295.655 44.785 295.795 44.940 ;
        RECT 294.660 44.645 295.795 44.785 ;
        RECT 294.660 44.600 294.950 44.645 ;
        RECT 300.715 44.505 300.855 44.985 ;
        RECT 308.905 44.925 309.225 45.185 ;
        RECT 303.815 44.785 304.105 44.830 ;
        RECT 306.595 44.785 306.885 44.830 ;
        RECT 308.455 44.785 308.745 44.830 ;
        RECT 303.815 44.645 308.745 44.785 ;
        RECT 303.815 44.600 304.105 44.645 ;
        RECT 306.595 44.600 306.885 44.645 ;
        RECT 308.455 44.600 308.745 44.645 ;
        RECT 272.105 44.305 279.235 44.445 ;
        RECT 272.105 44.245 272.425 44.305 ;
        RECT 281.320 44.260 281.610 44.490 ;
        RECT 300.625 44.245 300.945 44.505 ;
        RECT 162.095 43.625 311.135 44.105 ;
        RECT 173.665 43.425 173.985 43.485 ;
        RECT 173.065 43.285 173.985 43.425 ;
        RECT 173.065 42.745 173.205 43.285 ;
        RECT 173.665 43.225 173.985 43.285 ;
        RECT 175.520 43.425 175.810 43.470 ;
        RECT 176.425 43.425 176.745 43.485 ;
        RECT 175.520 43.285 176.745 43.425 ;
        RECT 175.520 43.240 175.810 43.285 ;
        RECT 176.425 43.225 176.745 43.285 ;
        RECT 178.725 43.425 179.045 43.485 ;
        RECT 180.120 43.425 180.410 43.470 ;
        RECT 178.725 43.285 180.410 43.425 ;
        RECT 178.725 43.225 179.045 43.285 ;
        RECT 180.120 43.240 180.410 43.285 ;
        RECT 181.945 43.225 182.265 43.485 ;
        RECT 189.320 43.425 189.610 43.470 ;
        RECT 190.685 43.425 191.005 43.485 ;
        RECT 189.320 43.285 191.005 43.425 ;
        RECT 189.320 43.240 189.610 43.285 ;
        RECT 190.685 43.225 191.005 43.285 ;
        RECT 197.125 43.425 197.445 43.485 ;
        RECT 201.725 43.425 202.045 43.485 ;
        RECT 202.595 43.425 202.885 43.470 ;
        RECT 213.685 43.425 214.005 43.485 ;
        RECT 216.460 43.425 216.750 43.470 ;
        RECT 225.185 43.425 225.505 43.485 ;
        RECT 197.125 43.285 225.505 43.425 ;
        RECT 197.125 43.225 197.445 43.285 ;
        RECT 201.725 43.225 202.045 43.285 ;
        RECT 202.595 43.240 202.885 43.285 ;
        RECT 213.685 43.225 214.005 43.285 ;
        RECT 216.460 43.240 216.750 43.285 ;
        RECT 225.185 43.225 225.505 43.285 ;
        RECT 226.120 43.425 226.410 43.470 ;
        RECT 230.705 43.425 231.025 43.485 ;
        RECT 226.120 43.285 231.025 43.425 ;
        RECT 226.120 43.240 226.410 43.285 ;
        RECT 230.705 43.225 231.025 43.285 ;
        RECT 232.545 43.425 232.865 43.485 ;
        RECT 243.600 43.425 243.890 43.470 ;
        RECT 232.545 43.285 243.890 43.425 ;
        RECT 232.545 43.225 232.865 43.285 ;
        RECT 243.600 43.240 243.890 43.285 ;
        RECT 270.280 43.425 270.570 43.470 ;
        RECT 271.185 43.425 271.505 43.485 ;
        RECT 270.280 43.285 271.505 43.425 ;
        RECT 270.280 43.240 270.570 43.285 ;
        RECT 271.185 43.225 271.505 43.285 ;
        RECT 276.335 43.285 281.535 43.425 ;
        RECT 174.600 43.085 174.890 43.130 ;
        RECT 191.110 43.085 191.400 43.130 ;
        RECT 193.000 43.085 193.290 43.130 ;
        RECT 196.120 43.085 196.410 43.130 ;
        RECT 174.600 42.945 184.475 43.085 ;
        RECT 174.600 42.900 174.890 42.945 ;
        RECT 170.995 42.605 173.205 42.745 ;
        RECT 176.885 42.745 177.205 42.805 ;
        RECT 178.280 42.745 178.570 42.790 ;
        RECT 176.885 42.605 178.570 42.745 ;
        RECT 170.995 42.450 171.135 42.605 ;
        RECT 176.885 42.545 177.205 42.605 ;
        RECT 178.280 42.560 178.570 42.605 ;
        RECT 178.815 42.465 178.955 42.945 ;
        RECT 170.920 42.220 171.210 42.450 ;
        RECT 171.840 42.405 172.130 42.450 ;
        RECT 173.665 42.405 173.985 42.465 ;
        RECT 171.840 42.265 173.985 42.405 ;
        RECT 171.840 42.220 172.130 42.265 ;
        RECT 173.665 42.205 173.985 42.265 ;
        RECT 178.725 42.205 179.045 42.465 ;
        RECT 181.040 42.385 181.330 42.450 ;
        RECT 183.785 42.405 184.105 42.465 ;
        RECT 184.335 42.450 184.475 42.945 ;
        RECT 191.110 42.945 196.410 43.085 ;
        RECT 191.110 42.900 191.400 42.945 ;
        RECT 193.000 42.900 193.290 42.945 ;
        RECT 196.120 42.900 196.410 42.945 ;
        RECT 185.180 42.745 185.470 42.790 ;
        RECT 197.215 42.745 197.355 43.225 ;
        RECT 202.150 43.085 202.440 43.130 ;
        RECT 204.040 43.085 204.330 43.130 ;
        RECT 207.160 43.085 207.450 43.130 ;
        RECT 202.150 42.945 207.450 43.085 ;
        RECT 202.150 42.900 202.440 42.945 ;
        RECT 204.040 42.900 204.330 42.945 ;
        RECT 207.160 42.900 207.450 42.945 ;
        RECT 213.225 42.885 213.545 43.145 ;
        RECT 218.250 43.085 218.540 43.130 ;
        RECT 220.140 43.085 220.430 43.130 ;
        RECT 223.260 43.085 223.550 43.130 ;
        RECT 218.250 42.945 223.550 43.085 ;
        RECT 218.250 42.900 218.540 42.945 ;
        RECT 220.140 42.900 220.430 42.945 ;
        RECT 223.260 42.900 223.550 42.945 ;
        RECT 231.280 43.085 231.570 43.130 ;
        RECT 234.400 43.085 234.690 43.130 ;
        RECT 236.290 43.085 236.580 43.130 ;
        RECT 258.305 43.085 258.625 43.145 ;
        RECT 231.280 42.945 236.580 43.085 ;
        RECT 231.280 42.900 231.570 42.945 ;
        RECT 234.400 42.900 234.690 42.945 ;
        RECT 236.290 42.900 236.580 42.945 ;
        RECT 254.255 42.945 258.625 43.085 ;
        RECT 185.180 42.605 197.355 42.745 ;
        RECT 201.280 42.745 201.570 42.790 ;
        RECT 204.485 42.745 204.805 42.805 ;
        RECT 201.280 42.605 204.805 42.745 ;
        RECT 185.180 42.560 185.470 42.605 ;
        RECT 201.280 42.560 201.570 42.605 ;
        RECT 204.485 42.545 204.805 42.605 ;
        RECT 211.400 42.745 211.690 42.790 ;
        RECT 211.860 42.745 212.150 42.790 ;
        RECT 214.145 42.745 214.465 42.805 ;
        RECT 226.565 42.745 226.885 42.805 ;
        RECT 233.465 42.745 233.785 42.805 ;
        RECT 211.400 42.605 214.465 42.745 ;
        RECT 211.400 42.560 211.690 42.605 ;
        RECT 211.860 42.560 212.150 42.605 ;
        RECT 214.145 42.545 214.465 42.605 ;
        RECT 224.355 42.605 233.785 42.745 ;
        RECT 181.575 42.385 184.105 42.405 ;
        RECT 181.040 42.265 184.105 42.385 ;
        RECT 181.040 42.245 181.715 42.265 ;
        RECT 181.040 42.220 181.330 42.245 ;
        RECT 183.785 42.205 184.105 42.265 ;
        RECT 184.260 42.220 184.550 42.450 ;
        RECT 186.100 42.220 186.390 42.450 ;
        RECT 177.360 42.065 177.650 42.110 ;
        RECT 179.645 42.065 179.965 42.125 ;
        RECT 186.175 42.065 186.315 42.220 ;
        RECT 190.225 42.205 190.545 42.465 ;
        RECT 190.705 42.405 190.995 42.450 ;
        RECT 192.540 42.405 192.830 42.450 ;
        RECT 196.120 42.405 196.410 42.450 ;
        RECT 190.705 42.265 196.410 42.405 ;
        RECT 190.705 42.220 190.995 42.265 ;
        RECT 192.540 42.220 192.830 42.265 ;
        RECT 196.120 42.220 196.410 42.265 ;
        RECT 177.360 41.925 179.965 42.065 ;
        RECT 177.360 41.880 177.650 41.925 ;
        RECT 179.645 41.865 179.965 41.925 ;
        RECT 180.195 41.925 186.315 42.065 ;
        RECT 169.985 41.525 170.305 41.785 ;
        RECT 177.805 41.725 178.125 41.785 ;
        RECT 180.195 41.725 180.335 41.925 ;
        RECT 191.605 41.865 191.925 42.125 ;
        RECT 193.900 42.065 194.550 42.110 ;
        RECT 196.665 42.065 196.985 42.125 ;
        RECT 197.200 42.110 197.490 42.425 ;
        RECT 201.745 42.405 202.035 42.450 ;
        RECT 203.580 42.405 203.870 42.450 ;
        RECT 207.160 42.405 207.450 42.450 ;
        RECT 201.745 42.265 207.450 42.405 ;
        RECT 201.745 42.220 202.035 42.265 ;
        RECT 203.580 42.220 203.870 42.265 ;
        RECT 207.160 42.220 207.450 42.265 ;
        RECT 197.200 42.065 197.790 42.110 ;
        RECT 193.900 41.925 197.790 42.065 ;
        RECT 193.900 41.880 194.550 41.925 ;
        RECT 196.665 41.865 196.985 41.925 ;
        RECT 197.500 41.880 197.790 41.925 ;
        RECT 200.360 42.065 200.650 42.110 ;
        RECT 200.805 42.065 201.125 42.125 ;
        RECT 208.240 42.110 208.530 42.425 ;
        RECT 216.445 42.405 216.765 42.465 ;
        RECT 217.380 42.405 217.670 42.450 ;
        RECT 216.445 42.265 217.670 42.405 ;
        RECT 216.445 42.205 216.765 42.265 ;
        RECT 217.380 42.220 217.670 42.265 ;
        RECT 217.845 42.405 218.135 42.450 ;
        RECT 219.680 42.405 219.970 42.450 ;
        RECT 223.260 42.405 223.550 42.450 ;
        RECT 224.355 42.425 224.495 42.605 ;
        RECT 226.565 42.545 226.885 42.605 ;
        RECT 233.465 42.545 233.785 42.605 ;
        RECT 237.160 42.745 237.450 42.790 ;
        RECT 238.985 42.745 239.305 42.805 ;
        RECT 237.160 42.605 239.305 42.745 ;
        RECT 237.160 42.560 237.450 42.605 ;
        RECT 238.985 42.545 239.305 42.605 ;
        RECT 246.820 42.745 247.110 42.790 ;
        RECT 250.945 42.745 251.265 42.805 ;
        RECT 246.820 42.605 251.265 42.745 ;
        RECT 246.820 42.560 247.110 42.605 ;
        RECT 250.945 42.545 251.265 42.605 ;
        RECT 217.845 42.265 223.550 42.405 ;
        RECT 217.845 42.220 218.135 42.265 ;
        RECT 219.680 42.220 219.970 42.265 ;
        RECT 223.260 42.220 223.550 42.265 ;
        RECT 200.360 41.925 201.125 42.065 ;
        RECT 200.360 41.880 200.650 41.925 ;
        RECT 200.805 41.865 201.125 41.925 ;
        RECT 204.940 42.065 205.590 42.110 ;
        RECT 208.240 42.065 208.830 42.110 ;
        RECT 209.085 42.065 209.405 42.125 ;
        RECT 211.385 42.065 211.705 42.125 ;
        RECT 215.080 42.065 215.370 42.110 ;
        RECT 204.940 41.925 211.705 42.065 ;
        RECT 204.940 41.880 205.590 41.925 ;
        RECT 208.540 41.880 208.830 41.925 ;
        RECT 209.085 41.865 209.405 41.925 ;
        RECT 211.385 41.865 211.705 41.925 ;
        RECT 214.235 41.925 215.370 42.065 ;
        RECT 177.805 41.585 180.335 41.725 ;
        RECT 183.800 41.725 184.090 41.770 ;
        RECT 189.765 41.725 190.085 41.785 ;
        RECT 214.235 41.770 214.375 41.925 ;
        RECT 215.080 41.880 215.370 41.925 ;
        RECT 218.745 41.865 219.065 42.125 ;
        RECT 224.340 42.110 224.630 42.425 ;
        RECT 227.025 42.205 227.345 42.465 ;
        RECT 230.200 42.110 230.490 42.425 ;
        RECT 231.280 42.405 231.570 42.450 ;
        RECT 234.860 42.405 235.150 42.450 ;
        RECT 236.695 42.405 236.985 42.450 ;
        RECT 231.280 42.265 236.985 42.405 ;
        RECT 231.280 42.220 231.570 42.265 ;
        RECT 234.860 42.220 235.150 42.265 ;
        RECT 236.695 42.220 236.985 42.265 ;
        RECT 240.365 42.205 240.685 42.465 ;
        RECT 247.265 42.405 247.585 42.465 ;
        RECT 254.255 42.450 254.395 42.945 ;
        RECT 258.305 42.885 258.625 42.945 ;
        RECT 261.950 43.085 262.240 43.130 ;
        RECT 263.840 43.085 264.130 43.130 ;
        RECT 266.960 43.085 267.250 43.130 ;
        RECT 261.950 42.945 267.250 43.085 ;
        RECT 261.950 42.900 262.240 42.945 ;
        RECT 263.840 42.900 264.130 42.945 ;
        RECT 266.960 42.900 267.250 42.945 ;
        RECT 267.505 43.085 267.825 43.145 ;
        RECT 276.335 43.085 276.475 43.285 ;
        RECT 267.505 42.945 276.475 43.085 ;
        RECT 267.505 42.885 267.825 42.945 ;
        RECT 277.165 42.885 277.485 43.145 ;
        RECT 280.845 42.885 281.165 43.145 ;
        RECT 281.395 43.085 281.535 43.285 ;
        RECT 282.225 43.225 282.545 43.485 ;
        RECT 289.125 43.225 289.445 43.485 ;
        RECT 291.885 43.425 292.205 43.485 ;
        RECT 294.185 43.425 294.505 43.485 ;
        RECT 291.885 43.285 294.505 43.425 ;
        RECT 291.885 43.225 292.205 43.285 ;
        RECT 294.185 43.225 294.505 43.285 ;
        RECT 302.940 43.425 303.230 43.470 ;
        RECT 304.305 43.425 304.625 43.485 ;
        RECT 302.940 43.285 304.625 43.425 ;
        RECT 302.940 43.240 303.230 43.285 ;
        RECT 303.015 43.085 303.155 43.240 ;
        RECT 304.305 43.225 304.625 43.285 ;
        RECT 305.225 43.425 305.545 43.485 ;
        RECT 306.160 43.425 306.450 43.470 ;
        RECT 305.225 43.285 306.450 43.425 ;
        RECT 305.225 43.225 305.545 43.285 ;
        RECT 306.160 43.240 306.450 43.285 ;
        RECT 281.395 42.945 303.155 43.085 ;
        RECT 260.605 42.745 260.925 42.805 ;
        RECT 255.635 42.605 260.925 42.745 ;
        RECT 255.635 42.450 255.775 42.605 ;
        RECT 253.720 42.405 254.010 42.450 ;
        RECT 247.265 42.265 254.010 42.405 ;
        RECT 247.265 42.205 247.585 42.265 ;
        RECT 253.720 42.220 254.010 42.265 ;
        RECT 254.180 42.220 254.470 42.450 ;
        RECT 255.560 42.220 255.850 42.450 ;
        RECT 256.465 42.205 256.785 42.465 ;
        RECT 257.220 42.405 257.510 42.450 ;
        RECT 257.220 42.220 257.615 42.405 ;
        RECT 233.465 42.110 233.785 42.125 ;
        RECT 221.040 42.065 221.690 42.110 ;
        RECT 224.340 42.065 224.930 42.110 ;
        RECT 221.040 41.925 224.930 42.065 ;
        RECT 221.040 41.880 221.690 41.925 ;
        RECT 224.640 41.880 224.930 41.925 ;
        RECT 229.900 42.065 230.490 42.110 ;
        RECT 233.140 42.065 233.790 42.110 ;
        RECT 235.780 42.065 236.070 42.110 ;
        RECT 229.900 41.925 233.790 42.065 ;
        RECT 229.900 41.880 230.190 41.925 ;
        RECT 233.140 41.880 233.790 41.925 ;
        RECT 234.015 41.925 236.070 42.065 ;
        RECT 233.465 41.865 233.785 41.880 ;
        RECT 183.800 41.585 190.085 41.725 ;
        RECT 177.805 41.525 178.125 41.585 ;
        RECT 183.800 41.540 184.090 41.585 ;
        RECT 189.765 41.525 190.085 41.585 ;
        RECT 214.160 41.540 214.450 41.770 ;
        RECT 227.945 41.725 228.265 41.785 ;
        RECT 234.015 41.725 234.155 41.925 ;
        RECT 235.780 41.880 236.070 41.925 ;
        RECT 254.640 42.065 254.930 42.110 ;
        RECT 257.475 42.065 257.615 42.220 ;
        RECT 257.845 42.205 258.165 42.465 ;
        RECT 258.880 42.450 259.020 42.605 ;
        RECT 260.605 42.545 260.925 42.605 ;
        RECT 262.460 42.745 262.750 42.790 ;
        RECT 265.665 42.745 265.985 42.805 ;
        RECT 262.460 42.605 265.985 42.745 ;
        RECT 262.460 42.560 262.750 42.605 ;
        RECT 265.665 42.545 265.985 42.605 ;
        RECT 269.820 42.745 270.110 42.790 ;
        RECT 273.960 42.745 274.250 42.790 ;
        RECT 269.820 42.605 274.250 42.745 ;
        RECT 277.255 42.745 277.395 42.885 ;
        RECT 280.935 42.745 281.075 42.885 ;
        RECT 277.255 42.605 279.240 42.745 ;
        RECT 269.820 42.560 270.110 42.605 ;
        RECT 273.960 42.560 274.250 42.605 ;
        RECT 258.805 42.220 259.095 42.450 ;
        RECT 261.080 42.220 261.370 42.450 ;
        RECT 261.545 42.405 261.835 42.450 ;
        RECT 263.380 42.405 263.670 42.450 ;
        RECT 266.960 42.405 267.250 42.450 ;
        RECT 261.545 42.265 267.250 42.405 ;
        RECT 261.545 42.220 261.835 42.265 ;
        RECT 263.380 42.220 263.670 42.265 ;
        RECT 266.960 42.220 267.250 42.265 ;
        RECT 254.640 41.925 257.615 42.065 ;
        RECT 254.640 41.880 254.930 41.925 ;
        RECT 257.475 41.785 257.615 41.925 ;
        RECT 258.305 41.865 258.625 42.125 ;
        RECT 259.225 42.065 259.545 42.125 ;
        RECT 261.155 42.065 261.295 42.220 ;
        RECT 259.225 41.925 261.295 42.065 ;
        RECT 264.740 42.065 265.390 42.110 ;
        RECT 265.665 42.065 265.985 42.125 ;
        RECT 268.040 42.110 268.330 42.425 ;
        RECT 268.885 42.405 269.205 42.465 ;
        RECT 273.040 42.405 273.330 42.450 ;
        RECT 268.885 42.265 273.330 42.405 ;
        RECT 268.885 42.205 269.205 42.265 ;
        RECT 273.040 42.220 273.330 42.265 ;
        RECT 276.705 42.405 277.025 42.465 ;
        RECT 279.100 42.450 279.240 42.605 ;
        RECT 280.475 42.605 281.075 42.745 ;
        RECT 284.065 42.745 284.385 42.805 ;
        RECT 285.000 42.745 285.290 42.790 ;
        RECT 284.065 42.605 285.290 42.745 ;
        RECT 278.560 42.405 278.850 42.450 ;
        RECT 276.705 42.265 278.850 42.405 ;
        RECT 276.705 42.205 277.025 42.265 ;
        RECT 278.560 42.220 278.850 42.265 ;
        RECT 279.025 42.220 279.315 42.450 ;
        RECT 279.465 42.405 279.785 42.465 ;
        RECT 280.475 42.450 280.615 42.605 ;
        RECT 284.065 42.545 284.385 42.605 ;
        RECT 285.000 42.560 285.290 42.605 ;
        RECT 297.865 42.545 298.185 42.805 ;
        RECT 305.225 42.745 305.545 42.805 ;
        RECT 298.415 42.605 305.915 42.745 ;
        RECT 298.415 42.465 298.555 42.605 ;
        RECT 305.225 42.545 305.545 42.605 ;
        RECT 279.940 42.405 280.230 42.450 ;
        RECT 279.465 42.265 280.230 42.405 ;
        RECT 279.465 42.205 279.785 42.265 ;
        RECT 279.940 42.220 280.230 42.265 ;
        RECT 280.400 42.220 280.690 42.450 ;
        RECT 280.885 42.220 281.175 42.450 ;
        RECT 268.040 42.065 268.630 42.110 ;
        RECT 264.740 41.925 268.630 42.065 ;
        RECT 259.225 41.865 259.545 41.925 ;
        RECT 264.740 41.880 265.390 41.925 ;
        RECT 265.665 41.865 265.985 41.925 ;
        RECT 268.340 41.880 268.630 41.925 ;
        RECT 272.565 42.065 272.885 42.125 ;
        RECT 280.960 42.065 281.100 42.220 ;
        RECT 285.905 42.205 286.225 42.465 ;
        RECT 296.960 42.405 297.250 42.450 ;
        RECT 298.325 42.405 298.645 42.465 ;
        RECT 296.960 42.265 298.645 42.405 ;
        RECT 296.960 42.220 297.250 42.265 ;
        RECT 298.325 42.205 298.645 42.265 ;
        RECT 300.625 42.205 300.945 42.465 ;
        RECT 305.775 42.450 305.915 42.605 ;
        RECT 305.700 42.220 305.990 42.450 ;
        RECT 281.305 42.065 281.625 42.125 ;
        RECT 283.145 42.065 283.465 42.125 ;
        RECT 289.585 42.065 289.905 42.125 ;
        RECT 272.565 41.925 289.905 42.065 ;
        RECT 272.565 41.865 272.885 41.925 ;
        RECT 281.305 41.865 281.625 41.925 ;
        RECT 283.145 41.865 283.465 41.925 ;
        RECT 289.585 41.865 289.905 41.925 ;
        RECT 292.360 42.065 292.650 42.110 ;
        RECT 300.715 42.065 300.855 42.205 ;
        RECT 292.360 41.925 300.855 42.065 ;
        RECT 292.360 41.880 292.650 41.925 ;
        RECT 302.480 41.880 302.770 42.110 ;
        RECT 227.945 41.585 234.155 41.725 ;
        RECT 234.845 41.725 235.165 41.785 ;
        RECT 237.620 41.725 237.910 41.770 ;
        RECT 234.845 41.585 237.910 41.725 ;
        RECT 227.945 41.525 228.265 41.585 ;
        RECT 234.845 41.525 235.165 41.585 ;
        RECT 237.620 41.540 237.910 41.585 ;
        RECT 251.405 41.725 251.725 41.785 ;
        RECT 252.800 41.725 253.090 41.770 ;
        RECT 251.405 41.585 253.090 41.725 ;
        RECT 251.405 41.525 251.725 41.585 ;
        RECT 252.800 41.540 253.090 41.585 ;
        RECT 257.385 41.525 257.705 41.785 ;
        RECT 259.700 41.725 259.990 41.770 ;
        RECT 261.985 41.725 262.305 41.785 ;
        RECT 259.700 41.585 262.305 41.725 ;
        RECT 259.700 41.540 259.990 41.585 ;
        RECT 261.985 41.525 262.305 41.585 ;
        RECT 281.765 41.525 282.085 41.785 ;
        RECT 289.125 41.725 289.445 41.785 ;
        RECT 292.435 41.725 292.575 41.880 ;
        RECT 289.125 41.585 292.575 41.725 ;
        RECT 295.580 41.725 295.870 41.770 ;
        RECT 296.025 41.725 296.345 41.785 ;
        RECT 295.580 41.585 296.345 41.725 ;
        RECT 289.125 41.525 289.445 41.585 ;
        RECT 295.580 41.540 295.870 41.585 ;
        RECT 296.025 41.525 296.345 41.585 ;
        RECT 296.945 41.725 297.265 41.785 ;
        RECT 302.555 41.725 302.695 41.880 ;
        RECT 296.945 41.585 302.695 41.725 ;
        RECT 296.945 41.525 297.265 41.585 ;
        RECT 162.095 40.905 311.935 41.385 ;
        RECT 169.985 40.705 170.305 40.765 ;
        RECT 165.935 40.565 170.305 40.705 ;
        RECT 165.935 40.410 166.075 40.565 ;
        RECT 169.985 40.505 170.305 40.565 ;
        RECT 173.220 40.520 173.510 40.750 ;
        RECT 165.860 40.180 166.150 40.410 ;
        RECT 168.140 40.365 168.790 40.410 ;
        RECT 171.740 40.365 172.030 40.410 ;
        RECT 168.140 40.225 172.030 40.365 ;
        RECT 173.295 40.365 173.435 40.520 ;
        RECT 173.665 40.505 173.985 40.765 ;
        RECT 177.805 40.705 178.125 40.765 ;
        RECT 174.675 40.565 178.125 40.705 ;
        RECT 174.675 40.365 174.815 40.565 ;
        RECT 177.805 40.505 178.125 40.565 ;
        RECT 179.185 40.505 179.505 40.765 ;
        RECT 179.645 40.705 179.965 40.765 ;
        RECT 182.880 40.705 183.170 40.750 ;
        RECT 179.645 40.565 183.170 40.705 ;
        RECT 179.645 40.505 179.965 40.565 ;
        RECT 182.880 40.520 183.170 40.565 ;
        RECT 186.560 40.520 186.850 40.750 ;
        RECT 190.700 40.705 190.990 40.750 ;
        RECT 191.605 40.705 191.925 40.765 ;
        RECT 190.700 40.565 191.925 40.705 ;
        RECT 190.700 40.520 190.990 40.565 ;
        RECT 173.295 40.225 174.815 40.365 ;
        RECT 175.160 40.365 175.450 40.410 ;
        RECT 178.400 40.365 179.050 40.410 ;
        RECT 179.275 40.365 179.415 40.505 ;
        RECT 175.160 40.225 179.415 40.365 ;
        RECT 181.040 40.365 181.330 40.410 ;
        RECT 186.635 40.365 186.775 40.520 ;
        RECT 191.605 40.505 191.925 40.565 ;
        RECT 193.920 40.520 194.210 40.750 ;
        RECT 195.760 40.705 196.050 40.750 ;
        RECT 200.805 40.705 201.125 40.765 ;
        RECT 195.760 40.565 201.125 40.705 ;
        RECT 195.760 40.520 196.050 40.565 ;
        RECT 193.995 40.365 194.135 40.520 ;
        RECT 200.805 40.505 201.125 40.565 ;
        RECT 201.725 40.505 202.045 40.765 ;
        RECT 213.225 40.505 213.545 40.765 ;
        RECT 218.745 40.705 219.065 40.765 ;
        RECT 219.680 40.705 219.970 40.750 ;
        RECT 222.440 40.705 222.730 40.750 ;
        RECT 218.745 40.565 219.970 40.705 ;
        RECT 218.745 40.505 219.065 40.565 ;
        RECT 219.680 40.520 219.970 40.565 ;
        RECT 220.675 40.565 222.730 40.705 ;
        RECT 201.815 40.365 201.955 40.505 ;
        RECT 181.040 40.225 186.775 40.365 ;
        RECT 189.855 40.225 194.135 40.365 ;
        RECT 197.215 40.225 201.955 40.365 ;
        RECT 203.580 40.365 203.870 40.410 ;
        RECT 205.880 40.365 206.170 40.410 ;
        RECT 203.580 40.225 206.170 40.365 ;
        RECT 168.140 40.180 168.790 40.225 ;
        RECT 171.440 40.180 172.030 40.225 ;
        RECT 175.160 40.180 175.750 40.225 ;
        RECT 178.400 40.180 179.050 40.225 ;
        RECT 181.040 40.180 181.330 40.225 ;
        RECT 164.945 40.025 165.235 40.070 ;
        RECT 166.780 40.025 167.070 40.070 ;
        RECT 170.360 40.025 170.650 40.070 ;
        RECT 164.945 39.885 170.650 40.025 ;
        RECT 164.945 39.840 165.235 39.885 ;
        RECT 166.780 39.840 167.070 39.885 ;
        RECT 170.360 39.840 170.650 39.885 ;
        RECT 171.440 40.025 171.730 40.180 ;
        RECT 171.440 39.885 173.205 40.025 ;
        RECT 171.440 39.865 171.730 39.885 ;
        RECT 164.480 39.500 164.770 39.730 ;
        RECT 173.065 39.685 173.205 39.885 ;
        RECT 175.460 39.865 175.750 40.180 ;
        RECT 176.540 40.025 176.830 40.070 ;
        RECT 180.120 40.025 180.410 40.070 ;
        RECT 181.955 40.025 182.245 40.070 ;
        RECT 176.540 39.885 182.245 40.025 ;
        RECT 176.540 39.840 176.830 39.885 ;
        RECT 180.120 39.840 180.410 39.885 ;
        RECT 181.955 39.840 182.245 39.885 ;
        RECT 182.420 40.025 182.710 40.070 ;
        RECT 182.420 39.885 187.235 40.025 ;
        RECT 182.420 39.840 182.710 39.885 ;
        RECT 178.265 39.685 178.585 39.745 ;
        RECT 173.065 39.545 178.585 39.685 ;
        RECT 164.555 39.005 164.695 39.500 ;
        RECT 178.265 39.485 178.585 39.545 ;
        RECT 185.625 39.485 185.945 39.745 ;
        RECT 187.095 39.685 187.235 39.885 ;
        RECT 187.465 39.825 187.785 40.085 ;
        RECT 189.855 40.070 189.995 40.225 ;
        RECT 189.780 39.840 190.070 40.070 ;
        RECT 192.065 39.825 192.385 40.085 ;
        RECT 190.225 39.685 190.545 39.745 ;
        RECT 187.095 39.545 190.545 39.685 ;
        RECT 190.225 39.485 190.545 39.545 ;
        RECT 194.825 39.685 195.145 39.745 ;
        RECT 197.215 39.730 197.355 40.225 ;
        RECT 203.580 40.180 203.870 40.225 ;
        RECT 205.880 40.180 206.170 40.225 ;
        RECT 208.160 40.365 208.810 40.410 ;
        RECT 211.760 40.365 212.050 40.410 ;
        RECT 208.160 40.225 212.050 40.365 ;
        RECT 208.160 40.180 208.810 40.225 ;
        RECT 211.460 40.180 212.050 40.225 ;
        RECT 211.460 40.085 211.750 40.180 ;
        RECT 203.105 39.825 203.425 40.085 ;
        RECT 204.965 40.025 205.255 40.070 ;
        RECT 206.800 40.025 207.090 40.070 ;
        RECT 210.380 40.025 210.670 40.070 ;
        RECT 204.965 39.885 210.670 40.025 ;
        RECT 204.965 39.840 205.255 39.885 ;
        RECT 206.800 39.840 207.090 39.885 ;
        RECT 210.380 39.840 210.670 39.885 ;
        RECT 211.385 40.025 211.750 40.085 ;
        RECT 214.145 40.025 214.465 40.085 ;
        RECT 220.675 40.070 220.815 40.565 ;
        RECT 222.440 40.520 222.730 40.565 ;
        RECT 224.265 40.505 224.585 40.765 ;
        RECT 225.185 40.505 225.505 40.765 ;
        RECT 227.960 40.705 228.250 40.750 ;
        RECT 229.785 40.705 230.105 40.765 ;
        RECT 227.960 40.565 230.105 40.705 ;
        RECT 227.960 40.520 228.250 40.565 ;
        RECT 229.785 40.505 230.105 40.565 ;
        RECT 230.245 40.505 230.565 40.765 ;
        RECT 234.385 40.505 234.705 40.765 ;
        RECT 234.845 40.505 235.165 40.765 ;
        RECT 241.745 40.705 242.065 40.765 ;
        RECT 259.225 40.705 259.545 40.765 ;
        RECT 241.745 40.565 259.545 40.705 ;
        RECT 241.745 40.505 242.065 40.565 ;
        RECT 211.385 39.885 214.465 40.025 ;
        RECT 211.385 39.865 211.750 39.885 ;
        RECT 211.385 39.825 211.705 39.865 ;
        RECT 214.145 39.825 214.465 39.885 ;
        RECT 220.600 39.840 220.890 40.070 ;
        RECT 221.060 39.840 221.350 40.070 ;
        RECT 196.220 39.685 196.510 39.730 ;
        RECT 194.825 39.545 196.510 39.685 ;
        RECT 194.825 39.485 195.145 39.545 ;
        RECT 196.220 39.500 196.510 39.545 ;
        RECT 197.140 39.500 197.430 39.730 ;
        RECT 200.805 39.485 201.125 39.745 ;
        RECT 204.485 39.485 204.805 39.745 ;
        RECT 165.350 39.345 165.640 39.390 ;
        RECT 167.240 39.345 167.530 39.390 ;
        RECT 170.360 39.345 170.650 39.390 ;
        RECT 165.350 39.205 170.650 39.345 ;
        RECT 165.350 39.160 165.640 39.205 ;
        RECT 167.240 39.160 167.530 39.205 ;
        RECT 170.360 39.160 170.650 39.205 ;
        RECT 176.540 39.345 176.830 39.390 ;
        RECT 179.660 39.345 179.950 39.390 ;
        RECT 181.550 39.345 181.840 39.390 ;
        RECT 176.540 39.205 181.840 39.345 ;
        RECT 176.540 39.160 176.830 39.205 ;
        RECT 179.660 39.160 179.950 39.205 ;
        RECT 181.550 39.160 181.840 39.205 ;
        RECT 165.845 39.005 166.165 39.065 ;
        RECT 164.555 38.865 166.165 39.005 ;
        RECT 165.845 38.805 166.165 38.865 ;
        RECT 189.765 39.005 190.085 39.065 ;
        RECT 191.160 39.005 191.450 39.050 ;
        RECT 189.765 38.865 191.450 39.005 ;
        RECT 189.765 38.805 190.085 38.865 ;
        RECT 191.160 38.820 191.450 38.865 ;
        RECT 198.045 38.805 198.365 39.065 ;
        RECT 204.575 39.005 204.715 39.485 ;
        RECT 205.370 39.345 205.660 39.390 ;
        RECT 207.260 39.345 207.550 39.390 ;
        RECT 210.380 39.345 210.670 39.390 ;
        RECT 205.370 39.205 210.670 39.345 ;
        RECT 221.135 39.345 221.275 39.840 ;
        RECT 224.725 39.485 225.045 39.745 ;
        RECT 225.275 39.730 225.415 40.505 ;
        RECT 230.720 40.365 231.010 40.410 ;
        RECT 243.600 40.365 243.890 40.410 ;
        RECT 246.820 40.365 247.110 40.410 ;
        RECT 230.720 40.225 247.110 40.365 ;
        RECT 230.720 40.180 231.010 40.225 ;
        RECT 243.600 40.180 243.890 40.225 ;
        RECT 246.820 40.180 247.110 40.225 ;
        RECT 227.040 40.025 227.330 40.070 ;
        RECT 228.865 40.025 229.185 40.085 ;
        RECT 248.735 40.070 248.875 40.565 ;
        RECT 259.225 40.505 259.545 40.565 ;
        RECT 268.885 40.505 269.205 40.765 ;
        RECT 276.260 40.705 276.550 40.750 ;
        RECT 280.845 40.705 281.165 40.765 ;
        RECT 276.260 40.565 281.165 40.705 ;
        RECT 276.260 40.520 276.550 40.565 ;
        RECT 280.845 40.505 281.165 40.565 ;
        RECT 281.780 40.705 282.070 40.750 ;
        RECT 285.905 40.705 286.225 40.765 ;
        RECT 281.780 40.565 286.225 40.705 ;
        RECT 281.780 40.520 282.070 40.565 ;
        RECT 285.905 40.505 286.225 40.565 ;
        RECT 289.585 40.705 289.905 40.765 ;
        RECT 293.725 40.705 294.045 40.765 ;
        RECT 289.585 40.565 294.045 40.705 ;
        RECT 289.585 40.505 289.905 40.565 ;
        RECT 293.725 40.505 294.045 40.565 ;
        RECT 295.105 40.505 295.425 40.765 ;
        RECT 308.445 40.705 308.765 40.765 ;
        RECT 307.155 40.565 308.765 40.705 ;
        RECT 250.040 40.365 250.330 40.410 ;
        RECT 251.405 40.365 251.725 40.425 ;
        RECT 252.325 40.410 252.645 40.425 ;
        RECT 250.040 40.225 251.725 40.365 ;
        RECT 250.040 40.180 250.330 40.225 ;
        RECT 251.405 40.165 251.725 40.225 ;
        RECT 252.320 40.365 252.970 40.410 ;
        RECT 255.920 40.365 256.210 40.410 ;
        RECT 252.320 40.225 256.210 40.365 ;
        RECT 252.320 40.180 252.970 40.225 ;
        RECT 255.620 40.180 256.210 40.225 ;
        RECT 257.385 40.365 257.705 40.425 ;
        RECT 257.860 40.365 258.150 40.410 ;
        RECT 257.385 40.225 258.150 40.365 ;
        RECT 252.325 40.165 252.645 40.180 ;
        RECT 227.040 39.885 229.185 40.025 ;
        RECT 227.040 39.840 227.330 39.885 ;
        RECT 228.865 39.825 229.185 39.885 ;
        RECT 246.360 40.025 246.650 40.070 ;
        RECT 246.360 39.885 248.415 40.025 ;
        RECT 246.360 39.840 246.650 39.885 ;
        RECT 225.200 39.685 225.490 39.730 ;
        RECT 231.180 39.685 231.470 39.730 ;
        RECT 235.320 39.685 235.610 39.730 ;
        RECT 225.200 39.545 235.610 39.685 ;
        RECT 225.200 39.500 225.490 39.545 ;
        RECT 231.180 39.500 231.470 39.545 ;
        RECT 235.320 39.500 235.610 39.545 ;
        RECT 240.825 39.485 241.145 39.745 ;
        RECT 247.725 39.485 248.045 39.745 ;
        RECT 248.275 39.685 248.415 39.885 ;
        RECT 248.660 39.840 248.950 40.070 ;
        RECT 249.125 40.025 249.415 40.070 ;
        RECT 250.960 40.025 251.250 40.070 ;
        RECT 254.540 40.025 254.830 40.070 ;
        RECT 249.125 39.885 254.830 40.025 ;
        RECT 249.125 39.840 249.415 39.885 ;
        RECT 250.960 39.840 251.250 39.885 ;
        RECT 254.540 39.840 254.830 39.885 ;
        RECT 255.620 39.865 255.910 40.180 ;
        RECT 257.385 40.165 257.705 40.225 ;
        RECT 257.860 40.180 258.150 40.225 ;
        RECT 258.305 40.365 258.625 40.425 ;
        RECT 268.975 40.365 269.115 40.505 ;
        RECT 258.305 40.225 269.115 40.365 ;
        RECT 271.180 40.365 271.830 40.410 ;
        RECT 272.105 40.365 272.425 40.425 ;
        RECT 274.780 40.365 275.070 40.410 ;
        RECT 271.180 40.225 275.070 40.365 ;
        RECT 258.305 40.165 258.625 40.225 ;
        RECT 271.180 40.180 271.830 40.225 ;
        RECT 272.105 40.165 272.425 40.225 ;
        RECT 274.480 40.180 275.070 40.225 ;
        RECT 277.625 40.365 277.945 40.425 ;
        RECT 280.385 40.365 280.675 40.410 ;
        RECT 295.195 40.365 295.335 40.505 ;
        RECT 307.155 40.410 307.295 40.565 ;
        RECT 308.445 40.505 308.765 40.565 ;
        RECT 277.625 40.225 280.675 40.365 ;
        RECT 261.985 40.025 262.305 40.085 ;
        RECT 264.300 40.025 264.590 40.070 ;
        RECT 261.985 39.885 264.590 40.025 ;
        RECT 261.985 39.825 262.305 39.885 ;
        RECT 264.300 39.840 264.590 39.885 ;
        RECT 267.985 40.025 268.275 40.070 ;
        RECT 269.820 40.025 270.110 40.070 ;
        RECT 273.400 40.025 273.690 40.070 ;
        RECT 267.985 39.885 273.690 40.025 ;
        RECT 267.985 39.840 268.275 39.885 ;
        RECT 269.820 39.840 270.110 39.885 ;
        RECT 273.400 39.840 273.690 39.885 ;
        RECT 274.480 39.865 274.770 40.180 ;
        RECT 277.625 40.165 277.945 40.225 ;
        RECT 280.385 40.180 280.675 40.225 ;
        RECT 292.895 40.225 295.335 40.365 ;
        RECT 301.200 40.365 301.490 40.410 ;
        RECT 304.440 40.365 305.090 40.410 ;
        RECT 301.200 40.225 305.090 40.365 ;
        RECT 278.545 39.825 278.865 40.085 ;
        RECT 279.300 40.025 279.590 40.070 ;
        RECT 279.300 39.840 279.695 40.025 ;
        RECT 257.400 39.685 257.690 39.730 ;
        RECT 260.620 39.685 260.910 39.730 ;
        RECT 248.275 39.545 256.005 39.685 ;
        RECT 232.560 39.345 232.850 39.390 ;
        RECT 221.135 39.205 232.850 39.345 ;
        RECT 205.370 39.160 205.660 39.205 ;
        RECT 207.260 39.160 207.550 39.205 ;
        RECT 210.380 39.160 210.670 39.205 ;
        RECT 232.560 39.160 232.850 39.205 ;
        RECT 249.530 39.345 249.820 39.390 ;
        RECT 251.420 39.345 251.710 39.390 ;
        RECT 254.540 39.345 254.830 39.390 ;
        RECT 249.530 39.205 254.830 39.345 ;
        RECT 255.865 39.345 256.005 39.545 ;
        RECT 257.400 39.545 260.910 39.685 ;
        RECT 257.400 39.500 257.690 39.545 ;
        RECT 260.620 39.500 260.910 39.545 ;
        RECT 264.745 39.685 265.065 39.745 ;
        RECT 267.520 39.685 267.810 39.730 ;
        RECT 264.745 39.545 267.810 39.685 ;
        RECT 264.745 39.485 265.065 39.545 ;
        RECT 267.520 39.500 267.810 39.545 ;
        RECT 268.900 39.685 269.190 39.730 ;
        RECT 271.185 39.685 271.505 39.745 ;
        RECT 268.900 39.545 271.505 39.685 ;
        RECT 279.555 39.685 279.695 39.840 ;
        RECT 279.925 39.825 280.245 40.085 ;
        RECT 281.305 40.070 281.625 40.085 ;
        RECT 281.090 39.840 281.625 40.070 ;
        RECT 281.305 39.825 281.625 39.840 ;
        RECT 282.225 39.825 282.545 40.085 ;
        RECT 290.505 39.825 290.825 40.085 ;
        RECT 291.885 39.825 292.205 40.085 ;
        RECT 282.315 39.685 282.455 39.825 ;
        RECT 279.555 39.545 282.455 39.685 ;
        RECT 268.900 39.500 269.190 39.545 ;
        RECT 271.185 39.485 271.505 39.545 ;
        RECT 268.390 39.345 268.680 39.390 ;
        RECT 270.280 39.345 270.570 39.390 ;
        RECT 273.400 39.345 273.690 39.390 ;
        RECT 255.865 39.205 262.215 39.345 ;
        RECT 249.530 39.160 249.820 39.205 ;
        RECT 251.420 39.160 251.710 39.205 ;
        RECT 254.540 39.160 254.830 39.205 ;
        RECT 205.865 39.005 206.185 39.065 ;
        RECT 204.575 38.865 206.185 39.005 ;
        RECT 205.865 38.805 206.185 38.865 ;
        RECT 221.980 39.005 222.270 39.050 ;
        RECT 227.945 39.005 228.265 39.065 ;
        RECT 221.980 38.865 228.265 39.005 ;
        RECT 221.980 38.820 222.270 38.865 ;
        RECT 227.945 38.805 228.265 38.865 ;
        RECT 228.405 38.805 228.725 39.065 ;
        RECT 244.505 38.805 244.825 39.065 ;
        RECT 249.105 39.005 249.425 39.065 ;
        RECT 252.325 39.005 252.645 39.065 ;
        RECT 249.105 38.865 252.645 39.005 ;
        RECT 249.105 38.805 249.425 38.865 ;
        RECT 252.325 38.805 252.645 38.865 ;
        RECT 261.525 38.805 261.845 39.065 ;
        RECT 262.075 39.005 262.215 39.205 ;
        RECT 268.390 39.205 273.690 39.345 ;
        RECT 268.390 39.160 268.680 39.205 ;
        RECT 270.280 39.160 270.570 39.205 ;
        RECT 273.400 39.160 273.690 39.205 ;
        RECT 279.925 39.345 280.245 39.405 ;
        RECT 292.895 39.390 293.035 40.225 ;
        RECT 301.200 40.180 301.790 40.225 ;
        RECT 304.440 40.180 305.090 40.225 ;
        RECT 307.080 40.180 307.370 40.410 ;
        RECT 295.105 39.825 295.425 40.085 ;
        RECT 301.500 40.025 301.790 40.180 ;
        RECT 302.005 40.025 302.325 40.085 ;
        RECT 301.500 39.885 302.325 40.025 ;
        RECT 301.500 39.865 301.790 39.885 ;
        RECT 302.005 39.825 302.325 39.885 ;
        RECT 302.580 40.025 302.870 40.070 ;
        RECT 306.160 40.025 306.450 40.070 ;
        RECT 307.995 40.025 308.285 40.070 ;
        RECT 302.580 39.885 308.285 40.025 ;
        RECT 302.580 39.840 302.870 39.885 ;
        RECT 306.160 39.840 306.450 39.885 ;
        RECT 307.995 39.840 308.285 39.885 ;
        RECT 308.460 40.025 308.750 40.070 ;
        RECT 308.905 40.025 309.225 40.085 ;
        RECT 308.460 39.885 309.225 40.025 ;
        RECT 308.460 39.840 308.750 39.885 ;
        RECT 308.905 39.825 309.225 39.885 ;
        RECT 296.485 39.485 296.805 39.745 ;
        RECT 292.820 39.345 293.110 39.390 ;
        RECT 279.925 39.205 293.110 39.345 ;
        RECT 279.925 39.145 280.245 39.205 ;
        RECT 292.820 39.160 293.110 39.205 ;
        RECT 302.580 39.345 302.870 39.390 ;
        RECT 305.700 39.345 305.990 39.390 ;
        RECT 307.590 39.345 307.880 39.390 ;
        RECT 302.580 39.205 307.880 39.345 ;
        RECT 302.580 39.160 302.870 39.205 ;
        RECT 305.700 39.160 305.990 39.205 ;
        RECT 307.590 39.160 307.880 39.205 ;
        RECT 270.725 39.005 271.045 39.065 ;
        RECT 262.075 38.865 271.045 39.005 ;
        RECT 270.725 38.805 271.045 38.865 ;
        RECT 299.705 38.805 300.025 39.065 ;
        RECT 162.095 38.185 311.135 38.665 ;
        RECT 180.120 37.985 180.410 38.030 ;
        RECT 187.465 37.985 187.785 38.045 ;
        RECT 180.120 37.845 187.785 37.985 ;
        RECT 180.120 37.800 180.410 37.845 ;
        RECT 187.465 37.785 187.785 37.845 ;
        RECT 195.760 37.985 196.050 38.030 ;
        RECT 200.805 37.985 201.125 38.045 ;
        RECT 195.760 37.845 201.125 37.985 ;
        RECT 195.760 37.800 196.050 37.845 ;
        RECT 200.805 37.785 201.125 37.845 ;
        RECT 212.765 37.985 213.085 38.045 ;
        RECT 214.620 37.985 214.910 38.030 ;
        RECT 212.765 37.845 214.910 37.985 ;
        RECT 212.765 37.785 213.085 37.845 ;
        RECT 214.620 37.800 214.910 37.845 ;
        RECT 224.725 37.985 225.045 38.045 ;
        RECT 227.040 37.985 227.330 38.030 ;
        RECT 224.725 37.845 227.330 37.985 ;
        RECT 224.725 37.785 225.045 37.845 ;
        RECT 227.040 37.800 227.330 37.845 ;
        RECT 228.865 37.985 229.185 38.045 ;
        RECT 230.720 37.985 231.010 38.030 ;
        RECT 228.865 37.845 231.010 37.985 ;
        RECT 228.865 37.785 229.185 37.845 ;
        RECT 230.720 37.800 231.010 37.845 ;
        RECT 240.825 37.985 241.145 38.045 ;
        RECT 241.300 37.985 241.590 38.030 ;
        RECT 247.725 37.985 248.045 38.045 ;
        RECT 240.825 37.845 241.590 37.985 ;
        RECT 240.825 37.785 241.145 37.845 ;
        RECT 241.300 37.800 241.590 37.845 ;
        RECT 241.835 37.845 248.045 37.985 ;
        RECT 166.730 37.645 167.020 37.690 ;
        RECT 168.620 37.645 168.910 37.690 ;
        RECT 171.740 37.645 172.030 37.690 ;
        RECT 166.730 37.505 172.030 37.645 ;
        RECT 166.730 37.460 167.020 37.505 ;
        RECT 168.620 37.460 168.910 37.505 ;
        RECT 171.740 37.460 172.030 37.505 ;
        RECT 174.600 37.645 174.890 37.690 ;
        RECT 185.625 37.645 185.945 37.705 ;
        RECT 174.600 37.505 185.945 37.645 ;
        RECT 174.600 37.460 174.890 37.505 ;
        RECT 185.625 37.445 185.945 37.505 ;
        RECT 187.890 37.645 188.180 37.690 ;
        RECT 189.780 37.645 190.070 37.690 ;
        RECT 192.900 37.645 193.190 37.690 ;
        RECT 187.890 37.505 193.190 37.645 ;
        RECT 187.890 37.460 188.180 37.505 ;
        RECT 189.780 37.460 190.070 37.505 ;
        RECT 192.900 37.460 193.190 37.505 ;
        RECT 206.750 37.645 207.040 37.690 ;
        RECT 208.640 37.645 208.930 37.690 ;
        RECT 211.760 37.645 212.050 37.690 ;
        RECT 241.835 37.645 241.975 37.845 ;
        RECT 247.725 37.785 248.045 37.845 ;
        RECT 253.705 37.985 254.025 38.045 ;
        RECT 267.520 37.985 267.810 38.030 ;
        RECT 253.705 37.845 267.810 37.985 ;
        RECT 253.705 37.785 254.025 37.845 ;
        RECT 267.520 37.800 267.810 37.845 ;
        RECT 271.185 37.785 271.505 38.045 ;
        RECT 283.605 37.985 283.925 38.045 ;
        RECT 285.000 37.985 285.290 38.030 ;
        RECT 289.585 37.985 289.905 38.045 ;
        RECT 283.605 37.845 289.905 37.985 ;
        RECT 283.605 37.785 283.925 37.845 ;
        RECT 285.000 37.800 285.290 37.845 ;
        RECT 289.585 37.785 289.905 37.845 ;
        RECT 295.105 37.985 295.425 38.045 ;
        RECT 296.500 37.985 296.790 38.030 ;
        RECT 295.105 37.845 296.790 37.985 ;
        RECT 295.105 37.785 295.425 37.845 ;
        RECT 296.500 37.800 296.790 37.845 ;
        RECT 305.225 37.985 305.545 38.045 ;
        RECT 305.700 37.985 305.990 38.030 ;
        RECT 305.225 37.845 305.990 37.985 ;
        RECT 305.225 37.785 305.545 37.845 ;
        RECT 305.700 37.800 305.990 37.845 ;
        RECT 206.750 37.505 212.050 37.645 ;
        RECT 206.750 37.460 207.040 37.505 ;
        RECT 208.640 37.460 208.930 37.505 ;
        RECT 211.760 37.460 212.050 37.505 ;
        RECT 234.015 37.505 241.975 37.645 ;
        RECT 244.160 37.645 244.450 37.690 ;
        RECT 247.280 37.645 247.570 37.690 ;
        RECT 249.170 37.645 249.460 37.690 ;
        RECT 244.160 37.505 249.460 37.645 ;
        RECT 176.885 37.305 177.205 37.365 ;
        RECT 177.360 37.305 177.650 37.350 ;
        RECT 176.885 37.165 177.650 37.305 ;
        RECT 176.885 37.105 177.205 37.165 ;
        RECT 177.360 37.120 177.650 37.165 ;
        RECT 177.820 37.305 178.110 37.350 ;
        RECT 178.725 37.305 179.045 37.365 ;
        RECT 177.820 37.165 179.045 37.305 ;
        RECT 177.820 37.120 178.110 37.165 ;
        RECT 165.845 36.765 166.165 37.025 ;
        RECT 166.325 36.965 166.615 37.010 ;
        RECT 168.160 36.965 168.450 37.010 ;
        RECT 171.740 36.965 172.030 37.010 ;
        RECT 166.325 36.825 172.030 36.965 ;
        RECT 166.325 36.780 166.615 36.825 ;
        RECT 168.160 36.780 168.450 36.825 ;
        RECT 171.740 36.780 172.030 36.825 ;
        RECT 167.225 36.425 167.545 36.685 ;
        RECT 172.820 36.670 173.110 36.985 ;
        RECT 177.435 36.965 177.575 37.120 ;
        RECT 178.725 37.105 179.045 37.165 ;
        RECT 179.645 37.105 179.965 37.365 ;
        RECT 187.020 37.305 187.310 37.350 ;
        RECT 190.225 37.305 190.545 37.365 ;
        RECT 187.020 37.165 190.545 37.305 ;
        RECT 187.020 37.120 187.310 37.165 ;
        RECT 190.225 37.105 190.545 37.165 ;
        RECT 205.865 37.105 206.185 37.365 ;
        RECT 225.645 37.305 225.965 37.365 ;
        RECT 234.015 37.350 234.155 37.505 ;
        RECT 244.160 37.460 244.450 37.505 ;
        RECT 247.280 37.460 247.570 37.505 ;
        RECT 249.170 37.460 249.460 37.505 ;
        RECT 257.040 37.645 257.330 37.690 ;
        RECT 260.160 37.645 260.450 37.690 ;
        RECT 262.050 37.645 262.340 37.690 ;
        RECT 257.040 37.505 262.340 37.645 ;
        RECT 257.040 37.460 257.330 37.505 ;
        RECT 260.160 37.460 260.450 37.505 ;
        RECT 262.050 37.460 262.340 37.505 ;
        RECT 274.495 37.505 281.995 37.645 ;
        RECT 233.940 37.305 234.230 37.350 ;
        RECT 225.645 37.165 234.230 37.305 ;
        RECT 225.645 37.105 225.965 37.165 ;
        RECT 233.940 37.120 234.230 37.165 ;
        RECT 234.845 37.105 235.165 37.365 ;
        RECT 241.745 37.305 242.065 37.365 ;
        RECT 248.660 37.305 248.950 37.350 ;
        RECT 261.065 37.305 261.385 37.365 ;
        RECT 262.920 37.305 263.210 37.350 ;
        RECT 264.745 37.305 265.065 37.365 ;
        RECT 274.495 37.350 274.635 37.505 ;
        RECT 281.855 37.365 281.995 37.505 ;
        RECT 282.225 37.445 282.545 37.705 ;
        RECT 287.250 37.645 287.540 37.690 ;
        RECT 289.140 37.645 289.430 37.690 ;
        RECT 292.260 37.645 292.550 37.690 ;
        RECT 284.155 37.505 286.135 37.645 ;
        RECT 241.745 37.165 248.950 37.305 ;
        RECT 241.745 37.105 242.065 37.165 ;
        RECT 248.660 37.120 248.950 37.165 ;
        RECT 250.115 37.165 265.065 37.305 ;
        RECT 179.735 36.965 179.875 37.105 ;
        RECT 177.435 36.825 179.875 36.965 ;
        RECT 183.325 36.765 183.645 37.025 ;
        RECT 187.485 36.965 187.775 37.010 ;
        RECT 189.320 36.965 189.610 37.010 ;
        RECT 192.900 36.965 193.190 37.010 ;
        RECT 187.485 36.825 193.190 36.965 ;
        RECT 187.485 36.780 187.775 36.825 ;
        RECT 189.320 36.780 189.610 36.825 ;
        RECT 192.900 36.780 193.190 36.825 ;
        RECT 169.520 36.625 170.170 36.670 ;
        RECT 172.820 36.625 173.410 36.670 ;
        RECT 177.805 36.625 178.125 36.685 ;
        RECT 169.520 36.485 178.125 36.625 ;
        RECT 169.520 36.440 170.170 36.485 ;
        RECT 173.120 36.440 173.410 36.485 ;
        RECT 177.805 36.425 178.125 36.485 ;
        RECT 178.265 36.625 178.585 36.685 ;
        RECT 180.580 36.625 180.870 36.670 ;
        RECT 178.265 36.485 180.870 36.625 ;
        RECT 178.265 36.425 178.585 36.485 ;
        RECT 180.580 36.440 180.870 36.485 ;
        RECT 188.400 36.625 188.690 36.670 ;
        RECT 189.765 36.625 190.085 36.685 ;
        RECT 193.980 36.670 194.270 36.985 ;
        RECT 197.585 36.965 197.905 37.025 ;
        RECT 199.900 36.965 200.190 37.010 ;
        RECT 197.585 36.825 200.190 36.965 ;
        RECT 197.585 36.765 197.905 36.825 ;
        RECT 199.900 36.780 200.190 36.825 ;
        RECT 206.345 36.965 206.635 37.010 ;
        RECT 208.180 36.965 208.470 37.010 ;
        RECT 211.760 36.965 212.050 37.010 ;
        RECT 206.345 36.825 212.050 36.965 ;
        RECT 206.345 36.780 206.635 36.825 ;
        RECT 208.180 36.780 208.470 36.825 ;
        RECT 211.760 36.780 212.050 36.825 ;
        RECT 188.400 36.485 190.085 36.625 ;
        RECT 188.400 36.440 188.690 36.485 ;
        RECT 189.765 36.425 190.085 36.485 ;
        RECT 190.680 36.625 191.330 36.670 ;
        RECT 193.980 36.625 194.570 36.670 ;
        RECT 200.345 36.625 200.665 36.685 ;
        RECT 190.680 36.485 200.665 36.625 ;
        RECT 190.680 36.440 191.330 36.485 ;
        RECT 194.280 36.440 194.570 36.485 ;
        RECT 200.345 36.425 200.665 36.485 ;
        RECT 207.245 36.425 207.565 36.685 ;
        RECT 212.840 36.670 213.130 36.985 ;
        RECT 221.505 36.765 221.825 37.025 ;
        RECT 222.885 36.965 223.205 37.025 ;
        RECT 224.740 36.965 225.030 37.010 ;
        RECT 222.885 36.825 225.030 36.965 ;
        RECT 222.885 36.765 223.205 36.825 ;
        RECT 224.740 36.780 225.030 36.825 ;
        RECT 230.245 36.765 230.565 37.025 ;
        RECT 232.545 36.765 232.865 37.025 ;
        RECT 233.020 36.965 233.310 37.010 ;
        RECT 234.935 36.965 235.075 37.105 ;
        RECT 233.020 36.825 235.075 36.965 ;
        RECT 236.240 36.965 236.530 37.010 ;
        RECT 238.525 36.965 238.845 37.025 ;
        RECT 250.115 37.010 250.255 37.165 ;
        RECT 261.065 37.105 261.385 37.165 ;
        RECT 262.920 37.120 263.210 37.165 ;
        RECT 264.745 37.105 265.065 37.165 ;
        RECT 274.420 37.120 274.710 37.350 ;
        RECT 278.085 37.305 278.405 37.365 ;
        RECT 274.955 37.165 277.855 37.305 ;
        RECT 240.380 36.965 240.670 37.010 ;
        RECT 236.240 36.825 240.670 36.965 ;
        RECT 233.020 36.780 233.310 36.825 ;
        RECT 236.240 36.780 236.530 36.825 ;
        RECT 238.525 36.765 238.845 36.825 ;
        RECT 240.380 36.780 240.670 36.825 ;
        RECT 209.540 36.625 210.190 36.670 ;
        RECT 212.840 36.625 213.430 36.670 ;
        RECT 214.145 36.625 214.465 36.685 ;
        RECT 220.125 36.625 220.445 36.685 ;
        RECT 243.080 36.670 243.370 36.985 ;
        RECT 244.160 36.965 244.450 37.010 ;
        RECT 247.740 36.965 248.030 37.010 ;
        RECT 249.575 36.965 249.865 37.010 ;
        RECT 244.160 36.825 249.865 36.965 ;
        RECT 244.160 36.780 244.450 36.825 ;
        RECT 247.740 36.780 248.030 36.825 ;
        RECT 249.575 36.780 249.865 36.825 ;
        RECT 250.040 36.780 250.330 37.010 ;
        RECT 252.325 36.965 252.645 37.025 ;
        RECT 255.085 36.965 255.405 37.025 ;
        RECT 255.960 36.965 256.250 36.985 ;
        RECT 252.325 36.825 256.250 36.965 ;
        RECT 209.540 36.485 220.445 36.625 ;
        RECT 209.540 36.440 210.190 36.485 ;
        RECT 213.140 36.440 213.430 36.485 ;
        RECT 194.825 36.285 195.145 36.345 ;
        RECT 197.140 36.285 197.430 36.330 ;
        RECT 194.825 36.145 197.430 36.285 ;
        RECT 194.825 36.085 195.145 36.145 ;
        RECT 197.140 36.100 197.430 36.145 ;
        RECT 212.305 36.285 212.625 36.345 ;
        RECT 213.775 36.285 213.915 36.485 ;
        RECT 214.145 36.425 214.465 36.485 ;
        RECT 220.125 36.425 220.445 36.485 ;
        RECT 242.780 36.625 243.370 36.670 ;
        RECT 246.020 36.625 246.670 36.670 ;
        RECT 249.105 36.625 249.425 36.685 ;
        RECT 242.780 36.485 249.425 36.625 ;
        RECT 242.780 36.440 243.070 36.485 ;
        RECT 246.020 36.440 246.670 36.485 ;
        RECT 249.105 36.425 249.425 36.485 ;
        RECT 212.305 36.145 213.915 36.285 ;
        RECT 212.305 36.085 212.625 36.145 ;
        RECT 220.585 36.085 220.905 36.345 ;
        RECT 221.045 36.285 221.365 36.345 ;
        RECT 221.980 36.285 222.270 36.330 ;
        RECT 221.045 36.145 222.270 36.285 ;
        RECT 221.045 36.085 221.365 36.145 ;
        RECT 221.980 36.100 222.270 36.145 ;
        RECT 238.065 36.085 238.385 36.345 ;
        RECT 242.205 36.285 242.525 36.345 ;
        RECT 250.115 36.285 250.255 36.780 ;
        RECT 252.325 36.765 252.645 36.825 ;
        RECT 255.085 36.765 255.405 36.825 ;
        RECT 255.960 36.670 256.250 36.825 ;
        RECT 257.040 36.965 257.330 37.010 ;
        RECT 260.620 36.965 260.910 37.010 ;
        RECT 262.455 36.965 262.745 37.010 ;
        RECT 257.040 36.825 262.745 36.965 ;
        RECT 257.040 36.780 257.330 36.825 ;
        RECT 260.620 36.780 260.910 36.825 ;
        RECT 262.455 36.780 262.745 36.825 ;
        RECT 266.140 36.965 266.430 37.010 ;
        RECT 266.140 36.825 269.805 36.965 ;
        RECT 266.140 36.780 266.430 36.825 ;
        RECT 255.660 36.625 256.250 36.670 ;
        RECT 258.900 36.625 259.550 36.670 ;
        RECT 255.660 36.485 259.550 36.625 ;
        RECT 255.660 36.440 255.950 36.485 ;
        RECT 258.900 36.440 259.550 36.485 ;
        RECT 261.525 36.425 261.845 36.685 ;
        RECT 269.665 36.625 269.805 36.825 ;
        RECT 270.725 36.765 271.045 37.025 ;
        RECT 274.955 37.010 275.095 37.165 ;
        RECT 274.880 36.780 275.170 37.010 ;
        RECT 272.565 36.625 272.885 36.685 ;
        RECT 269.665 36.485 272.885 36.625 ;
        RECT 272.565 36.425 272.885 36.485 ;
        RECT 242.205 36.145 250.255 36.285 ;
        RECT 254.180 36.285 254.470 36.330 ;
        RECT 258.305 36.285 258.625 36.345 ;
        RECT 254.180 36.145 258.625 36.285 ;
        RECT 242.205 36.085 242.525 36.145 ;
        RECT 254.180 36.100 254.470 36.145 ;
        RECT 258.305 36.085 258.625 36.145 ;
        RECT 267.045 36.085 267.365 36.345 ;
        RECT 269.805 36.285 270.125 36.345 ;
        RECT 274.955 36.285 275.095 36.780 ;
        RECT 276.245 36.765 276.565 37.025 ;
        RECT 277.715 36.965 277.855 37.165 ;
        RECT 278.085 37.165 278.775 37.305 ;
        RECT 278.085 37.105 278.405 37.165 ;
        RECT 278.635 36.965 278.775 37.165 ;
        RECT 281.765 37.105 282.085 37.365 ;
        RECT 284.155 37.305 284.295 37.505 ;
        RECT 283.235 37.165 284.295 37.305 ;
        RECT 282.240 36.965 282.530 37.010 ;
        RECT 277.715 36.825 278.315 36.965 ;
        RECT 278.635 36.825 282.530 36.965 ;
        RECT 275.340 36.625 275.630 36.670 ;
        RECT 278.175 36.625 278.315 36.825 ;
        RECT 282.240 36.780 282.530 36.825 ;
        RECT 279.465 36.625 279.785 36.685 ;
        RECT 275.340 36.485 277.855 36.625 ;
        RECT 278.175 36.485 279.785 36.625 ;
        RECT 275.340 36.440 275.630 36.485 ;
        RECT 269.805 36.145 275.095 36.285 ;
        RECT 269.805 36.085 270.125 36.145 ;
        RECT 277.165 36.085 277.485 36.345 ;
        RECT 277.715 36.285 277.855 36.485 ;
        RECT 279.465 36.425 279.785 36.485 ;
        RECT 279.925 36.625 280.245 36.685 ;
        RECT 283.235 36.670 283.375 37.165 ;
        RECT 283.605 36.765 283.925 37.025 ;
        RECT 285.995 36.685 286.135 37.505 ;
        RECT 287.250 37.505 292.550 37.645 ;
        RECT 287.250 37.460 287.540 37.505 ;
        RECT 289.140 37.460 289.430 37.505 ;
        RECT 292.260 37.460 292.550 37.505 ;
        RECT 295.580 37.460 295.870 37.690 ;
        RECT 296.025 37.645 296.345 37.705 ;
        RECT 302.005 37.645 302.325 37.705 ;
        RECT 296.025 37.505 302.325 37.645 ;
        RECT 290.505 37.305 290.825 37.365 ;
        RECT 295.655 37.305 295.795 37.460 ;
        RECT 296.025 37.445 296.345 37.505 ;
        RECT 302.005 37.445 302.325 37.505 ;
        RECT 290.505 37.165 295.795 37.305 ;
        RECT 290.505 37.105 290.825 37.165 ;
        RECT 286.365 36.765 286.685 37.025 ;
        RECT 286.845 36.965 287.135 37.010 ;
        RECT 288.680 36.965 288.970 37.010 ;
        RECT 292.260 36.965 292.550 37.010 ;
        RECT 286.845 36.825 292.550 36.965 ;
        RECT 286.845 36.780 287.135 36.825 ;
        RECT 288.680 36.780 288.970 36.825 ;
        RECT 292.260 36.780 292.550 36.825 ;
        RECT 293.340 36.965 293.630 36.985 ;
        RECT 296.115 36.965 296.255 37.445 ;
        RECT 296.485 37.105 296.805 37.365 ;
        RECT 299.705 37.305 300.025 37.365 ;
        RECT 300.180 37.305 300.470 37.350 ;
        RECT 299.705 37.165 300.470 37.305 ;
        RECT 299.705 37.105 300.025 37.165 ;
        RECT 300.180 37.120 300.470 37.165 ;
        RECT 293.340 36.825 296.255 36.965 ;
        RECT 296.575 36.965 296.715 37.105 ;
        RECT 304.305 36.965 304.625 37.025 ;
        RECT 306.160 36.965 306.450 37.010 ;
        RECT 296.575 36.825 299.935 36.965 ;
        RECT 280.400 36.625 280.690 36.670 ;
        RECT 279.925 36.485 280.690 36.625 ;
        RECT 279.925 36.425 280.245 36.485 ;
        RECT 280.400 36.440 280.690 36.485 ;
        RECT 283.160 36.440 283.450 36.670 ;
        RECT 285.905 36.425 286.225 36.685 ;
        RECT 293.340 36.670 293.630 36.825 ;
        RECT 287.760 36.440 288.050 36.670 ;
        RECT 290.040 36.625 290.690 36.670 ;
        RECT 293.340 36.625 293.930 36.670 ;
        RECT 290.040 36.485 293.930 36.625 ;
        RECT 290.040 36.440 290.690 36.485 ;
        RECT 293.640 36.440 293.930 36.485 ;
        RECT 280.015 36.285 280.155 36.425 ;
        RECT 277.715 36.145 280.155 36.285 ;
        RECT 281.305 36.085 281.625 36.345 ;
        RECT 283.605 36.285 283.925 36.345 ;
        RECT 284.080 36.285 284.370 36.330 ;
        RECT 283.605 36.145 284.370 36.285 ;
        RECT 283.605 36.085 283.925 36.145 ;
        RECT 284.080 36.100 284.370 36.145 ;
        RECT 284.920 36.285 285.210 36.330 ;
        RECT 287.835 36.285 287.975 36.440 ;
        RECT 295.105 36.425 295.425 36.685 ;
        RECT 296.575 36.670 296.715 36.825 ;
        RECT 296.420 36.485 296.715 36.670 ;
        RECT 296.420 36.440 296.710 36.485 ;
        RECT 297.420 36.440 297.710 36.670 ;
        RECT 297.880 36.625 298.170 36.670 ;
        RECT 298.325 36.625 298.645 36.685 ;
        RECT 297.880 36.485 298.645 36.625 ;
        RECT 297.880 36.440 298.170 36.485 ;
        RECT 295.195 36.285 295.335 36.425 ;
        RECT 297.495 36.285 297.635 36.440 ;
        RECT 298.325 36.425 298.645 36.485 ;
        RECT 298.785 36.425 299.105 36.685 ;
        RECT 299.795 36.670 299.935 36.825 ;
        RECT 304.305 36.825 306.450 36.965 ;
        RECT 304.305 36.765 304.625 36.825 ;
        RECT 306.160 36.780 306.450 36.825 ;
        RECT 299.720 36.440 300.010 36.670 ;
        RECT 284.920 36.145 297.635 36.285 ;
        RECT 284.920 36.100 285.210 36.145 ;
        RECT 303.385 36.085 303.705 36.345 ;
        RECT 162.095 35.465 311.935 35.945 ;
        RECT 165.845 35.265 166.165 35.325 ;
        RECT 177.345 35.265 177.665 35.325 ;
        RECT 165.845 35.125 177.665 35.265 ;
        RECT 165.845 35.065 166.165 35.125 ;
        RECT 167.315 34.630 167.455 35.125 ;
        RECT 177.345 35.065 177.665 35.125 ;
        RECT 178.265 35.065 178.585 35.325 ;
        RECT 178.740 35.265 179.030 35.310 ;
        RECT 179.185 35.265 179.505 35.325 ;
        RECT 178.740 35.125 179.505 35.265 ;
        RECT 178.740 35.080 179.030 35.125 ;
        RECT 179.185 35.065 179.505 35.125 ;
        RECT 183.325 35.065 183.645 35.325 ;
        RECT 192.065 35.265 192.385 35.325 ;
        RECT 193.460 35.265 193.750 35.310 ;
        RECT 192.065 35.125 193.750 35.265 ;
        RECT 192.065 35.065 192.385 35.125 ;
        RECT 193.460 35.080 193.750 35.125 ;
        RECT 204.025 35.065 204.345 35.325 ;
        RECT 207.245 35.265 207.565 35.325 ;
        RECT 208.180 35.265 208.470 35.310 ;
        RECT 207.245 35.125 208.470 35.265 ;
        RECT 207.245 35.065 207.565 35.125 ;
        RECT 208.180 35.080 208.470 35.125 ;
        RECT 209.545 35.065 209.865 35.325 ;
        RECT 211.400 35.265 211.690 35.310 ;
        RECT 212.765 35.265 213.085 35.325 ;
        RECT 211.400 35.125 213.085 35.265 ;
        RECT 211.400 35.080 211.690 35.125 ;
        RECT 212.765 35.065 213.085 35.125 ;
        RECT 220.600 35.265 220.890 35.310 ;
        RECT 221.045 35.265 221.365 35.325 ;
        RECT 220.600 35.125 221.365 35.265 ;
        RECT 220.600 35.080 220.890 35.125 ;
        RECT 221.045 35.065 221.365 35.125 ;
        RECT 221.505 35.265 221.825 35.325 ;
        RECT 222.440 35.265 222.730 35.310 ;
        RECT 221.505 35.125 222.730 35.265 ;
        RECT 221.505 35.065 221.825 35.125 ;
        RECT 222.440 35.080 222.730 35.125 ;
        RECT 224.725 35.065 225.045 35.325 ;
        RECT 225.645 35.065 225.965 35.325 ;
        RECT 238.065 35.265 238.385 35.325 ;
        RECT 227.575 35.125 232.315 35.265 ;
        RECT 170.900 34.925 171.550 34.970 ;
        RECT 174.500 34.925 174.790 34.970 ;
        RECT 177.805 34.925 178.125 34.985 ;
        RECT 170.900 34.785 178.125 34.925 ;
        RECT 170.900 34.740 171.550 34.785 ;
        RECT 174.200 34.740 174.790 34.785 ;
        RECT 167.240 34.400 167.530 34.630 ;
        RECT 167.705 34.585 167.995 34.630 ;
        RECT 169.540 34.585 169.830 34.630 ;
        RECT 173.120 34.585 173.410 34.630 ;
        RECT 167.705 34.445 173.410 34.585 ;
        RECT 167.705 34.400 167.995 34.445 ;
        RECT 169.540 34.400 169.830 34.445 ;
        RECT 173.120 34.400 173.410 34.445 ;
        RECT 174.200 34.425 174.490 34.740 ;
        RECT 177.805 34.725 178.125 34.785 ;
        RECT 183.415 34.585 183.555 35.065 ;
        RECT 191.160 34.925 191.450 34.970 ;
        RECT 198.045 34.925 198.365 34.985 ;
        RECT 191.160 34.785 198.365 34.925 ;
        RECT 191.160 34.740 191.450 34.785 ;
        RECT 198.045 34.725 198.365 34.785 ;
        RECT 203.580 34.925 203.870 34.970 ;
        RECT 210.465 34.925 210.785 34.985 ;
        RECT 211.860 34.925 212.150 34.970 ;
        RECT 222.885 34.925 223.205 34.985 ;
        RECT 203.580 34.785 212.150 34.925 ;
        RECT 203.580 34.740 203.870 34.785 ;
        RECT 210.465 34.725 210.785 34.785 ;
        RECT 211.860 34.740 212.150 34.785 ;
        RECT 217.915 34.785 223.205 34.925 ;
        RECT 176.055 34.445 183.555 34.585 ;
        RECT 190.685 34.585 191.005 34.645 ;
        RECT 191.620 34.585 191.910 34.630 ;
        RECT 190.685 34.445 191.910 34.585 ;
        RECT 168.605 34.045 168.925 34.305 ;
        RECT 176.055 34.290 176.195 34.445 ;
        RECT 190.685 34.385 191.005 34.445 ;
        RECT 191.620 34.400 191.910 34.445 ;
        RECT 194.825 34.385 195.145 34.645 ;
        RECT 205.880 34.585 206.170 34.630 ;
        RECT 209.100 34.585 209.390 34.630 ;
        RECT 209.545 34.585 209.865 34.645 ;
        RECT 213.225 34.585 213.545 34.645 ;
        RECT 217.915 34.630 218.055 34.785 ;
        RECT 222.885 34.725 223.205 34.785 ;
        RECT 205.880 34.445 208.855 34.585 ;
        RECT 205.880 34.400 206.170 34.445 ;
        RECT 175.980 34.060 176.270 34.290 ;
        RECT 179.660 34.060 179.950 34.290 ;
        RECT 180.105 34.245 180.425 34.305 ;
        RECT 190.240 34.245 190.530 34.290 ;
        RECT 195.285 34.245 195.605 34.305 ;
        RECT 180.105 34.105 195.605 34.245 ;
        RECT 168.110 33.905 168.400 33.950 ;
        RECT 170.000 33.905 170.290 33.950 ;
        RECT 173.120 33.905 173.410 33.950 ;
        RECT 168.110 33.765 173.410 33.905 ;
        RECT 168.110 33.720 168.400 33.765 ;
        RECT 170.000 33.720 170.290 33.765 ;
        RECT 173.120 33.720 173.410 33.765 ;
        RECT 178.725 33.905 179.045 33.965 ;
        RECT 179.735 33.905 179.875 34.060 ;
        RECT 180.105 34.045 180.425 34.105 ;
        RECT 190.240 34.060 190.530 34.105 ;
        RECT 195.285 34.045 195.605 34.105 ;
        RECT 200.805 34.045 201.125 34.305 ;
        RECT 206.325 34.045 206.645 34.305 ;
        RECT 207.260 34.245 207.550 34.290 ;
        RECT 208.715 34.245 208.855 34.445 ;
        RECT 209.100 34.445 209.865 34.585 ;
        RECT 209.100 34.400 209.390 34.445 ;
        RECT 209.545 34.385 209.865 34.445 ;
        RECT 210.095 34.445 213.545 34.585 ;
        RECT 210.095 34.245 210.235 34.445 ;
        RECT 213.225 34.385 213.545 34.445 ;
        RECT 217.840 34.400 218.130 34.630 ;
        RECT 220.140 34.585 220.430 34.630 ;
        RECT 224.265 34.585 224.585 34.645 ;
        RECT 220.140 34.445 224.585 34.585 ;
        RECT 220.140 34.400 220.430 34.445 ;
        RECT 224.265 34.385 224.585 34.445 ;
        RECT 206.875 34.105 207.935 34.245 ;
        RECT 208.715 34.105 210.235 34.245 ;
        RECT 212.780 34.245 213.070 34.290 ;
        RECT 213.685 34.245 214.005 34.305 ;
        RECT 212.780 34.105 214.005 34.245 ;
        RECT 191.605 33.905 191.925 33.965 ;
        RECT 206.875 33.905 207.015 34.105 ;
        RECT 207.260 34.060 207.550 34.105 ;
        RECT 178.725 33.765 207.015 33.905 ;
        RECT 178.725 33.705 179.045 33.765 ;
        RECT 191.605 33.705 191.925 33.765 ;
        RECT 176.425 33.365 176.745 33.625 ;
        RECT 193.905 33.365 194.225 33.625 ;
        RECT 207.795 33.565 207.935 34.105 ;
        RECT 212.780 34.060 213.070 34.105 ;
        RECT 213.685 34.045 214.005 34.105 ;
        RECT 221.060 34.060 221.350 34.290 ;
        RECT 221.965 34.245 222.285 34.305 ;
        RECT 225.735 34.290 225.875 35.065 ;
        RECT 227.575 34.985 227.715 35.125 ;
        RECT 227.485 34.725 227.805 34.985 ;
        RECT 229.785 34.925 230.105 34.985 ;
        RECT 231.640 34.925 231.930 34.970 ;
        RECT 229.785 34.785 231.930 34.925 ;
        RECT 232.175 34.925 232.315 35.125 ;
        RECT 233.555 35.125 238.385 35.265 ;
        RECT 233.555 34.925 233.695 35.125 ;
        RECT 238.065 35.065 238.385 35.125 ;
        RECT 239.000 35.265 239.290 35.310 ;
        RECT 240.365 35.265 240.685 35.325 ;
        RECT 239.000 35.125 240.685 35.265 ;
        RECT 239.000 35.080 239.290 35.125 ;
        RECT 240.365 35.065 240.685 35.125 ;
        RECT 241.745 35.065 242.065 35.325 ;
        RECT 244.505 35.065 244.825 35.325 ;
        RECT 250.945 35.065 251.265 35.325 ;
        RECT 255.085 35.065 255.405 35.325 ;
        RECT 260.605 35.265 260.925 35.325 ;
        RECT 260.605 35.125 283.605 35.265 ;
        RECT 260.605 35.065 260.925 35.125 ;
        RECT 233.920 34.925 234.570 34.970 ;
        RECT 237.520 34.925 237.810 34.970 ;
        RECT 244.595 34.925 244.735 35.065 ;
        RECT 232.175 34.785 237.810 34.925 ;
        RECT 229.785 34.725 230.105 34.785 ;
        RECT 231.640 34.740 231.930 34.785 ;
        RECT 233.920 34.740 234.570 34.785 ;
        RECT 237.220 34.740 237.810 34.785 ;
        RECT 240.915 34.785 244.735 34.925 ;
        RECT 245.880 34.925 246.530 34.970 ;
        RECT 249.480 34.925 249.770 34.970 ;
        RECT 245.880 34.785 249.770 34.925 ;
        RECT 230.725 34.585 231.015 34.630 ;
        RECT 232.560 34.585 232.850 34.630 ;
        RECT 236.140 34.585 236.430 34.630 ;
        RECT 230.725 34.445 236.430 34.585 ;
        RECT 230.725 34.400 231.015 34.445 ;
        RECT 232.560 34.400 232.850 34.445 ;
        RECT 236.140 34.400 236.430 34.445 ;
        RECT 237.220 34.425 237.510 34.740 ;
        RECT 240.915 34.630 241.055 34.785 ;
        RECT 245.880 34.740 246.530 34.785 ;
        RECT 249.180 34.740 249.770 34.785 ;
        RECT 249.180 34.645 249.470 34.740 ;
        RECT 240.840 34.400 241.130 34.630 ;
        RECT 242.205 34.385 242.525 34.645 ;
        RECT 242.685 34.585 242.975 34.630 ;
        RECT 244.520 34.585 244.810 34.630 ;
        RECT 248.100 34.585 248.390 34.630 ;
        RECT 242.685 34.445 248.390 34.585 ;
        RECT 242.685 34.400 242.975 34.445 ;
        RECT 244.520 34.400 244.810 34.445 ;
        RECT 248.100 34.400 248.390 34.445 ;
        RECT 249.105 34.425 249.470 34.645 ;
        RECT 251.035 34.585 251.175 35.065 ;
        RECT 255.175 34.925 255.315 35.065 ;
        RECT 265.665 34.925 265.985 34.985 ;
        RECT 255.175 34.785 265.985 34.925 ;
        RECT 265.665 34.725 265.985 34.785 ;
        RECT 269.805 34.725 270.125 34.985 ;
        RECT 271.760 34.925 272.050 34.970 ;
        RECT 275.000 34.925 275.650 34.970 ;
        RECT 271.760 34.785 275.650 34.925 ;
        RECT 271.760 34.740 272.350 34.785 ;
        RECT 275.000 34.740 275.650 34.785 ;
        RECT 277.640 34.925 277.930 34.970 ;
        RECT 280.845 34.925 281.165 34.985 ;
        RECT 277.640 34.785 281.165 34.925 ;
        RECT 283.465 34.925 283.605 35.125 ;
        RECT 285.905 35.065 286.225 35.325 ;
        RECT 287.760 35.080 288.050 35.310 ;
        RECT 289.585 35.265 289.905 35.325 ;
        RECT 291.900 35.265 292.190 35.310 ;
        RECT 298.325 35.265 298.645 35.325 ;
        RECT 300.165 35.265 300.485 35.325 ;
        RECT 289.585 35.125 298.645 35.265 ;
        RECT 285.000 34.925 285.290 34.970 ;
        RECT 283.465 34.785 285.290 34.925 ;
        RECT 277.640 34.740 277.930 34.785 ;
        RECT 272.060 34.645 272.350 34.740 ;
        RECT 280.845 34.725 281.165 34.785 ;
        RECT 285.000 34.740 285.290 34.785 ;
        RECT 254.180 34.585 254.470 34.630 ;
        RECT 251.035 34.445 254.470 34.585 ;
        RECT 249.105 34.385 249.425 34.425 ;
        RECT 254.180 34.400 254.470 34.445 ;
        RECT 265.205 34.585 265.525 34.645 ;
        RECT 268.440 34.585 268.730 34.630 ;
        RECT 265.205 34.445 268.730 34.585 ;
        RECT 265.205 34.385 265.525 34.445 ;
        RECT 268.440 34.400 268.730 34.445 ;
        RECT 268.900 34.585 269.190 34.630 ;
        RECT 268.900 34.445 269.805 34.585 ;
        RECT 268.900 34.400 269.190 34.445 ;
        RECT 225.660 34.245 225.950 34.290 ;
        RECT 221.965 34.105 225.950 34.245 ;
        RECT 221.135 33.905 221.275 34.060 ;
        RECT 221.965 34.045 222.285 34.105 ;
        RECT 225.660 34.060 225.950 34.105 ;
        RECT 227.025 34.045 227.345 34.305 ;
        RECT 229.325 34.245 229.645 34.305 ;
        RECT 230.260 34.245 230.550 34.290 ;
        RECT 229.325 34.105 230.550 34.245 ;
        RECT 229.325 34.045 229.645 34.105 ;
        RECT 230.260 34.060 230.550 34.105 ;
        RECT 243.585 34.045 243.905 34.305 ;
        RECT 228.865 33.905 229.185 33.965 ;
        RECT 212.395 33.765 229.185 33.905 ;
        RECT 212.395 33.565 212.535 33.765 ;
        RECT 228.865 33.705 229.185 33.765 ;
        RECT 231.130 33.905 231.420 33.950 ;
        RECT 233.020 33.905 233.310 33.950 ;
        RECT 236.140 33.905 236.430 33.950 ;
        RECT 231.130 33.765 236.430 33.905 ;
        RECT 231.130 33.720 231.420 33.765 ;
        RECT 233.020 33.720 233.310 33.765 ;
        RECT 236.140 33.720 236.430 33.765 ;
        RECT 243.090 33.905 243.380 33.950 ;
        RECT 244.980 33.905 245.270 33.950 ;
        RECT 248.100 33.905 248.390 33.950 ;
        RECT 243.090 33.765 248.390 33.905 ;
        RECT 268.515 33.905 268.655 34.400 ;
        RECT 269.665 34.245 269.805 34.445 ;
        RECT 272.060 34.425 272.425 34.645 ;
        RECT 272.105 34.385 272.425 34.425 ;
        RECT 273.140 34.585 273.430 34.630 ;
        RECT 276.720 34.585 277.010 34.630 ;
        RECT 278.555 34.585 278.845 34.630 ;
        RECT 273.140 34.445 278.845 34.585 ;
        RECT 273.140 34.400 273.430 34.445 ;
        RECT 276.720 34.400 277.010 34.445 ;
        RECT 278.555 34.400 278.845 34.445 ;
        RECT 279.005 34.585 279.325 34.645 ;
        RECT 285.995 34.585 286.135 35.065 ;
        RECT 286.840 34.925 287.130 34.970 ;
        RECT 287.835 34.925 287.975 35.080 ;
        RECT 289.585 35.065 289.905 35.125 ;
        RECT 291.900 35.080 292.190 35.125 ;
        RECT 298.325 35.065 298.645 35.125 ;
        RECT 298.875 35.125 300.485 35.265 ;
        RECT 296.945 34.925 297.265 34.985 ;
        RECT 298.875 34.970 299.015 35.125 ;
        RECT 300.165 35.065 300.485 35.125 ;
        RECT 303.385 35.265 303.705 35.325 ;
        RECT 303.385 35.125 307.295 35.265 ;
        RECT 303.385 35.065 303.705 35.125 ;
        RECT 297.880 34.925 298.170 34.970 ;
        RECT 286.840 34.785 287.975 34.925 ;
        RECT 290.595 34.785 296.255 34.925 ;
        RECT 286.840 34.740 287.130 34.785 ;
        RECT 290.595 34.630 290.735 34.785 ;
        RECT 296.115 34.630 296.255 34.785 ;
        RECT 296.945 34.785 298.170 34.925 ;
        RECT 296.945 34.725 297.265 34.785 ;
        RECT 297.880 34.740 298.170 34.785 ;
        RECT 298.800 34.740 299.090 34.970 ;
        RECT 301.200 34.925 301.490 34.970 ;
        RECT 302.005 34.925 302.325 34.985 ;
        RECT 307.155 34.970 307.295 35.125 ;
        RECT 304.440 34.925 305.090 34.970 ;
        RECT 301.200 34.785 305.090 34.925 ;
        RECT 301.200 34.740 301.790 34.785 ;
        RECT 290.520 34.585 290.810 34.630 ;
        RECT 279.005 34.445 283.605 34.585 ;
        RECT 285.995 34.445 290.810 34.585 ;
        RECT 279.005 34.385 279.325 34.445 ;
        RECT 270.280 34.245 270.570 34.290 ;
        RECT 279.925 34.245 280.245 34.305 ;
        RECT 269.665 34.105 280.245 34.245 ;
        RECT 270.280 34.060 270.570 34.105 ;
        RECT 279.925 34.045 280.245 34.105 ;
        RECT 273.140 33.905 273.430 33.950 ;
        RECT 276.260 33.905 276.550 33.950 ;
        RECT 278.150 33.905 278.440 33.950 ;
        RECT 268.515 33.765 272.795 33.905 ;
        RECT 243.090 33.720 243.380 33.765 ;
        RECT 244.980 33.720 245.270 33.765 ;
        RECT 248.100 33.720 248.390 33.765 ;
        RECT 207.795 33.425 212.535 33.565 ;
        RECT 213.225 33.565 213.545 33.625 ;
        RECT 214.620 33.565 214.910 33.610 ;
        RECT 213.225 33.425 214.910 33.565 ;
        RECT 213.225 33.365 213.545 33.425 ;
        RECT 214.620 33.380 214.910 33.425 ;
        RECT 215.985 33.565 216.305 33.625 ;
        RECT 218.300 33.565 218.590 33.610 ;
        RECT 215.985 33.425 218.590 33.565 ;
        RECT 215.985 33.365 216.305 33.425 ;
        RECT 218.300 33.380 218.590 33.425 ;
        RECT 224.265 33.565 224.585 33.625 ;
        RECT 229.800 33.565 230.090 33.610 ;
        RECT 233.925 33.565 234.245 33.625 ;
        RECT 224.265 33.425 234.245 33.565 ;
        RECT 224.265 33.365 224.585 33.425 ;
        RECT 229.800 33.380 230.090 33.425 ;
        RECT 233.925 33.365 234.245 33.425 ;
        RECT 251.405 33.365 251.725 33.625 ;
        RECT 269.345 33.365 269.665 33.625 ;
        RECT 272.655 33.565 272.795 33.765 ;
        RECT 273.140 33.765 278.440 33.905 ;
        RECT 283.465 33.905 283.605 34.445 ;
        RECT 290.520 34.400 290.810 34.445 ;
        RECT 292.360 34.400 292.650 34.630 ;
        RECT 296.040 34.400 296.330 34.630 ;
        RECT 301.500 34.425 301.790 34.740 ;
        RECT 302.005 34.725 302.325 34.785 ;
        RECT 304.440 34.740 305.090 34.785 ;
        RECT 307.080 34.740 307.370 34.970 ;
        RECT 302.580 34.585 302.870 34.630 ;
        RECT 306.160 34.585 306.450 34.630 ;
        RECT 307.995 34.585 308.285 34.630 ;
        RECT 302.580 34.445 308.285 34.585 ;
        RECT 302.580 34.400 302.870 34.445 ;
        RECT 306.160 34.400 306.450 34.445 ;
        RECT 307.995 34.400 308.285 34.445 ;
        RECT 308.460 34.585 308.750 34.630 ;
        RECT 308.905 34.585 309.225 34.645 ;
        RECT 308.460 34.445 309.225 34.585 ;
        RECT 308.460 34.400 308.750 34.445 ;
        RECT 285.445 34.245 285.765 34.305 ;
        RECT 289.140 34.245 289.430 34.290 ;
        RECT 292.435 34.245 292.575 34.400 ;
        RECT 285.445 34.105 292.575 34.245 ;
        RECT 296.115 34.245 296.255 34.400 ;
        RECT 308.905 34.385 309.225 34.445 ;
        RECT 298.785 34.245 299.105 34.305 ;
        RECT 299.720 34.245 300.010 34.290 ;
        RECT 296.115 34.105 300.010 34.245 ;
        RECT 285.445 34.045 285.765 34.105 ;
        RECT 289.140 34.060 289.430 34.105 ;
        RECT 298.785 34.045 299.105 34.105 ;
        RECT 299.720 34.060 300.010 34.105 ;
        RECT 286.365 33.905 286.685 33.965 ;
        RECT 288.665 33.905 288.985 33.965 ;
        RECT 290.965 33.905 291.285 33.965 ;
        RECT 283.465 33.765 291.285 33.905 ;
        RECT 273.140 33.720 273.430 33.765 ;
        RECT 276.260 33.720 276.550 33.765 ;
        RECT 278.150 33.720 278.440 33.765 ;
        RECT 286.365 33.705 286.685 33.765 ;
        RECT 288.665 33.705 288.985 33.765 ;
        RECT 290.965 33.705 291.285 33.765 ;
        RECT 302.580 33.905 302.870 33.950 ;
        RECT 305.700 33.905 305.990 33.950 ;
        RECT 307.590 33.905 307.880 33.950 ;
        RECT 302.580 33.765 307.880 33.905 ;
        RECT 302.580 33.720 302.870 33.765 ;
        RECT 305.700 33.720 305.990 33.765 ;
        RECT 307.590 33.720 307.880 33.765 ;
        RECT 275.785 33.565 276.105 33.625 ;
        RECT 272.655 33.425 276.105 33.565 ;
        RECT 275.785 33.365 276.105 33.425 ;
        RECT 282.700 33.565 282.990 33.610 ;
        RECT 284.065 33.565 284.385 33.625 ;
        RECT 282.700 33.425 284.385 33.565 ;
        RECT 282.700 33.380 282.990 33.425 ;
        RECT 284.065 33.365 284.385 33.425 ;
        RECT 289.125 33.365 289.445 33.625 ;
        RECT 293.280 33.565 293.570 33.610 ;
        RECT 293.725 33.565 294.045 33.625 ;
        RECT 293.280 33.425 294.045 33.565 ;
        RECT 293.280 33.380 293.570 33.425 ;
        RECT 293.725 33.365 294.045 33.425 ;
        RECT 162.095 32.745 311.135 33.225 ;
        RECT 167.225 32.345 167.545 32.605 ;
        RECT 168.605 32.545 168.925 32.605 ;
        RECT 170.920 32.545 171.210 32.590 ;
        RECT 168.605 32.405 171.210 32.545 ;
        RECT 168.605 32.345 168.925 32.405 ;
        RECT 170.920 32.360 171.210 32.405 ;
        RECT 178.725 32.345 179.045 32.605 ;
        RECT 190.175 32.545 190.465 32.590 ;
        RECT 193.905 32.545 194.225 32.605 ;
        RECT 190.175 32.405 194.225 32.545 ;
        RECT 190.175 32.360 190.465 32.405 ;
        RECT 193.905 32.345 194.225 32.405 ;
        RECT 197.585 32.345 197.905 32.605 ;
        RECT 200.805 32.545 201.125 32.605 ;
        RECT 205.420 32.545 205.710 32.590 ;
        RECT 200.805 32.405 205.710 32.545 ;
        RECT 200.805 32.345 201.125 32.405 ;
        RECT 205.420 32.360 205.710 32.405 ;
        RECT 212.870 32.545 213.160 32.590 ;
        RECT 214.620 32.545 214.910 32.590 ;
        RECT 212.870 32.405 214.910 32.545 ;
        RECT 212.870 32.360 213.160 32.405 ;
        RECT 214.620 32.360 214.910 32.405 ;
        RECT 218.695 32.545 218.985 32.590 ;
        RECT 220.585 32.545 220.905 32.605 ;
        RECT 218.695 32.405 220.905 32.545 ;
        RECT 218.695 32.360 218.985 32.405 ;
        RECT 220.585 32.345 220.905 32.405 ;
        RECT 227.025 32.345 227.345 32.605 ;
        RECT 243.585 32.545 243.905 32.605 ;
        RECT 244.060 32.545 244.350 32.590 ;
        RECT 228.955 32.405 243.355 32.545 ;
        RECT 167.315 32.205 167.455 32.345 ;
        RECT 169.080 32.205 169.370 32.250 ;
        RECT 167.315 32.065 169.370 32.205 ;
        RECT 169.080 32.020 169.370 32.065 ;
        RECT 176.425 31.865 176.745 31.925 ;
        RECT 178.815 31.910 178.955 32.345 ;
        RECT 228.955 32.265 229.095 32.405 ;
        RECT 182.520 32.205 182.810 32.250 ;
        RECT 185.640 32.205 185.930 32.250 ;
        RECT 187.530 32.205 187.820 32.250 ;
        RECT 182.520 32.065 187.820 32.205 ;
        RECT 182.520 32.020 182.810 32.065 ;
        RECT 185.640 32.020 185.930 32.065 ;
        RECT 187.530 32.020 187.820 32.065 ;
        RECT 189.730 32.205 190.020 32.250 ;
        RECT 191.620 32.205 191.910 32.250 ;
        RECT 194.740 32.205 195.030 32.250 ;
        RECT 207.705 32.205 208.025 32.265 ;
        RECT 189.730 32.065 195.030 32.205 ;
        RECT 189.730 32.020 190.020 32.065 ;
        RECT 191.620 32.020 191.910 32.065 ;
        RECT 194.740 32.020 195.030 32.065 ;
        RECT 204.115 32.065 208.025 32.205 ;
        RECT 170.075 31.725 176.745 31.865 ;
        RECT 170.075 31.570 170.215 31.725 ;
        RECT 176.425 31.665 176.745 31.725 ;
        RECT 178.740 31.680 179.030 31.910 ;
        RECT 187.005 31.665 187.325 31.925 ;
        RECT 188.400 31.865 188.690 31.910 ;
        RECT 188.860 31.865 189.150 31.910 ;
        RECT 190.225 31.865 190.545 31.925 ;
        RECT 188.400 31.725 190.545 31.865 ;
        RECT 188.400 31.680 188.690 31.725 ;
        RECT 188.860 31.680 189.150 31.725 ;
        RECT 190.225 31.665 190.545 31.725 ;
        RECT 192.985 31.865 193.305 31.925 ;
        RECT 204.115 31.865 204.255 32.065 ;
        RECT 207.705 32.005 208.025 32.065 ;
        RECT 208.280 32.205 208.570 32.250 ;
        RECT 211.400 32.205 211.690 32.250 ;
        RECT 213.290 32.205 213.580 32.250 ;
        RECT 208.280 32.065 213.580 32.205 ;
        RECT 208.280 32.020 208.570 32.065 ;
        RECT 211.400 32.020 211.690 32.065 ;
        RECT 213.290 32.020 213.580 32.065 ;
        RECT 218.250 32.205 218.540 32.250 ;
        RECT 220.140 32.205 220.430 32.250 ;
        RECT 223.260 32.205 223.550 32.250 ;
        RECT 218.250 32.065 223.550 32.205 ;
        RECT 218.250 32.020 218.540 32.065 ;
        RECT 220.140 32.020 220.430 32.065 ;
        RECT 223.260 32.020 223.550 32.065 ;
        RECT 228.865 32.005 229.185 32.265 ;
        RECT 229.900 32.205 230.190 32.250 ;
        RECT 233.020 32.205 233.310 32.250 ;
        RECT 234.910 32.205 235.200 32.250 ;
        RECT 229.900 32.065 235.200 32.205 ;
        RECT 243.215 32.205 243.355 32.405 ;
        RECT 243.585 32.405 244.350 32.545 ;
        RECT 243.585 32.345 243.905 32.405 ;
        RECT 244.060 32.360 244.350 32.405 ;
        RECT 265.205 32.345 265.525 32.605 ;
        RECT 272.670 32.545 272.960 32.590 ;
        RECT 276.705 32.545 277.025 32.605 ;
        RECT 272.670 32.405 277.025 32.545 ;
        RECT 272.670 32.360 272.960 32.405 ;
        RECT 276.705 32.345 277.025 32.405 ;
        RECT 279.555 32.405 284.295 32.545 ;
        RECT 260.605 32.205 260.925 32.265 ;
        RECT 243.215 32.065 260.925 32.205 ;
        RECT 229.900 32.020 230.190 32.065 ;
        RECT 233.020 32.020 233.310 32.065 ;
        RECT 234.910 32.020 235.200 32.065 ;
        RECT 216.445 31.865 216.765 31.925 ;
        RECT 217.380 31.865 217.670 31.910 ;
        RECT 229.325 31.865 229.645 31.925 ;
        RECT 248.275 31.910 248.415 32.065 ;
        RECT 260.605 32.005 260.925 32.065 ;
        RECT 268.080 32.205 268.370 32.250 ;
        RECT 271.200 32.205 271.490 32.250 ;
        RECT 273.090 32.205 273.380 32.250 ;
        RECT 268.080 32.065 273.380 32.205 ;
        RECT 268.080 32.020 268.370 32.065 ;
        RECT 271.200 32.020 271.490 32.065 ;
        RECT 273.090 32.020 273.380 32.065 ;
        RECT 235.780 31.865 236.070 31.910 ;
        RECT 192.985 31.725 204.255 31.865 ;
        RECT 204.575 31.725 215.295 31.865 ;
        RECT 192.985 31.665 193.305 31.725 ;
        RECT 170.000 31.340 170.290 31.570 ;
        RECT 171.840 31.525 172.130 31.570 ;
        RECT 171.840 31.385 173.205 31.525 ;
        RECT 171.840 31.340 172.130 31.385 ;
        RECT 173.065 30.845 173.205 31.385 ;
        RECT 177.820 31.185 178.110 31.230 ;
        RECT 178.265 31.185 178.585 31.245 ;
        RECT 181.440 31.230 181.730 31.545 ;
        RECT 182.520 31.525 182.810 31.570 ;
        RECT 186.100 31.525 186.390 31.570 ;
        RECT 187.935 31.525 188.225 31.570 ;
        RECT 182.520 31.385 188.225 31.525 ;
        RECT 182.520 31.340 182.810 31.385 ;
        RECT 186.100 31.340 186.390 31.385 ;
        RECT 187.935 31.340 188.225 31.385 ;
        RECT 189.325 31.525 189.615 31.570 ;
        RECT 191.160 31.525 191.450 31.570 ;
        RECT 194.740 31.525 195.030 31.570 ;
        RECT 189.325 31.385 195.030 31.525 ;
        RECT 189.325 31.340 189.615 31.385 ;
        RECT 191.160 31.340 191.450 31.385 ;
        RECT 194.740 31.340 195.030 31.385 ;
        RECT 195.820 31.230 196.110 31.545 ;
        RECT 177.820 31.045 178.585 31.185 ;
        RECT 177.820 31.000 178.110 31.045 ;
        RECT 178.265 30.985 178.585 31.045 ;
        RECT 181.140 31.185 181.730 31.230 ;
        RECT 184.380 31.185 185.030 31.230 ;
        RECT 192.520 31.185 193.170 31.230 ;
        RECT 195.820 31.185 196.410 31.230 ;
        RECT 196.665 31.185 196.985 31.245 ;
        RECT 204.575 31.230 204.715 31.725 ;
        RECT 207.200 31.230 207.490 31.545 ;
        RECT 208.280 31.525 208.570 31.570 ;
        RECT 211.860 31.525 212.150 31.570 ;
        RECT 213.695 31.525 213.985 31.570 ;
        RECT 208.280 31.385 213.985 31.525 ;
        RECT 208.280 31.340 208.570 31.385 ;
        RECT 211.860 31.340 212.150 31.385 ;
        RECT 213.695 31.340 213.985 31.385 ;
        RECT 214.160 31.340 214.450 31.570 ;
        RECT 181.140 31.045 191.375 31.185 ;
        RECT 181.140 31.000 181.430 31.045 ;
        RECT 184.380 31.000 185.030 31.045 ;
        RECT 175.520 30.845 175.810 30.890 ;
        RECT 173.065 30.705 175.810 30.845 ;
        RECT 175.520 30.660 175.810 30.705 ;
        RECT 177.360 30.845 177.650 30.890 ;
        RECT 179.660 30.845 179.950 30.890 ;
        RECT 190.685 30.845 191.005 30.905 ;
        RECT 177.360 30.705 191.005 30.845 ;
        RECT 191.235 30.845 191.375 31.045 ;
        RECT 192.520 31.045 203.795 31.185 ;
        RECT 192.520 31.000 193.170 31.045 ;
        RECT 196.120 31.000 196.410 31.045 ;
        RECT 196.665 30.985 196.985 31.045 ;
        RECT 196.755 30.845 196.895 30.985 ;
        RECT 191.235 30.705 196.895 30.845 ;
        RECT 200.345 30.845 200.665 30.905 ;
        RECT 203.120 30.845 203.410 30.890 ;
        RECT 200.345 30.705 203.410 30.845 ;
        RECT 203.655 30.845 203.795 31.045 ;
        RECT 204.500 31.000 204.790 31.230 ;
        RECT 206.900 31.185 207.490 31.230 ;
        RECT 210.140 31.185 210.790 31.230 ;
        RECT 212.305 31.185 212.625 31.245 ;
        RECT 206.900 31.045 212.625 31.185 ;
        RECT 206.900 31.000 207.190 31.045 ;
        RECT 210.140 31.000 210.790 31.045 ;
        RECT 212.305 30.985 212.625 31.045 ;
        RECT 214.235 30.905 214.375 31.340 ;
        RECT 215.155 31.185 215.295 31.725 ;
        RECT 216.445 31.725 236.070 31.865 ;
        RECT 216.445 31.665 216.765 31.725 ;
        RECT 217.380 31.680 217.670 31.725 ;
        RECT 229.325 31.665 229.645 31.725 ;
        RECT 235.780 31.680 236.070 31.725 ;
        RECT 248.200 31.680 248.490 31.910 ;
        RECT 251.405 31.665 251.725 31.925 ;
        RECT 215.525 31.325 215.845 31.585 ;
        RECT 215.985 31.525 216.305 31.585 ;
        RECT 216.920 31.525 217.210 31.570 ;
        RECT 215.985 31.385 217.210 31.525 ;
        RECT 215.985 31.325 216.305 31.385 ;
        RECT 216.920 31.340 217.210 31.385 ;
        RECT 217.845 31.525 218.135 31.570 ;
        RECT 219.680 31.525 219.970 31.570 ;
        RECT 223.260 31.525 223.550 31.570 ;
        RECT 217.845 31.385 223.550 31.525 ;
        RECT 217.845 31.340 218.135 31.385 ;
        RECT 219.680 31.340 219.970 31.385 ;
        RECT 223.260 31.340 223.550 31.385 ;
        RECT 224.340 31.230 224.630 31.545 ;
        RECT 221.040 31.185 221.690 31.230 ;
        RECT 224.340 31.185 224.930 31.230 ;
        RECT 227.485 31.185 227.805 31.245 ;
        RECT 228.820 31.230 229.110 31.545 ;
        RECT 229.900 31.525 230.190 31.570 ;
        RECT 233.480 31.525 233.770 31.570 ;
        RECT 235.315 31.525 235.605 31.570 ;
        RECT 229.900 31.385 235.605 31.525 ;
        RECT 229.900 31.340 230.190 31.385 ;
        RECT 233.480 31.340 233.770 31.385 ;
        RECT 235.315 31.340 235.605 31.385 ;
        RECT 236.225 31.325 236.545 31.585 ;
        RECT 238.065 31.325 238.385 31.585 ;
        RECT 244.980 31.525 245.270 31.570 ;
        RECT 247.740 31.525 248.030 31.570 ;
        RECT 251.495 31.525 251.635 31.665 ;
        RECT 244.980 31.385 245.655 31.525 ;
        RECT 244.980 31.340 245.270 31.385 ;
        RECT 215.155 31.045 224.930 31.185 ;
        RECT 205.405 30.845 205.725 30.905 ;
        RECT 203.655 30.705 205.725 30.845 ;
        RECT 177.360 30.660 177.650 30.705 ;
        RECT 179.660 30.660 179.950 30.705 ;
        RECT 190.685 30.645 191.005 30.705 ;
        RECT 200.345 30.645 200.665 30.705 ;
        RECT 203.120 30.660 203.410 30.705 ;
        RECT 205.405 30.645 205.725 30.705 ;
        RECT 205.865 30.845 206.185 30.905 ;
        RECT 214.145 30.845 214.465 30.905 ;
        RECT 205.865 30.705 214.465 30.845 ;
        RECT 205.865 30.645 206.185 30.705 ;
        RECT 214.145 30.645 214.465 30.705 ;
        RECT 215.985 30.645 216.305 30.905 ;
        RECT 220.675 30.845 220.815 31.045 ;
        RECT 221.040 31.000 221.690 31.045 ;
        RECT 224.640 31.000 224.930 31.045 ;
        RECT 225.735 31.045 227.805 31.185 ;
        RECT 225.735 30.845 225.875 31.045 ;
        RECT 227.485 30.985 227.805 31.045 ;
        RECT 228.520 31.185 229.110 31.230 ;
        RECT 231.760 31.185 232.410 31.230 ;
        RECT 228.520 31.045 233.695 31.185 ;
        RECT 228.520 31.000 228.810 31.045 ;
        RECT 231.760 31.000 232.410 31.045 ;
        RECT 233.555 30.905 233.695 31.045 ;
        RECT 234.385 30.985 234.705 31.245 ;
        RECT 220.675 30.705 225.875 30.845 ;
        RECT 226.120 30.845 226.410 30.890 ;
        RECT 230.245 30.845 230.565 30.905 ;
        RECT 226.120 30.705 230.565 30.845 ;
        RECT 226.120 30.660 226.410 30.705 ;
        RECT 230.245 30.645 230.565 30.705 ;
        RECT 233.465 30.645 233.785 30.905 ;
        RECT 245.515 30.890 245.655 31.385 ;
        RECT 247.740 31.385 251.635 31.525 ;
        RECT 247.740 31.340 248.030 31.385 ;
        RECT 253.705 31.325 254.025 31.585 ;
        RECT 260.695 31.570 260.835 32.005 ;
        RECT 279.555 31.925 279.695 32.405 ;
        RECT 279.925 32.205 280.245 32.265 ;
        RECT 283.605 32.205 283.925 32.265 ;
        RECT 279.925 32.065 282.915 32.205 ;
        RECT 279.925 32.005 280.245 32.065 ;
        RECT 273.960 31.865 274.250 31.910 ;
        RECT 279.005 31.865 279.325 31.925 ;
        RECT 273.960 31.725 279.325 31.865 ;
        RECT 273.960 31.680 274.250 31.725 ;
        RECT 279.005 31.665 279.325 31.725 ;
        RECT 279.465 31.865 279.785 31.925 ;
        RECT 281.320 31.865 281.610 31.910 ;
        RECT 279.465 31.725 281.610 31.865 ;
        RECT 279.465 31.665 279.785 31.725 ;
        RECT 281.320 31.680 281.610 31.725 ;
        RECT 282.225 31.665 282.545 31.925 ;
        RECT 260.620 31.340 260.910 31.570 ;
        RECT 265.665 31.525 265.985 31.585 ;
        RECT 267.000 31.525 267.290 31.545 ;
        RECT 265.665 31.385 267.290 31.525 ;
        RECT 265.665 31.325 265.985 31.385 ;
        RECT 247.280 31.185 247.570 31.230 ;
        RECT 253.795 31.185 253.935 31.325 ;
        RECT 267.000 31.230 267.290 31.385 ;
        RECT 268.080 31.525 268.370 31.570 ;
        RECT 271.660 31.525 271.950 31.570 ;
        RECT 273.495 31.525 273.785 31.570 ;
        RECT 268.080 31.385 273.785 31.525 ;
        RECT 268.080 31.340 268.370 31.385 ;
        RECT 271.660 31.340 271.950 31.385 ;
        RECT 273.495 31.340 273.785 31.385 ;
        RECT 274.880 31.525 275.170 31.570 ;
        RECT 276.245 31.525 276.565 31.585 ;
        RECT 274.880 31.385 276.565 31.525 ;
        RECT 274.880 31.340 275.170 31.385 ;
        RECT 276.245 31.325 276.565 31.385 ;
        RECT 280.860 31.525 281.150 31.570 ;
        RECT 282.315 31.525 282.455 31.665 ;
        RECT 282.775 31.570 282.915 32.065 ;
        RECT 283.465 32.005 283.925 32.205 ;
        RECT 283.465 31.865 283.605 32.005 ;
        RECT 283.235 31.725 283.605 31.865 ;
        RECT 280.860 31.385 282.455 31.525 ;
        RECT 280.860 31.340 281.150 31.385 ;
        RECT 282.700 31.340 282.990 31.570 ;
        RECT 247.280 31.045 253.935 31.185 ;
        RECT 257.860 31.185 258.150 31.230 ;
        RECT 258.780 31.185 259.070 31.230 ;
        RECT 257.860 31.045 259.070 31.185 ;
        RECT 247.280 31.000 247.570 31.045 ;
        RECT 257.860 31.000 258.150 31.045 ;
        RECT 258.780 31.000 259.070 31.045 ;
        RECT 259.700 31.000 259.990 31.230 ;
        RECT 266.700 31.185 267.290 31.230 ;
        RECT 269.940 31.185 270.590 31.230 ;
        RECT 266.700 31.045 270.590 31.185 ;
        RECT 266.700 31.000 266.990 31.045 ;
        RECT 269.940 31.000 270.590 31.045 ;
        RECT 272.565 31.185 272.885 31.245 ;
        RECT 279.005 31.185 279.325 31.245 ;
        RECT 280.400 31.185 280.690 31.230 ;
        RECT 283.235 31.185 283.375 31.725 ;
        RECT 283.620 31.525 283.910 31.570 ;
        RECT 284.155 31.525 284.295 32.405 ;
        RECT 285.445 32.345 285.765 32.605 ;
        RECT 292.910 32.545 293.200 32.590 ;
        RECT 293.725 32.545 294.045 32.605 ;
        RECT 292.910 32.405 294.045 32.545 ;
        RECT 292.910 32.360 293.200 32.405 ;
        RECT 293.725 32.345 294.045 32.405 ;
        RECT 294.645 32.345 294.965 32.605 ;
        RECT 288.320 32.205 288.610 32.250 ;
        RECT 291.440 32.205 291.730 32.250 ;
        RECT 293.330 32.205 293.620 32.250 ;
        RECT 288.320 32.065 293.620 32.205 ;
        RECT 288.320 32.020 288.610 32.065 ;
        RECT 291.440 32.020 291.730 32.065 ;
        RECT 293.330 32.020 293.620 32.065 ;
        RECT 297.520 32.205 297.810 32.250 ;
        RECT 300.640 32.205 300.930 32.250 ;
        RECT 302.530 32.205 302.820 32.250 ;
        RECT 297.520 32.065 302.820 32.205 ;
        RECT 297.520 32.020 297.810 32.065 ;
        RECT 300.640 32.020 300.930 32.065 ;
        RECT 302.530 32.020 302.820 32.065 ;
        RECT 290.965 31.865 291.285 31.925 ;
        RECT 294.200 31.865 294.490 31.910 ;
        RECT 303.400 31.865 303.690 31.910 ;
        RECT 308.445 31.865 308.765 31.925 ;
        RECT 290.965 31.725 308.765 31.865 ;
        RECT 290.965 31.665 291.285 31.725 ;
        RECT 294.200 31.680 294.490 31.725 ;
        RECT 303.400 31.680 303.690 31.725 ;
        RECT 308.445 31.665 308.765 31.725 ;
        RECT 287.285 31.545 287.605 31.585 ;
        RECT 283.620 31.385 284.295 31.525 ;
        RECT 283.620 31.340 283.910 31.385 ;
        RECT 287.240 31.325 287.605 31.545 ;
        RECT 288.320 31.525 288.610 31.570 ;
        RECT 291.900 31.525 292.190 31.570 ;
        RECT 293.735 31.525 294.025 31.570 ;
        RECT 288.320 31.385 294.025 31.525 ;
        RECT 288.320 31.340 288.610 31.385 ;
        RECT 291.900 31.340 292.190 31.385 ;
        RECT 293.735 31.340 294.025 31.385 ;
        RECT 287.240 31.230 287.530 31.325 ;
        RECT 296.440 31.230 296.730 31.545 ;
        RECT 297.520 31.525 297.810 31.570 ;
        RECT 301.100 31.525 301.390 31.570 ;
        RECT 302.935 31.525 303.225 31.570 ;
        RECT 297.520 31.385 303.225 31.525 ;
        RECT 297.520 31.340 297.810 31.385 ;
        RECT 301.100 31.340 301.390 31.385 ;
        RECT 302.935 31.340 303.225 31.385 ;
        RECT 303.845 31.525 304.165 31.585 ;
        RECT 307.080 31.525 307.370 31.570 ;
        RECT 303.845 31.385 307.370 31.525 ;
        RECT 303.845 31.325 304.165 31.385 ;
        RECT 307.080 31.340 307.370 31.385 ;
        RECT 272.565 31.045 278.775 31.185 ;
        RECT 245.440 30.660 245.730 30.890 ;
        RECT 247.725 30.845 248.045 30.905 ;
        RECT 256.480 30.845 256.770 30.890 ;
        RECT 247.725 30.705 256.770 30.845 ;
        RECT 259.775 30.845 259.915 31.000 ;
        RECT 272.565 30.985 272.885 31.045 ;
        RECT 269.345 30.845 269.665 30.905 ;
        RECT 259.775 30.705 269.665 30.845 ;
        RECT 247.725 30.645 248.045 30.705 ;
        RECT 256.480 30.660 256.770 30.705 ;
        RECT 269.345 30.645 269.665 30.705 ;
        RECT 277.625 30.645 277.945 30.905 ;
        RECT 278.635 30.890 278.775 31.045 ;
        RECT 279.005 31.045 283.375 31.185 ;
        RECT 286.940 31.185 287.530 31.230 ;
        RECT 290.180 31.185 290.830 31.230 ;
        RECT 286.940 31.045 290.830 31.185 ;
        RECT 279.005 30.985 279.325 31.045 ;
        RECT 280.400 31.000 280.690 31.045 ;
        RECT 282.315 30.905 282.455 31.045 ;
        RECT 286.940 31.000 287.230 31.045 ;
        RECT 290.180 31.000 290.830 31.045 ;
        RECT 296.140 31.185 296.730 31.230 ;
        RECT 299.380 31.185 300.030 31.230 ;
        RECT 302.020 31.185 302.310 31.230 ;
        RECT 304.320 31.185 304.610 31.230 ;
        RECT 296.140 31.045 301.315 31.185 ;
        RECT 296.140 31.000 296.430 31.045 ;
        RECT 299.380 31.000 300.030 31.045 ;
        RECT 278.560 30.660 278.850 30.890 ;
        RECT 282.225 30.645 282.545 30.905 ;
        RECT 282.685 30.645 283.005 30.905 ;
        RECT 301.175 30.845 301.315 31.045 ;
        RECT 302.020 31.045 304.610 31.185 ;
        RECT 302.020 31.000 302.310 31.045 ;
        RECT 304.320 31.000 304.610 31.045 ;
        RECT 305.225 30.985 305.545 31.245 ;
        RECT 305.315 30.845 305.455 30.985 ;
        RECT 301.175 30.705 305.455 30.845 ;
        RECT 162.095 30.025 311.935 30.505 ;
        RECT 187.005 29.625 187.325 29.885 ;
        RECT 192.985 29.825 193.305 29.885 ;
        RECT 189.855 29.685 193.305 29.825 ;
        RECT 189.855 29.485 189.995 29.685 ;
        RECT 192.985 29.625 193.305 29.685 ;
        RECT 193.460 29.825 193.750 29.870 ;
        RECT 194.365 29.825 194.685 29.885 ;
        RECT 193.460 29.685 194.685 29.825 ;
        RECT 193.460 29.640 193.750 29.685 ;
        RECT 194.365 29.625 194.685 29.685 ;
        RECT 194.825 29.825 195.145 29.885 ;
        RECT 195.760 29.825 196.050 29.870 ;
        RECT 194.825 29.685 196.050 29.825 ;
        RECT 194.825 29.625 195.145 29.685 ;
        RECT 195.760 29.640 196.050 29.685 ;
        RECT 210.465 29.625 210.785 29.885 ;
        RECT 212.780 29.825 213.070 29.870 ;
        RECT 215.065 29.825 215.385 29.885 ;
        RECT 215.985 29.825 216.305 29.885 ;
        RECT 212.780 29.685 215.385 29.825 ;
        RECT 212.780 29.640 213.070 29.685 ;
        RECT 215.065 29.625 215.385 29.685 ;
        RECT 215.615 29.685 216.305 29.825 ;
        RECT 165.015 29.345 189.995 29.485 ;
        RECT 190.225 29.485 190.545 29.545 ;
        RECT 200.360 29.485 200.650 29.530 ;
        RECT 201.725 29.485 202.045 29.545 ;
        RECT 190.225 29.345 199.195 29.485 ;
        RECT 165.015 29.190 165.155 29.345 ;
        RECT 190.225 29.285 190.545 29.345 ;
        RECT 164.940 28.960 165.230 29.190 ;
        RECT 186.085 28.945 186.405 29.205 ;
        RECT 199.055 29.190 199.195 29.345 ;
        RECT 200.360 29.345 202.045 29.485 ;
        RECT 200.360 29.300 200.650 29.345 ;
        RECT 201.725 29.285 202.045 29.345 ;
        RECT 202.640 29.485 203.290 29.530 ;
        RECT 206.240 29.485 206.530 29.530 ;
        RECT 202.640 29.345 206.530 29.485 ;
        RECT 202.640 29.300 203.290 29.345 ;
        RECT 205.940 29.300 206.530 29.345 ;
        RECT 210.940 29.485 211.230 29.530 ;
        RECT 213.225 29.485 213.545 29.545 ;
        RECT 215.615 29.530 215.755 29.685 ;
        RECT 215.985 29.625 216.305 29.685 ;
        RECT 222.885 29.625 223.205 29.885 ;
        RECT 231.640 29.640 231.930 29.870 ;
        RECT 232.545 29.825 232.865 29.885 ;
        RECT 233.480 29.825 233.770 29.870 ;
        RECT 232.545 29.685 233.770 29.825 ;
        RECT 210.940 29.345 213.545 29.485 ;
        RECT 210.940 29.300 211.230 29.345 ;
        RECT 193.920 29.145 194.210 29.190 ;
        RECT 190.315 29.005 194.210 29.145 ;
        RECT 190.315 28.185 190.455 29.005 ;
        RECT 193.920 28.960 194.210 29.005 ;
        RECT 198.980 28.960 199.270 29.190 ;
        RECT 199.445 29.145 199.735 29.190 ;
        RECT 201.280 29.145 201.570 29.190 ;
        RECT 204.860 29.145 205.150 29.190 ;
        RECT 199.445 29.005 205.150 29.145 ;
        RECT 199.445 28.960 199.735 29.005 ;
        RECT 201.280 28.960 201.570 29.005 ;
        RECT 204.860 28.960 205.150 29.005 ;
        RECT 205.405 29.145 205.725 29.205 ;
        RECT 205.940 29.145 206.230 29.300 ;
        RECT 213.225 29.285 213.545 29.345 ;
        RECT 215.540 29.300 215.830 29.530 ;
        RECT 217.820 29.485 218.470 29.530 ;
        RECT 221.420 29.485 221.710 29.530 ;
        RECT 217.820 29.345 221.710 29.485 ;
        RECT 217.820 29.300 218.470 29.345 ;
        RECT 221.120 29.300 221.710 29.345 ;
        RECT 205.405 29.005 206.230 29.145 ;
        RECT 205.405 28.945 205.725 29.005 ;
        RECT 205.940 28.985 206.230 29.005 ;
        RECT 214.145 28.945 214.465 29.205 ;
        RECT 214.625 29.145 214.915 29.190 ;
        RECT 216.460 29.145 216.750 29.190 ;
        RECT 220.040 29.145 220.330 29.190 ;
        RECT 214.625 29.005 220.330 29.145 ;
        RECT 214.625 28.960 214.915 29.005 ;
        RECT 216.460 28.960 216.750 29.005 ;
        RECT 220.040 28.960 220.330 29.005 ;
        RECT 220.585 29.145 220.905 29.205 ;
        RECT 221.120 29.145 221.410 29.300 ;
        RECT 229.800 29.145 230.090 29.190 ;
        RECT 231.715 29.145 231.855 29.640 ;
        RECT 232.545 29.625 232.865 29.685 ;
        RECT 233.480 29.640 233.770 29.685 ;
        RECT 233.925 29.625 234.245 29.885 ;
        RECT 277.165 29.625 277.485 29.885 ;
        RECT 277.625 29.825 277.945 29.885 ;
        RECT 277.625 29.685 280.615 29.825 ;
        RECT 277.625 29.625 277.945 29.685 ;
        RECT 267.505 29.485 267.825 29.545 ;
        RECT 272.105 29.530 272.425 29.545 ;
        RECT 269.360 29.485 269.650 29.530 ;
        RECT 267.505 29.345 269.650 29.485 ;
        RECT 267.505 29.285 267.825 29.345 ;
        RECT 269.360 29.300 269.650 29.345 ;
        RECT 271.640 29.485 272.425 29.530 ;
        RECT 275.240 29.485 275.530 29.530 ;
        RECT 271.640 29.345 275.530 29.485 ;
        RECT 271.640 29.300 272.425 29.345 ;
        RECT 272.105 29.285 272.425 29.300 ;
        RECT 274.940 29.300 275.530 29.345 ;
        RECT 220.585 29.005 222.195 29.145 ;
        RECT 220.585 28.945 220.905 29.005 ;
        RECT 221.120 28.985 221.410 29.005 ;
        RECT 193.000 28.805 193.290 28.850 ;
        RECT 195.285 28.805 195.605 28.865 ;
        RECT 203.105 28.805 203.425 28.865 ;
        RECT 210.020 28.805 210.310 28.850 ;
        RECT 193.000 28.665 210.695 28.805 ;
        RECT 193.000 28.620 193.290 28.665 ;
        RECT 195.285 28.605 195.605 28.665 ;
        RECT 203.105 28.605 203.425 28.665 ;
        RECT 210.020 28.620 210.310 28.665 ;
        RECT 199.850 28.465 200.140 28.510 ;
        RECT 201.740 28.465 202.030 28.510 ;
        RECT 204.860 28.465 205.150 28.510 ;
        RECT 199.850 28.325 205.150 28.465 ;
        RECT 199.850 28.280 200.140 28.325 ;
        RECT 201.740 28.280 202.030 28.325 ;
        RECT 204.860 28.280 205.150 28.325 ;
        RECT 164.005 27.925 164.325 28.185 ;
        RECT 190.225 28.125 190.545 28.185 ;
        RECT 206.325 28.125 206.645 28.185 ;
        RECT 207.720 28.125 208.010 28.170 ;
        RECT 190.225 27.985 208.010 28.125 ;
        RECT 210.555 28.125 210.695 28.665 ;
        RECT 215.030 28.465 215.320 28.510 ;
        RECT 216.920 28.465 217.210 28.510 ;
        RECT 220.040 28.465 220.330 28.510 ;
        RECT 215.030 28.325 220.330 28.465 ;
        RECT 215.030 28.280 215.320 28.325 ;
        RECT 216.920 28.280 217.210 28.325 ;
        RECT 220.040 28.280 220.330 28.325 ;
        RECT 221.045 28.265 221.365 28.525 ;
        RECT 222.055 28.465 222.195 29.005 ;
        RECT 229.800 29.005 231.855 29.145 ;
        RECT 264.745 29.145 265.065 29.205 ;
        RECT 267.980 29.145 268.270 29.190 ;
        RECT 264.745 29.005 268.270 29.145 ;
        RECT 229.800 28.960 230.090 29.005 ;
        RECT 264.745 28.945 265.065 29.005 ;
        RECT 267.980 28.960 268.270 29.005 ;
        RECT 268.445 29.145 268.735 29.190 ;
        RECT 270.280 29.145 270.570 29.190 ;
        RECT 273.860 29.145 274.150 29.190 ;
        RECT 268.445 29.005 274.150 29.145 ;
        RECT 268.445 28.960 268.735 29.005 ;
        RECT 270.280 28.960 270.570 29.005 ;
        RECT 273.860 28.960 274.150 29.005 ;
        RECT 274.940 28.985 275.230 29.300 ;
        RECT 277.255 29.145 277.395 29.625 ;
        RECT 279.610 29.485 279.900 29.530 ;
        RECT 279.555 29.300 279.900 29.485 ;
        RECT 278.100 29.145 278.390 29.190 ;
        RECT 277.255 29.005 278.390 29.145 ;
        RECT 278.100 28.960 278.390 29.005 ;
        RECT 278.545 28.945 278.865 29.205 ;
        RECT 279.020 28.960 279.310 29.190 ;
        RECT 228.865 28.805 229.185 28.865 ;
        RECT 234.400 28.805 234.690 28.850 ;
        RECT 228.865 28.665 234.690 28.805 ;
        RECT 228.865 28.605 229.185 28.665 ;
        RECT 234.400 28.620 234.690 28.665 ;
        RECT 269.345 28.805 269.665 28.865 ;
        RECT 276.705 28.805 277.025 28.865 ;
        RECT 277.180 28.805 277.470 28.850 ;
        RECT 269.345 28.665 274.635 28.805 ;
        RECT 269.345 28.605 269.665 28.665 ;
        RECT 233.465 28.465 233.785 28.525 ;
        RECT 222.055 28.325 233.785 28.465 ;
        RECT 233.465 28.265 233.785 28.325 ;
        RECT 268.850 28.465 269.140 28.510 ;
        RECT 270.740 28.465 271.030 28.510 ;
        RECT 273.860 28.465 274.150 28.510 ;
        RECT 268.850 28.325 274.150 28.465 ;
        RECT 274.495 28.465 274.635 28.665 ;
        RECT 276.705 28.665 277.470 28.805 ;
        RECT 276.705 28.605 277.025 28.665 ;
        RECT 277.180 28.620 277.470 28.665 ;
        RECT 279.095 28.465 279.235 28.960 ;
        RECT 279.555 28.805 279.695 29.300 ;
        RECT 280.475 29.190 280.615 29.685 ;
        RECT 280.845 29.625 281.165 29.885 ;
        RECT 281.305 29.625 281.625 29.885 ;
        RECT 282.225 29.625 282.545 29.885 ;
        RECT 282.685 29.625 283.005 29.885 ;
        RECT 295.105 29.625 295.425 29.885 ;
        RECT 299.720 29.825 300.010 29.870 ;
        RECT 303.845 29.825 304.165 29.885 ;
        RECT 299.720 29.685 304.165 29.825 ;
        RECT 299.720 29.640 300.010 29.685 ;
        RECT 303.845 29.625 304.165 29.685 ;
        RECT 305.225 29.625 305.545 29.885 ;
        RECT 280.400 28.960 280.690 29.190 ;
        RECT 281.395 29.145 281.535 29.625 ;
        RECT 282.315 29.190 282.455 29.625 ;
        RECT 282.775 29.190 282.915 29.625 ;
        RECT 283.145 29.530 283.465 29.545 ;
        RECT 283.145 29.300 283.580 29.530 ;
        RECT 301.200 29.485 301.490 29.530 ;
        RECT 304.440 29.485 305.090 29.530 ;
        RECT 305.315 29.485 305.455 29.625 ;
        RECT 301.200 29.345 305.455 29.485 ;
        RECT 305.685 29.485 306.005 29.545 ;
        RECT 307.080 29.485 307.370 29.530 ;
        RECT 305.685 29.345 307.370 29.485 ;
        RECT 301.200 29.300 301.790 29.345 ;
        RECT 304.440 29.300 305.090 29.345 ;
        RECT 283.145 29.285 283.465 29.300 ;
        RECT 281.780 29.145 282.070 29.190 ;
        RECT 281.395 29.005 282.070 29.145 ;
        RECT 281.780 28.960 282.070 29.005 ;
        RECT 282.240 28.960 282.530 29.190 ;
        RECT 282.700 28.960 282.990 29.190 ;
        RECT 283.235 28.805 283.375 29.285 ;
        RECT 284.065 28.945 284.385 29.205 ;
        RECT 295.580 29.145 295.870 29.190 ;
        RECT 297.865 29.145 298.185 29.205 ;
        RECT 295.580 29.005 298.185 29.145 ;
        RECT 295.580 28.960 295.870 29.005 ;
        RECT 297.865 28.945 298.185 29.005 ;
        RECT 301.500 28.985 301.790 29.300 ;
        RECT 305.685 29.285 306.005 29.345 ;
        RECT 307.080 29.300 307.370 29.345 ;
        RECT 302.580 29.145 302.870 29.190 ;
        RECT 306.160 29.145 306.450 29.190 ;
        RECT 307.995 29.145 308.285 29.190 ;
        RECT 302.580 29.005 308.285 29.145 ;
        RECT 302.580 28.960 302.870 29.005 ;
        RECT 306.160 28.960 306.450 29.005 ;
        RECT 307.995 28.960 308.285 29.005 ;
        RECT 308.445 28.945 308.765 29.205 ;
        RECT 279.555 28.665 283.375 28.805 ;
        RECT 274.495 28.325 279.235 28.465 ;
        RECT 268.850 28.280 269.140 28.325 ;
        RECT 270.740 28.280 271.030 28.325 ;
        RECT 273.860 28.280 274.150 28.325 ;
        RECT 279.465 28.265 279.785 28.525 ;
        RECT 302.580 28.465 302.870 28.510 ;
        RECT 305.700 28.465 305.990 28.510 ;
        RECT 307.590 28.465 307.880 28.510 ;
        RECT 302.580 28.325 307.880 28.465 ;
        RECT 302.580 28.280 302.870 28.325 ;
        RECT 305.700 28.280 305.990 28.325 ;
        RECT 307.590 28.280 307.880 28.325 ;
        RECT 221.135 28.125 221.275 28.265 ;
        RECT 210.555 27.985 221.275 28.125 ;
        RECT 230.720 28.125 231.010 28.170 ;
        RECT 234.385 28.125 234.705 28.185 ;
        RECT 230.720 27.985 234.705 28.125 ;
        RECT 190.225 27.925 190.545 27.985 ;
        RECT 206.325 27.925 206.645 27.985 ;
        RECT 207.720 27.940 208.010 27.985 ;
        RECT 230.720 27.940 231.010 27.985 ;
        RECT 234.385 27.925 234.705 27.985 ;
        RECT 276.720 28.125 277.010 28.170 ;
        RECT 279.555 28.125 279.695 28.265 ;
        RECT 276.720 27.985 279.695 28.125 ;
        RECT 276.720 27.940 277.010 27.985 ;
        RECT 162.095 27.305 311.135 27.785 ;
        RECT 186.085 27.105 186.405 27.165 ;
        RECT 188.400 27.105 188.690 27.150 ;
        RECT 186.085 26.965 188.690 27.105 ;
        RECT 186.085 26.905 186.405 26.965 ;
        RECT 188.400 26.920 188.690 26.965 ;
        RECT 201.725 26.905 202.045 27.165 ;
        RECT 205.405 26.905 205.725 27.165 ;
        RECT 265.665 27.105 265.985 27.165 ;
        RECT 271.660 27.105 271.950 27.150 ;
        RECT 265.665 26.965 271.950 27.105 ;
        RECT 265.665 26.905 265.985 26.965 ;
        RECT 271.660 26.920 271.950 26.965 ;
        RECT 190.685 26.225 191.005 26.485 ;
        RECT 191.605 26.225 191.925 26.485 ;
        RECT 190.225 25.885 190.545 26.145 ;
        RECT 202.660 26.085 202.950 26.130 ;
        RECT 204.025 26.085 204.345 26.145 ;
        RECT 202.660 25.945 204.345 26.085 ;
        RECT 202.660 25.900 202.950 25.945 ;
        RECT 204.025 25.885 204.345 25.945 ;
        RECT 266.585 26.085 266.905 26.145 ;
        RECT 273.040 26.085 273.330 26.130 ;
        RECT 266.585 25.945 273.330 26.085 ;
        RECT 266.585 25.885 266.905 25.945 ;
        RECT 273.040 25.900 273.330 25.945 ;
        RECT 199.885 25.745 200.205 25.805 ;
        RECT 204.960 25.745 205.250 25.790 ;
        RECT 199.885 25.605 205.250 25.745 ;
        RECT 199.885 25.545 200.205 25.605 ;
        RECT 204.960 25.560 205.250 25.605 ;
        RECT 162.095 24.585 311.935 25.065 ;
        RECT 162.095 21.865 311.135 22.345 ;
        RECT 162.095 19.145 311.935 19.625 ;
        RECT 135.120 14.050 138.400 18.845 ;
        RECT 146.290 14.050 155.900 18.845 ;
        RECT 162.095 16.425 311.135 16.905 ;
        RECT 135.120 4.900 155.900 14.050 ;
        RECT 162.095 13.705 311.935 14.185 ;
        RECT 4.100 4.100 155.900 4.900 ;
      LAYER met2 ;
        RECT 45.340 224.760 45.740 225.560 ;
        RECT 64.710 225.410 217.040 225.710 ;
        RECT 64.710 225.310 65.510 225.410 ;
        RECT 59.190 224.760 59.990 225.160 ;
        RECT 67.470 224.810 207.380 225.110 ;
        RECT 67.470 224.710 68.270 224.810 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.210 197.720 224.510 ;
        RECT 70.230 224.110 71.030 224.210 ;
        RECT 72.990 223.610 188.060 223.910 ;
        RECT 72.990 223.510 73.790 223.610 ;
        RECT 75.700 223.010 178.400 223.310 ;
        RECT 75.700 222.910 76.500 223.010 ;
        RECT 78.545 222.410 168.740 222.710 ;
        RECT 78.545 222.310 79.345 222.410 ;
        RECT 83.980 221.810 164.500 222.110 ;
        RECT 83.980 221.710 84.780 221.810 ;
        RECT 86.740 221.210 163.500 221.510 ;
        RECT 164.100 221.310 164.500 221.810 ;
        RECT 86.740 221.110 87.540 221.210 ;
        RECT 92.260 220.610 162.500 220.910 ;
        RECT 163.100 220.710 163.500 221.210 ;
        RECT 92.260 220.510 93.060 220.610 ;
        RECT 162.100 220.110 162.500 220.610 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.495 208.765 51.905 210.765 ;
        RECT 9.495 205.765 45.165 207.765 ;
        RECT 51.315 207.460 51.905 208.765 ;
        RECT 9.495 202.765 48.270 204.765 ;
        RECT 9.495 198.745 48.270 200.745 ;
        RECT 9.495 195.745 45.165 197.745 ;
        RECT 9.495 192.745 46.670 194.745 ;
        RECT 9.495 187.420 15.245 188.980 ;
        RECT 16.515 188.295 45.165 190.295 ;
        RECT 52.860 188.465 54.245 190.570 ;
        RECT 16.515 184.775 56.920 186.775 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.495 182.570 15.245 184.130 ;
        RECT 16.515 181.255 46.670 183.255 ;
        RECT 5.910 176.050 7.510 179.250 ;
        RECT 57.020 178.865 57.820 178.990 ;
        RECT 9.500 177.365 58.420 178.865 ;
        RECT 53.870 176.720 54.670 176.890 ;
        RECT 9.500 175.220 54.670 176.720 ;
        RECT 9.500 172.820 54.670 174.320 ;
        RECT 53.870 172.640 54.670 172.820 ;
        RECT 52.220 171.920 53.020 172.040 ;
        RECT 9.500 170.420 53.020 171.920 ;
        RECT 63.470 170.855 65.220 217.105 ;
        RECT 66.220 170.855 67.970 217.105 ;
        RECT 68.970 170.855 70.720 217.105 ;
        RECT 71.720 170.855 73.470 217.105 ;
        RECT 74.470 170.855 76.220 217.105 ;
        RECT 77.220 170.855 78.970 217.105 ;
        RECT 79.970 170.115 81.970 217.845 ;
        RECT 106.340 217.515 107.940 219.915 ;
        RECT 109.240 219.705 111.675 220.105 ;
        RECT 113.270 219.705 115.705 220.105 ;
        RECT 117.300 219.705 119.735 220.105 ;
        RECT 121.330 219.705 123.765 220.105 ;
        RECT 125.360 219.705 127.795 220.105 ;
        RECT 129.390 219.705 131.825 220.105 ;
        RECT 133.420 219.705 135.855 220.105 ;
        RECT 137.450 219.705 139.885 220.105 ;
        RECT 141.480 219.705 143.915 220.105 ;
        RECT 145.510 219.705 147.945 220.105 ;
        RECT 149.540 219.705 151.975 220.105 ;
        RECT 109.240 217.705 109.640 219.705 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 111.820 217.295 112.220 219.305 ;
        RECT 113.270 217.705 113.670 219.705 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 115.850 217.295 116.250 219.305 ;
        RECT 117.300 217.705 117.700 219.705 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 119.880 217.295 120.280 219.305 ;
        RECT 121.330 217.705 121.730 219.705 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 123.910 217.295 124.310 219.305 ;
        RECT 125.360 217.705 125.760 219.705 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 127.940 217.295 128.340 219.305 ;
        RECT 129.390 217.705 129.790 219.705 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 131.970 217.295 132.370 219.305 ;
        RECT 133.420 217.705 133.820 219.705 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 136.000 217.295 136.400 219.305 ;
        RECT 137.450 217.705 137.850 219.705 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 140.030 217.295 140.430 219.305 ;
        RECT 141.480 217.705 141.880 219.705 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 144.060 217.295 144.460 219.305 ;
        RECT 145.510 217.705 145.910 219.705 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 148.090 217.295 148.490 219.305 ;
        RECT 149.540 217.705 149.940 219.705 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 152.120 217.295 152.520 219.305 ;
        RECT 82.970 170.855 84.720 217.105 ;
        RECT 85.720 170.855 87.470 217.105 ;
        RECT 88.470 170.855 90.220 217.105 ;
        RECT 91.220 170.855 92.970 217.105 ;
        RECT 93.970 170.855 95.720 217.105 ;
        RECT 96.720 170.855 98.470 217.105 ;
        RECT 109.785 216.895 112.220 217.295 ;
        RECT 113.815 216.895 116.250 217.295 ;
        RECT 117.845 216.895 120.280 217.295 ;
        RECT 121.875 216.895 124.310 217.295 ;
        RECT 125.905 216.895 128.340 217.295 ;
        RECT 129.935 216.895 132.370 217.295 ;
        RECT 133.965 216.895 136.400 217.295 ;
        RECT 137.995 216.895 140.430 217.295 ;
        RECT 142.025 216.895 144.460 217.295 ;
        RECT 146.055 216.895 148.490 217.295 ;
        RECT 150.085 216.895 152.520 217.295 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 111.820 205.955 112.220 206.755 ;
        RECT 115.850 205.955 116.250 206.755 ;
        RECT 119.880 205.955 120.280 206.755 ;
        RECT 123.910 205.955 124.310 206.755 ;
        RECT 127.940 205.955 128.340 206.755 ;
        RECT 131.970 205.955 132.370 206.755 ;
        RECT 136.000 205.955 136.400 206.755 ;
        RECT 140.030 205.955 140.430 206.755 ;
        RECT 144.060 205.955 144.460 206.755 ;
        RECT 148.090 205.955 148.490 206.755 ;
        RECT 152.120 205.955 152.520 206.755 ;
        RECT 109.240 204.745 111.675 205.545 ;
        RECT 113.270 204.745 115.705 205.545 ;
        RECT 117.300 204.745 119.735 205.545 ;
        RECT 121.330 204.745 123.765 205.545 ;
        RECT 125.360 204.745 127.795 205.545 ;
        RECT 129.390 204.745 131.825 205.545 ;
        RECT 133.420 204.745 135.855 205.545 ;
        RECT 137.450 204.745 139.885 205.545 ;
        RECT 141.480 204.745 143.915 205.545 ;
        RECT 145.510 204.745 147.945 205.545 ;
        RECT 149.540 204.745 151.975 205.545 ;
        RECT 108.540 202.425 108.940 202.625 ;
        RECT 109.785 202.425 110.385 204.345 ;
        RECT 108.540 202.025 110.385 202.425 ;
        RECT 108.540 201.825 108.940 202.025 ;
        RECT 109.785 199.970 110.385 202.025 ;
        RECT 111.075 199.970 111.675 204.745 ;
        RECT 112.570 202.425 112.970 202.625 ;
        RECT 113.815 202.425 114.415 204.345 ;
        RECT 112.570 202.025 114.415 202.425 ;
        RECT 112.570 201.825 112.970 202.025 ;
        RECT 113.815 199.970 114.415 202.025 ;
        RECT 115.105 199.970 115.705 204.745 ;
        RECT 116.600 202.425 117.000 202.625 ;
        RECT 117.845 202.425 118.445 204.345 ;
        RECT 116.600 202.025 118.445 202.425 ;
        RECT 116.600 201.825 117.000 202.025 ;
        RECT 117.845 199.970 118.445 202.025 ;
        RECT 119.135 199.970 119.735 204.745 ;
        RECT 120.630 202.425 121.030 202.625 ;
        RECT 121.875 202.425 122.475 204.345 ;
        RECT 120.630 202.025 122.475 202.425 ;
        RECT 120.630 201.825 121.030 202.025 ;
        RECT 121.875 199.970 122.475 202.025 ;
        RECT 123.165 199.970 123.765 204.745 ;
        RECT 124.660 202.425 125.060 202.625 ;
        RECT 125.905 202.425 126.505 204.345 ;
        RECT 124.660 202.025 126.505 202.425 ;
        RECT 124.660 201.825 125.060 202.025 ;
        RECT 125.905 199.970 126.505 202.025 ;
        RECT 127.195 199.970 127.795 204.745 ;
        RECT 128.690 202.425 129.090 202.625 ;
        RECT 129.935 202.425 130.535 204.345 ;
        RECT 128.690 202.025 130.535 202.425 ;
        RECT 128.690 201.825 129.090 202.025 ;
        RECT 129.935 199.970 130.535 202.025 ;
        RECT 131.225 199.970 131.825 204.745 ;
        RECT 132.720 202.425 133.120 202.625 ;
        RECT 133.965 202.425 134.565 204.345 ;
        RECT 132.720 202.025 134.565 202.425 ;
        RECT 132.720 201.825 133.120 202.025 ;
        RECT 133.965 199.970 134.565 202.025 ;
        RECT 135.255 199.970 135.855 204.745 ;
        RECT 136.750 202.425 137.150 202.625 ;
        RECT 137.995 202.425 138.595 204.345 ;
        RECT 136.750 202.025 138.595 202.425 ;
        RECT 136.750 201.825 137.150 202.025 ;
        RECT 137.995 199.970 138.595 202.025 ;
        RECT 139.285 199.970 139.885 204.745 ;
        RECT 140.780 202.425 141.180 202.625 ;
        RECT 142.025 202.425 142.625 204.345 ;
        RECT 140.780 202.025 142.625 202.425 ;
        RECT 140.780 201.825 141.180 202.025 ;
        RECT 142.025 199.970 142.625 202.025 ;
        RECT 143.315 199.970 143.915 204.745 ;
        RECT 144.810 202.425 145.210 202.625 ;
        RECT 146.055 202.425 146.655 204.345 ;
        RECT 144.810 202.025 146.655 202.425 ;
        RECT 144.810 201.825 145.210 202.025 ;
        RECT 146.055 199.970 146.655 202.025 ;
        RECT 147.345 199.970 147.945 204.745 ;
        RECT 148.840 202.425 149.240 202.625 ;
        RECT 150.085 202.425 150.685 204.345 ;
        RECT 148.840 202.025 150.685 202.425 ;
        RECT 148.840 201.825 149.240 202.025 ;
        RECT 150.085 199.970 150.685 202.025 ;
        RECT 151.375 199.970 151.975 204.745 ;
        RECT 168.460 202.290 168.740 222.410 ;
        RECT 178.120 202.290 178.400 223.010 ;
        RECT 187.780 202.290 188.060 223.610 ;
        RECT 197.440 202.290 197.720 224.210 ;
        RECT 207.100 202.290 207.380 224.810 ;
        RECT 216.760 202.290 217.040 225.410 ;
        RECT 246.615 225.060 247.015 225.660 ;
        RECT 226.420 224.460 226.700 224.510 ;
        RECT 236.020 224.460 236.420 225.060 ;
        RECT 226.360 223.860 226.760 224.460 ;
        RECT 226.420 202.290 226.700 223.860 ;
        RECT 236.080 202.290 236.360 224.460 ;
        RECT 246.665 218.450 246.965 225.060 ;
        RECT 246.615 217.650 247.015 218.450 ;
        RECT 168.530 201.140 168.670 202.290 ;
        RECT 173.635 201.305 175.175 201.675 ;
        RECT 178.190 201.140 178.330 202.290 ;
        RECT 187.850 201.140 187.990 202.290 ;
        RECT 192.145 201.305 193.685 201.675 ;
        RECT 197.510 201.140 197.650 202.290 ;
        RECT 207.170 201.140 207.310 202.290 ;
        RECT 210.655 201.305 212.195 201.675 ;
        RECT 216.830 201.140 216.970 202.290 ;
        RECT 226.490 201.140 226.630 202.290 ;
        RECT 229.165 201.305 230.705 201.675 ;
        RECT 236.150 201.140 236.290 202.290 ;
        RECT 168.470 200.820 168.730 201.140 ;
        RECT 178.130 200.820 178.390 201.140 ;
        RECT 187.790 200.820 188.050 201.140 ;
        RECT 197.450 200.820 197.710 201.140 ;
        RECT 207.110 200.820 207.370 201.140 ;
        RECT 216.770 200.820 217.030 201.140 ;
        RECT 226.430 200.820 226.690 201.140 ;
        RECT 236.090 200.820 236.350 201.140 ;
        RECT 166.630 199.800 166.890 200.120 ;
        RECT 178.590 199.800 178.850 200.120 ;
        RECT 189.630 199.800 189.890 200.120 ;
        RECT 199.290 199.800 199.550 200.120 ;
        RECT 208.950 199.800 209.210 200.120 ;
        RECT 226.890 199.800 227.150 200.120 ;
        RECT 236.090 199.800 236.350 200.120 ;
        RECT 109.240 194.440 109.640 199.685 ;
        RECT 109.240 194.040 110.255 194.440 ;
        RECT 109.240 191.285 109.640 192.885 ;
        RECT 110.530 187.540 110.930 198.905 ;
        RECT 111.820 194.440 112.220 199.685 ;
        RECT 111.205 194.040 112.220 194.440 ;
        RECT 113.270 194.440 113.670 199.685 ;
        RECT 113.270 194.040 114.285 194.440 ;
        RECT 111.820 191.285 112.220 192.885 ;
        RECT 113.270 191.285 113.670 192.885 ;
        RECT 114.560 187.540 114.960 198.905 ;
        RECT 115.850 194.440 116.250 199.685 ;
        RECT 115.235 194.040 116.250 194.440 ;
        RECT 117.300 194.440 117.700 199.685 ;
        RECT 117.300 194.040 118.315 194.440 ;
        RECT 115.850 191.285 116.250 192.885 ;
        RECT 117.300 191.285 117.700 192.885 ;
        RECT 118.590 187.540 118.990 198.905 ;
        RECT 119.880 194.440 120.280 199.685 ;
        RECT 119.265 194.040 120.280 194.440 ;
        RECT 121.330 194.440 121.730 199.685 ;
        RECT 121.330 194.040 122.345 194.440 ;
        RECT 119.880 191.285 120.280 192.885 ;
        RECT 121.330 191.285 121.730 192.885 ;
        RECT 122.620 187.540 123.020 198.905 ;
        RECT 123.910 194.440 124.310 199.685 ;
        RECT 123.295 194.040 124.310 194.440 ;
        RECT 125.360 194.440 125.760 199.685 ;
        RECT 125.360 194.040 126.375 194.440 ;
        RECT 123.910 191.285 124.310 192.885 ;
        RECT 125.360 191.285 125.760 192.885 ;
        RECT 126.650 187.540 127.050 198.905 ;
        RECT 127.940 194.440 128.340 199.685 ;
        RECT 127.325 194.040 128.340 194.440 ;
        RECT 129.390 194.440 129.790 199.685 ;
        RECT 129.390 194.040 130.405 194.440 ;
        RECT 127.940 191.285 128.340 192.885 ;
        RECT 129.390 191.285 129.790 192.885 ;
        RECT 130.680 187.540 131.080 198.905 ;
        RECT 131.970 194.440 132.370 199.685 ;
        RECT 131.355 194.040 132.370 194.440 ;
        RECT 133.420 194.440 133.820 199.685 ;
        RECT 133.420 194.040 134.435 194.440 ;
        RECT 131.970 191.285 132.370 192.885 ;
        RECT 133.420 191.285 133.820 192.885 ;
        RECT 134.710 187.540 135.110 198.905 ;
        RECT 136.000 194.440 136.400 199.685 ;
        RECT 135.385 194.040 136.400 194.440 ;
        RECT 137.450 194.440 137.850 199.685 ;
        RECT 137.450 194.040 138.465 194.440 ;
        RECT 136.000 191.285 136.400 192.885 ;
        RECT 137.450 191.285 137.850 192.885 ;
        RECT 138.740 187.540 139.140 198.905 ;
        RECT 140.030 194.440 140.430 199.685 ;
        RECT 139.415 194.040 140.430 194.440 ;
        RECT 141.480 194.440 141.880 199.685 ;
        RECT 141.480 194.040 142.495 194.440 ;
        RECT 140.030 191.285 140.430 192.885 ;
        RECT 141.480 191.285 141.880 192.885 ;
        RECT 142.770 187.540 143.170 198.905 ;
        RECT 144.060 194.440 144.460 199.685 ;
        RECT 143.445 194.040 144.460 194.440 ;
        RECT 145.510 194.440 145.910 199.685 ;
        RECT 145.510 194.040 146.525 194.440 ;
        RECT 144.060 191.285 144.460 192.885 ;
        RECT 145.510 191.285 145.910 192.885 ;
        RECT 146.800 187.540 147.200 198.905 ;
        RECT 148.090 194.440 148.490 199.685 ;
        RECT 147.475 194.040 148.490 194.440 ;
        RECT 149.540 194.440 149.940 199.685 ;
        RECT 149.540 194.040 150.555 194.440 ;
        RECT 148.090 191.285 148.490 192.885 ;
        RECT 149.540 191.285 149.940 192.885 ;
        RECT 150.830 187.540 151.230 198.905 ;
        RECT 152.120 194.440 152.520 199.685 ;
        RECT 166.690 197.935 166.830 199.800 ;
        RECT 169.850 199.460 170.110 199.780 ;
        RECT 166.620 197.565 166.900 197.935 ;
        RECT 151.505 194.040 152.520 194.440 ;
        RECT 152.120 191.285 152.520 192.885 ;
        RECT 168.930 191.300 169.190 191.620 ;
        RECT 166.630 188.920 166.890 189.240 ;
        RECT 161.590 188.380 162.390 188.430 ;
        RECT 166.690 188.415 166.830 188.920 ;
        RECT 158.335 188.080 162.390 188.380 ;
        RECT 109.240 184.370 109.640 184.770 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 158.335 187.580 158.735 188.080 ;
        RECT 161.590 188.030 162.390 188.080 ;
        RECT 166.620 188.045 166.900 188.415 ;
        RECT 167.550 185.860 167.810 186.180 ;
        RECT 167.610 184.820 167.750 185.860 ;
        RECT 167.550 184.500 167.810 184.820 ;
        RECT 109.240 183.970 154.345 184.370 ;
        RECT 153.945 183.570 154.345 183.970 ;
        RECT 166.630 183.480 166.890 183.800 ;
        RECT 168.010 183.480 168.270 183.800 ;
        RECT 161.590 178.860 162.390 178.910 ;
        RECT 157.560 178.560 162.390 178.860 ;
        RECT 115.265 175.815 117.965 176.215 ;
        RECT 119.885 175.815 122.585 176.215 ;
        RECT 124.505 175.815 127.205 176.215 ;
        RECT 129.125 175.815 131.825 176.215 ;
        RECT 133.745 175.815 136.445 176.215 ;
        RECT 138.365 175.815 141.065 176.215 ;
        RECT 142.985 175.815 145.685 176.215 ;
        RECT 147.605 175.815 150.305 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 157.560 178.060 157.960 178.560 ;
        RECT 161.590 178.510 162.390 178.560 ;
        RECT 166.690 176.320 166.830 183.480 ;
        RECT 167.090 181.100 167.350 181.420 ;
        RECT 167.150 178.895 167.290 181.100 ;
        RECT 167.080 178.525 167.360 178.895 ;
        RECT 167.550 178.040 167.810 178.360 ;
        RECT 166.630 176.000 166.890 176.320 ;
        RECT 167.610 175.640 167.750 178.040 ;
        RECT 168.070 176.660 168.210 183.480 ;
        RECT 168.460 183.285 168.740 183.655 ;
        RECT 168.530 179.380 168.670 183.285 ;
        RECT 168.990 182.100 169.130 191.300 ;
        RECT 169.910 190.260 170.050 199.460 ;
        RECT 172.150 199.120 172.410 199.440 ;
        RECT 171.230 191.640 171.490 191.960 ;
        RECT 169.850 189.940 170.110 190.260 ;
        RECT 170.760 188.725 171.040 189.095 ;
        RECT 169.840 188.045 170.120 188.415 ;
        RECT 170.310 188.240 170.570 188.560 ;
        RECT 169.910 186.860 170.050 188.045 ;
        RECT 170.370 186.860 170.510 188.240 ;
        RECT 170.830 187.540 170.970 188.725 ;
        RECT 171.290 188.470 171.430 191.640 ;
        RECT 171.690 188.470 171.950 188.560 ;
        RECT 171.290 188.330 171.950 188.470 ;
        RECT 171.690 188.240 171.950 188.330 ;
        RECT 170.770 187.220 171.030 187.540 ;
        RECT 171.750 186.860 171.890 188.240 ;
        RECT 169.850 186.540 170.110 186.860 ;
        RECT 170.310 186.540 170.570 186.860 ;
        RECT 171.690 186.540 171.950 186.860 ;
        RECT 169.850 185.520 170.110 185.840 ;
        RECT 168.930 181.780 169.190 182.100 ;
        RECT 169.390 181.100 169.650 181.420 ;
        RECT 168.930 180.080 169.190 180.400 ;
        RECT 168.470 179.060 168.730 179.380 ;
        RECT 168.990 178.360 169.130 180.080 ;
        RECT 169.450 179.040 169.590 181.100 ;
        RECT 169.390 178.720 169.650 179.040 ;
        RECT 169.910 178.360 170.050 185.520 ;
        RECT 170.370 184.820 170.510 186.540 ;
        RECT 170.770 186.260 171.030 186.520 ;
        RECT 170.770 186.200 171.430 186.260 ;
        RECT 170.830 186.120 171.430 186.200 ;
        RECT 170.770 185.520 171.030 185.840 ;
        RECT 170.310 184.500 170.570 184.820 ;
        RECT 170.830 183.800 170.970 185.520 ;
        RECT 170.770 183.480 171.030 183.800 ;
        RECT 170.310 182.800 170.570 183.120 ;
        RECT 170.370 181.420 170.510 182.800 ;
        RECT 170.310 181.100 170.570 181.420 ;
        RECT 170.770 181.100 171.030 181.420 ;
        RECT 170.830 179.380 170.970 181.100 ;
        RECT 170.770 179.060 171.030 179.380 ;
        RECT 168.930 178.040 169.190 178.360 ;
        RECT 169.850 178.040 170.110 178.360 ;
        RECT 168.010 176.340 168.270 176.660 ;
        RECT 171.290 176.060 171.430 186.120 ;
        RECT 171.750 181.420 171.890 186.540 ;
        RECT 172.210 184.820 172.350 199.120 ;
        RECT 173.635 195.865 175.175 196.235 ;
        RECT 176.750 193.680 177.010 194.000 ;
        RECT 175.370 191.980 175.630 192.300 ;
        RECT 175.830 191.980 176.090 192.300 ;
        RECT 173.070 190.960 173.330 191.280 ;
        RECT 172.610 188.920 172.870 189.240 ;
        RECT 172.150 184.500 172.410 184.820 ;
        RECT 172.670 184.050 172.810 188.920 ;
        RECT 173.130 184.390 173.270 190.960 ;
        RECT 173.635 190.425 175.175 190.795 ;
        RECT 175.430 189.775 175.570 191.980 ;
        RECT 175.360 189.405 175.640 189.775 ;
        RECT 174.910 188.920 175.170 189.240 ;
        RECT 173.530 188.240 173.790 188.560 ;
        RECT 173.590 187.620 173.730 188.240 ;
        RECT 173.590 187.480 174.190 187.620 ;
        RECT 174.050 186.860 174.190 187.480 ;
        RECT 174.970 187.200 175.110 188.920 ;
        RECT 174.910 186.880 175.170 187.200 ;
        RECT 173.990 186.540 174.250 186.860 ;
        RECT 175.360 186.685 175.640 187.055 ;
        RECT 175.370 186.540 175.630 186.685 ;
        RECT 173.635 184.985 175.175 185.355 ;
        RECT 173.130 184.250 173.730 184.390 ;
        RECT 173.990 184.335 174.250 184.480 ;
        RECT 172.670 183.910 173.270 184.050 ;
        RECT 172.610 183.140 172.870 183.460 ;
        RECT 172.670 182.975 172.810 183.140 ;
        RECT 172.600 182.605 172.880 182.975 ;
        RECT 171.690 181.100 171.950 181.420 ;
        RECT 172.610 180.420 172.870 180.740 ;
        RECT 172.670 178.700 172.810 180.420 ;
        RECT 173.130 179.290 173.270 183.910 ;
        RECT 173.590 181.420 173.730 184.250 ;
        RECT 173.980 183.965 174.260 184.335 ;
        RECT 175.430 184.220 175.570 186.540 ;
        RECT 174.510 184.080 175.570 184.220 ;
        RECT 175.890 184.220 176.030 191.980 ;
        RECT 176.290 190.960 176.550 191.280 ;
        RECT 176.350 190.260 176.490 190.960 ;
        RECT 176.290 189.940 176.550 190.260 ;
        RECT 176.810 188.560 176.950 193.680 ;
        RECT 178.650 192.980 178.790 199.800 ;
        RECT 182.270 199.120 182.530 199.440 ;
        RECT 180.430 194.360 180.690 194.680 ;
        RECT 179.970 194.020 180.230 194.340 ;
        RECT 178.590 192.660 178.850 192.980 ;
        RECT 178.590 191.980 178.850 192.300 ;
        RECT 176.750 188.240 177.010 188.560 ;
        RECT 177.200 188.045 177.480 188.415 ;
        RECT 177.670 188.240 177.930 188.560 ;
        RECT 178.130 188.240 178.390 188.560 ;
        RECT 176.750 186.540 177.010 186.860 ;
        RECT 176.290 186.200 176.550 186.520 ;
        RECT 176.350 184.730 176.490 186.200 ;
        RECT 176.810 185.840 176.950 186.540 ;
        RECT 176.750 185.520 177.010 185.840 ;
        RECT 176.350 184.590 176.950 184.730 ;
        RECT 175.890 184.080 176.490 184.220 ;
        RECT 174.510 183.370 174.650 184.080 ;
        RECT 175.370 183.480 175.630 183.800 ;
        RECT 175.830 183.480 176.090 183.800 ;
        RECT 174.050 183.230 174.650 183.370 ;
        RECT 174.050 181.420 174.190 183.230 ;
        RECT 173.530 181.100 173.790 181.420 ;
        RECT 173.990 181.100 174.250 181.420 ;
        RECT 174.050 180.740 174.190 181.100 ;
        RECT 173.990 180.420 174.250 180.740 ;
        RECT 173.635 179.545 175.175 179.915 ;
        RECT 175.430 179.380 175.570 183.480 ;
        RECT 175.890 179.380 176.030 183.480 ;
        RECT 173.130 179.150 175.110 179.290 ;
        RECT 172.610 178.380 172.870 178.700 ;
        RECT 172.670 176.430 173.270 176.570 ;
        RECT 172.670 176.060 172.810 176.430 ;
        RECT 173.130 176.290 173.270 176.430 ;
        RECT 174.050 176.430 174.650 176.570 ;
        RECT 174.050 176.290 174.190 176.430 ;
        RECT 171.290 175.920 172.810 176.060 ;
        RECT 167.550 175.320 167.810 175.640 ;
        RECT 114.835 172.120 118.395 174.820 ;
        RECT 119.155 172.120 123.015 174.820 ;
        RECT 123.775 172.120 127.635 174.820 ;
        RECT 128.395 172.120 132.255 174.820 ;
        RECT 133.015 172.120 136.875 174.820 ;
        RECT 137.635 172.120 141.495 174.820 ;
        RECT 142.255 172.120 146.115 174.820 ;
        RECT 146.875 172.120 150.735 174.820 ;
        RECT 57.020 169.775 57.820 169.890 ;
        RECT 9.500 168.275 58.420 169.775 ;
        RECT 9.500 165.715 56.920 166.715 ;
        RECT 103.350 164.990 103.750 170.890 ;
        RECT 105.930 168.490 106.330 170.890 ;
        RECT 9.500 163.915 55.070 164.915 ;
        RECT 102.625 164.590 103.750 164.990 ;
        RECT 104.640 164.790 105.040 167.190 ;
        RECT 107.380 164.990 107.780 170.890 ;
        RECT 109.960 168.490 110.360 170.890 ;
        RECT 115.625 169.795 117.605 170.845 ;
        RECT 119.155 169.795 119.755 172.120 ;
        RECT 115.625 169.195 119.755 169.795 ;
        RECT 120.245 169.795 122.225 170.845 ;
        RECT 123.775 169.795 124.375 172.120 ;
        RECT 120.245 169.195 124.375 169.795 ;
        RECT 124.865 169.795 126.845 170.845 ;
        RECT 128.395 169.795 128.995 172.120 ;
        RECT 124.865 169.195 128.995 169.795 ;
        RECT 129.485 169.795 131.465 170.845 ;
        RECT 133.015 169.795 133.615 172.120 ;
        RECT 129.485 169.195 133.615 169.795 ;
        RECT 134.105 169.795 136.085 170.845 ;
        RECT 137.635 169.795 138.235 172.120 ;
        RECT 134.105 169.195 138.235 169.795 ;
        RECT 138.725 169.795 140.705 170.845 ;
        RECT 142.255 169.795 142.855 172.120 ;
        RECT 138.725 169.195 142.855 169.795 ;
        RECT 143.345 169.795 145.325 170.845 ;
        RECT 146.875 169.795 147.475 172.120 ;
        RECT 143.345 169.195 147.475 169.795 ;
        RECT 115.625 168.145 117.605 169.195 ;
        RECT 120.245 168.145 122.225 169.195 ;
        RECT 124.865 168.145 126.845 169.195 ;
        RECT 129.485 168.145 131.465 169.195 ;
        RECT 134.105 168.145 136.085 169.195 ;
        RECT 138.725 168.145 140.705 169.195 ;
        RECT 143.345 168.145 145.325 169.195 ;
        RECT 147.965 168.145 150.345 170.845 ;
        RECT 106.655 164.590 107.780 164.990 ;
        RECT 108.670 164.790 109.070 167.190 ;
        RECT 9.500 162.115 51.610 163.115 ;
        RECT 9.500 159.815 53.170 161.315 ;
        RECT 2.705 157.015 51.610 159.015 ;
        RECT 2.705 1.285 3.505 157.015 ;
        RECT 9.500 154.715 53.170 156.215 ;
        RECT 9.500 152.915 51.610 153.915 ;
        RECT 9.500 151.115 55.070 152.115 ;
        RECT 74.940 151.875 86.100 155.595 ;
        RECT 9.500 149.315 56.520 150.315 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 148.155 78.660 151.875 ;
        RECT 80.100 149.595 80.930 150.425 ;
        RECT 82.380 148.155 86.100 151.875 ;
        RECT 102.625 149.850 103.025 164.590 ;
        RECT 103.350 162.940 104.365 163.340 ;
        RECT 105.315 162.940 106.330 163.340 ;
        RECT 103.350 159.695 103.750 162.940 ;
        RECT 105.930 160.395 106.330 162.940 ;
        RECT 104.190 159.795 106.330 160.395 ;
        RECT 104.190 159.410 104.495 159.795 ;
        RECT 105.930 159.695 106.330 159.795 ;
        RECT 103.895 154.535 104.495 159.410 ;
        RECT 105.185 155.035 105.785 159.410 ;
        RECT 103.895 153.935 106.330 154.535 ;
        RECT 103.350 150.640 103.750 153.565 ;
        RECT 105.930 152.190 106.330 153.935 ;
        RECT 103.895 151.790 106.330 152.190 ;
        RECT 103.895 151.015 104.495 151.790 ;
        RECT 105.185 150.640 105.785 151.415 ;
        RECT 103.350 150.240 105.785 150.640 ;
        RECT 106.655 149.850 107.055 164.590 ;
        RECT 107.380 162.940 108.395 163.340 ;
        RECT 109.345 162.940 110.360 163.340 ;
        RECT 107.380 159.695 107.780 162.940 ;
        RECT 109.960 160.395 110.360 162.940 ;
        RECT 108.220 159.795 110.360 160.395 ;
        RECT 108.220 159.410 108.525 159.795 ;
        RECT 109.960 159.695 110.360 159.795 ;
        RECT 107.925 154.535 108.525 159.410 ;
        RECT 109.215 155.035 109.815 159.410 ;
        RECT 107.925 153.935 110.360 154.535 ;
        RECT 107.380 150.640 107.780 153.565 ;
        RECT 109.960 152.190 110.360 153.935 ;
        RECT 107.925 151.790 110.360 152.190 ;
        RECT 107.925 151.015 108.525 151.790 ;
        RECT 109.215 150.640 109.815 151.415 ;
        RECT 107.380 150.240 109.815 150.640 ;
        RECT 102.625 149.450 103.750 149.850 ;
        RECT 74.940 144.435 86.100 148.155 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 11.195 139.800 23.015 140.200 ;
        RECT 11.195 137.185 11.795 139.800 ;
        RECT 14.860 138.370 21.050 138.770 ;
        RECT 14.860 137.585 15.260 138.370 ;
        RECT 20.650 137.970 21.050 138.370 ;
        RECT 14.130 137.185 16.020 137.585 ;
        RECT 16.805 137.185 18.955 137.585 ;
        RECT 16.805 136.875 17.205 137.185 ;
        RECT 11.940 136.275 15.275 136.875 ;
        RECT 16.165 136.275 17.205 136.875 ;
        RECT 5.910 132.225 7.510 135.425 ;
        RECT 13.485 133.130 14.085 135.875 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 16.805 129.110 17.205 136.275 ;
        RECT 19.100 136.125 20.750 136.725 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 19.100 128.925 19.500 136.125 ;
        RECT 22.615 134.120 23.015 139.800 ;
        RECT 24.255 135.155 25.755 143.745 ;
        RECT 27.765 135.155 29.265 143.745 ;
        RECT 36.055 135.155 37.555 143.745 ;
        RECT 44.345 135.155 45.845 143.745 ;
        RECT 52.635 135.155 54.135 143.745 ;
        RECT 56.145 135.155 57.645 143.745 ;
        RECT 103.350 143.435 103.750 149.450 ;
        RECT 104.640 147.135 105.040 149.535 ;
        RECT 106.655 149.450 107.780 149.850 ;
        RECT 105.930 143.435 106.330 145.835 ;
        RECT 107.380 143.435 107.780 149.450 ;
        RECT 108.670 147.135 109.070 149.535 ;
        RECT 109.960 143.435 110.360 145.835 ;
        RECT 116.310 143.410 116.910 168.145 ;
        RECT 120.930 147.550 121.530 168.145 ;
        RECT 125.550 159.440 126.150 168.145 ;
        RECT 125.550 158.840 128.940 159.440 ;
        RECT 120.930 146.950 126.935 147.550 ;
        RECT 122.645 144.030 124.245 144.830 ;
        RECT 128.340 144.540 128.940 158.840 ;
        RECT 130.170 148.610 130.770 168.145 ;
        RECT 134.795 164.330 135.395 168.145 ;
        RECT 133.685 163.140 134.485 163.740 ;
        RECT 133.785 155.610 134.385 163.140 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 139.410 157.075 140.010 168.145 ;
        RECT 144.035 163.040 144.635 168.145 ;
        RECT 146.855 164.430 147.655 165.030 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 141.615 158.550 142.415 159.150 ;
        RECT 138.070 156.475 140.010 157.075 ;
        RECT 133.285 155.010 134.885 155.610 ;
        RECT 133.275 151.400 134.875 152.200 ;
        RECT 133.275 150.230 134.875 151.030 ;
        RECT 138.070 149.760 138.670 156.475 ;
        RECT 141.715 152.110 142.315 158.550 ;
        RECT 141.215 151.905 142.815 152.110 ;
        RECT 140.950 151.505 143.050 151.905 ;
        RECT 133.285 149.160 138.670 149.760 ;
        RECT 130.170 148.010 134.430 148.610 ;
        RECT 130.615 146.830 132.215 147.630 ;
        RECT 133.285 147.410 134.885 148.010 ;
        RECT 138.525 147.310 140.125 148.110 ;
        RECT 128.340 143.940 134.885 144.540 ;
        RECT 138.525 143.820 140.125 144.620 ;
        RECT 116.310 142.810 132.215 143.410 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 141.990 142.815 142.790 ;
        RECT 146.955 142.730 147.555 164.430 ;
        RECT 148.655 158.450 149.255 168.145 ;
        RECT 146.455 142.640 148.055 142.730 ;
        RECT 146.195 142.240 148.295 142.640 ;
        RECT 146.455 142.130 148.055 142.240 ;
        RECT 104.640 139.365 152.360 140.165 ;
        RECT 97.200 137.420 147.750 138.220 ;
        RECT 107.380 135.525 132.465 136.325 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 56.145 133.555 77.110 135.155 ;
        RECT 80.120 133.320 137.265 134.120 ;
        RECT 137.945 133.410 144.375 133.810 ;
        RECT 21.615 131.745 135.665 132.545 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 142.980 131.990 143.630 132.590 ;
        RECT 27.065 129.995 134.065 130.795 ;
        RECT 19.100 128.125 101.315 128.925 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 142.980 126.815 143.230 131.990 ;
        RECT 144.025 131.050 144.375 133.410 ;
        RECT 143.725 129.545 144.425 131.050 ;
        RECT 153.945 129.545 154.345 129.945 ;
        RECT 143.725 129.145 154.345 129.545 ;
        RECT 143.725 127.640 144.425 129.145 ;
        RECT 142.980 126.215 143.630 126.815 ;
        RECT 10.025 122.800 70.175 123.810 ;
        RECT 71.775 122.750 114.165 123.850 ;
        RECT 10.025 120.300 70.175 122.300 ;
        RECT 71.775 121.250 114.165 122.350 ;
        RECT 115.905 121.575 128.935 123.145 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 10.025 117.800 70.175 119.800 ;
        RECT 71.775 119.750 114.165 120.850 ;
        RECT 71.775 118.250 114.165 119.350 ;
        RECT 10.025 115.300 70.175 117.300 ;
        RECT 71.775 116.750 114.165 117.850 ;
        RECT 115.905 117.075 128.935 118.645 ;
        RECT 141.900 116.370 150.745 117.170 ;
        RECT 71.775 115.250 114.165 116.350 ;
        RECT 10.025 112.780 70.175 114.800 ;
        RECT 71.775 112.730 114.165 114.850 ;
        RECT 136.465 114.770 144.870 115.570 ;
        RECT 173.060 115.285 173.340 176.290 ;
        RECT 115.905 112.615 128.935 114.185 ;
        RECT 10.025 110.280 70.175 112.280 ;
        RECT 71.775 111.230 114.165 112.330 ;
        RECT 133.265 111.795 141.675 112.595 ;
        RECT 10.025 107.780 70.175 109.780 ;
        RECT 71.775 109.730 114.165 110.830 ;
        RECT 140.875 110.315 141.675 111.795 ;
        RECT 144.070 110.315 144.870 114.770 ;
        RECT 164.025 115.005 173.340 115.285 ;
        RECT 71.775 108.230 114.165 109.330 ;
        RECT 115.905 108.115 128.935 109.685 ;
        RECT 139.560 109.515 142.995 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 10.025 105.280 70.175 107.280 ;
        RECT 71.775 106.730 114.165 107.830 ;
        RECT 71.775 105.230 114.165 106.330 ;
        RECT 10.025 103.770 70.175 104.780 ;
        RECT 71.775 103.730 114.165 104.830 ;
        RECT 115.905 103.655 128.935 105.225 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 10.025 91.525 128.935 92.775 ;
        RECT 10.025 89.640 128.935 91.140 ;
        RECT 10.025 85.640 128.935 88.640 ;
        RECT 136.295 86.115 138.400 90.215 ;
        RECT 10.025 83.140 128.935 84.640 ;
        RECT 10.025 81.505 128.935 82.755 ;
        RECT 10.025 79.620 128.935 81.120 ;
        RECT 136.295 80.265 138.400 85.535 ;
        RECT 139.560 82.025 140.860 109.515 ;
        RECT 141.695 91.385 142.995 109.515 ;
        RECT 141.290 90.795 143.395 91.385 ;
        RECT 139.155 81.435 141.260 82.025 ;
        RECT 10.025 75.620 128.935 78.620 ;
        RECT 136.295 75.585 138.400 79.685 ;
        RECT 10.025 73.120 128.935 74.620 ;
        RECT 10.025 71.485 128.935 72.735 ;
        RECT 10.025 69.600 128.935 71.100 ;
        RECT 136.295 70.905 138.400 75.005 ;
        RECT 10.025 65.600 128.935 68.600 ;
        RECT 136.295 66.225 138.400 70.325 ;
        RECT 10.025 63.100 128.935 64.600 ;
        RECT 10.025 61.465 128.935 62.715 ;
        RECT 10.025 59.580 128.935 61.080 ;
        RECT 136.295 60.375 138.400 65.645 ;
        RECT 10.025 55.580 128.935 58.580 ;
        RECT 136.295 55.695 138.400 59.795 ;
        RECT 10.025 53.080 128.935 54.580 ;
        RECT 10.025 51.445 128.935 52.695 ;
        RECT 136.295 51.015 138.400 55.115 ;
        RECT 12.915 45.565 14.515 47.165 ;
        RECT 90.715 45.565 92.315 47.165 ;
        RECT 136.295 46.335 138.400 50.435 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 136.295 40.485 138.400 45.755 ;
        RECT 143.835 42.245 145.135 110.315 ;
        RECT 164.025 109.225 164.305 115.005 ;
        RECT 173.980 114.705 174.260 176.290 ;
        RECT 174.510 176.175 174.650 176.430 ;
        RECT 174.970 176.290 175.110 179.150 ;
        RECT 175.370 179.060 175.630 179.380 ;
        RECT 175.830 179.060 176.090 179.380 ;
        RECT 176.350 178.780 176.490 184.080 ;
        RECT 176.810 181.760 176.950 184.590 ;
        RECT 176.750 181.440 177.010 181.760 ;
        RECT 176.750 180.760 177.010 181.080 ;
        RECT 175.890 178.640 176.490 178.780 ;
        RECT 176.810 178.700 176.950 180.760 ;
        RECT 175.890 176.290 176.030 178.640 ;
        RECT 176.750 178.380 177.010 178.700 ;
        RECT 177.270 177.420 177.410 188.045 ;
        RECT 177.730 179.040 177.870 188.240 ;
        RECT 178.190 184.820 178.330 188.240 ;
        RECT 178.650 184.820 178.790 191.980 ;
        RECT 180.030 191.960 180.170 194.020 ;
        RECT 180.490 191.960 180.630 194.360 ;
        RECT 182.330 192.300 182.470 199.120 ;
        RECT 182.890 198.585 184.430 198.955 ;
        RECT 189.690 195.700 189.830 199.800 ;
        RECT 192.145 195.865 193.685 196.235 ;
        RECT 189.630 195.380 189.890 195.700 ;
        RECT 190.550 195.040 190.810 195.360 ;
        RECT 191.010 195.215 191.270 195.360 ;
        RECT 182.890 193.145 184.430 193.515 ;
        RECT 190.610 192.980 190.750 195.040 ;
        RECT 191.000 194.845 191.280 195.215 ;
        RECT 192.390 194.700 192.650 195.020 ;
        RECT 190.550 192.660 190.810 192.980 ;
        RECT 190.090 192.320 190.350 192.640 ;
        RECT 191.470 192.320 191.730 192.640 ;
        RECT 182.270 191.980 182.530 192.300 ;
        RECT 184.570 191.980 184.830 192.300 ;
        RECT 185.030 192.210 185.290 192.300 ;
        RECT 185.030 192.070 187.990 192.210 ;
        RECT 185.030 191.980 185.290 192.070 ;
        RECT 179.970 191.640 180.230 191.960 ;
        RECT 180.430 191.640 180.690 191.960 ;
        RECT 180.490 190.260 180.630 191.640 ;
        RECT 181.810 191.530 182.070 191.620 ;
        RECT 180.950 191.390 182.070 191.530 ;
        RECT 180.430 189.940 180.690 190.260 ;
        RECT 179.050 189.150 179.310 189.240 ;
        RECT 179.050 189.010 179.710 189.150 ;
        RECT 180.430 189.095 180.690 189.240 ;
        RECT 179.050 188.920 179.310 189.010 ;
        RECT 179.050 187.220 179.310 187.540 ;
        RECT 179.110 186.860 179.250 187.220 ;
        RECT 179.050 186.540 179.310 186.860 ;
        RECT 179.110 186.375 179.250 186.540 ;
        RECT 179.040 186.005 179.320 186.375 ;
        RECT 178.130 184.500 178.390 184.820 ;
        RECT 178.590 184.500 178.850 184.820 ;
        RECT 179.570 184.730 179.710 189.010 ;
        RECT 180.420 188.725 180.700 189.095 ;
        RECT 180.430 188.240 180.690 188.560 ;
        RECT 180.490 186.940 180.630 188.240 ;
        RECT 180.950 187.540 181.090 191.390 ;
        RECT 181.810 191.300 182.070 191.390 ;
        RECT 182.330 191.280 182.470 191.980 ;
        RECT 182.270 190.960 182.530 191.280 ;
        RECT 182.270 189.600 182.530 189.920 ;
        RECT 181.350 188.920 181.610 189.240 ;
        RECT 180.890 187.220 181.150 187.540 ;
        RECT 180.030 186.860 180.630 186.940 ;
        RECT 179.970 186.800 180.630 186.860 ;
        RECT 179.970 186.540 180.230 186.800 ;
        RECT 180.890 186.540 181.150 186.860 ;
        RECT 180.430 185.860 180.690 186.180 ;
        RECT 180.490 185.695 180.630 185.860 ;
        RECT 180.420 185.325 180.700 185.695 ;
        RECT 179.110 184.590 179.710 184.730 ;
        RECT 178.130 183.480 178.390 183.800 ;
        RECT 178.190 182.100 178.330 183.480 ;
        RECT 178.590 182.975 178.850 183.120 ;
        RECT 178.580 182.605 178.860 182.975 ;
        RECT 179.110 182.860 179.250 184.590 ;
        RECT 180.950 184.480 181.090 186.540 ;
        RECT 180.890 184.160 181.150 184.480 ;
        RECT 180.950 183.800 181.090 184.160 ;
        RECT 179.970 183.480 180.230 183.800 ;
        RECT 180.890 183.480 181.150 183.800 ;
        RECT 179.110 182.720 179.710 182.860 ;
        RECT 178.580 182.180 178.860 182.295 ;
        RECT 178.130 181.780 178.390 182.100 ;
        RECT 178.580 182.040 179.250 182.180 ;
        RECT 178.580 181.925 178.860 182.040 ;
        RECT 177.670 178.720 177.930 179.040 ;
        RECT 179.110 178.270 179.250 182.040 ;
        RECT 179.570 181.500 179.710 182.720 ;
        RECT 180.030 182.100 180.170 183.480 ;
        RECT 180.430 183.140 180.690 183.460 ;
        RECT 180.490 182.100 180.630 183.140 ;
        RECT 180.880 182.605 181.160 182.975 ;
        RECT 179.970 181.780 180.230 182.100 ;
        RECT 180.430 181.780 180.690 182.100 ;
        RECT 179.570 181.360 180.630 181.500 ;
        RECT 179.970 180.935 180.230 181.080 ;
        RECT 179.960 180.565 180.240 180.935 ;
        RECT 180.030 178.360 180.170 180.565 ;
        RECT 179.110 178.130 179.710 178.270 ;
        RECT 177.270 177.280 177.870 177.420 ;
        RECT 176.350 176.600 176.950 176.740 ;
        RECT 176.350 176.320 176.490 176.600 ;
        RECT 174.440 175.805 174.720 176.175 ;
        RECT 166.325 114.425 174.260 114.705 ;
        RECT 166.325 109.225 166.605 114.425 ;
        RECT 174.900 114.125 175.180 176.290 ;
        RECT 168.625 113.845 175.180 114.125 ;
        RECT 168.625 109.225 168.905 113.845 ;
        RECT 175.820 113.545 176.100 176.290 ;
        RECT 176.290 176.000 176.550 176.320 ;
        RECT 176.810 176.290 176.950 176.600 ;
        RECT 177.730 176.290 177.870 177.280 ;
        RECT 178.190 176.660 178.790 176.740 ;
        RECT 178.130 176.600 178.790 176.660 ;
        RECT 178.130 176.340 178.390 176.600 ;
        RECT 178.650 176.290 178.790 176.600 ;
        RECT 179.570 176.290 179.710 178.130 ;
        RECT 179.970 178.040 180.230 178.360 ;
        RECT 180.490 176.290 180.630 181.360 ;
        RECT 180.950 179.380 181.090 182.605 ;
        RECT 180.890 179.060 181.150 179.380 ;
        RECT 180.890 177.360 181.150 177.680 ;
        RECT 180.950 176.660 181.090 177.360 ;
        RECT 180.890 176.340 181.150 176.660 ;
        RECT 181.410 176.290 181.550 188.920 ;
        RECT 181.810 188.240 182.070 188.560 ;
        RECT 181.870 180.400 182.010 188.240 ;
        RECT 182.330 187.540 182.470 189.600 ;
        RECT 182.890 187.705 184.430 188.075 ;
        RECT 182.270 187.220 182.530 187.540 ;
        RECT 183.650 187.220 183.910 187.540 ;
        RECT 182.270 186.540 182.530 186.860 ;
        RECT 182.330 185.015 182.470 186.540 ;
        RECT 182.730 185.520 182.990 185.840 ;
        RECT 183.190 185.520 183.450 185.840 ;
        RECT 182.260 184.645 182.540 185.015 ;
        RECT 182.270 183.710 182.530 183.800 ;
        RECT 182.790 183.710 182.930 185.520 ;
        RECT 182.270 183.570 182.930 183.710 ;
        RECT 182.270 183.480 182.530 183.570 ;
        RECT 182.330 181.420 182.470 183.480 ;
        RECT 183.250 183.120 183.390 185.520 ;
        RECT 183.710 184.820 183.850 187.220 ;
        RECT 184.630 187.200 184.770 191.980 ;
        RECT 185.030 188.920 185.290 189.240 ;
        RECT 185.490 188.920 185.750 189.240 ;
        RECT 187.330 188.920 187.590 189.240 ;
        RECT 184.570 186.880 184.830 187.200 ;
        RECT 184.560 186.260 184.840 186.375 ;
        RECT 184.170 186.120 184.840 186.260 ;
        RECT 183.650 184.500 183.910 184.820 ;
        RECT 184.170 184.480 184.310 186.120 ;
        RECT 184.560 186.005 184.840 186.120 ;
        RECT 184.570 185.520 184.830 185.840 ;
        RECT 184.110 184.160 184.370 184.480 ;
        RECT 183.190 182.800 183.450 183.120 ;
        RECT 182.890 182.265 184.430 182.635 ;
        RECT 184.110 181.440 184.370 181.760 ;
        RECT 182.270 181.100 182.530 181.420 ;
        RECT 181.810 180.080 182.070 180.400 ;
        RECT 181.810 178.950 182.070 179.040 ;
        RECT 182.330 178.950 182.470 181.100 ;
        RECT 182.720 180.565 183.000 180.935 ;
        RECT 181.810 178.810 182.470 178.950 ;
        RECT 181.810 178.720 182.070 178.810 ;
        RECT 182.790 178.700 182.930 180.565 ;
        RECT 183.640 179.885 183.920 180.255 ;
        RECT 182.730 178.380 182.990 178.700 ;
        RECT 181.810 178.040 182.070 178.360 ;
        RECT 181.870 176.320 182.010 178.040 ;
        RECT 182.270 177.700 182.530 178.020 ;
        RECT 170.925 113.265 176.100 113.545 ;
        RECT 170.925 109.225 171.205 113.265 ;
        RECT 176.740 112.965 177.020 176.290 ;
        RECT 173.225 112.685 177.020 112.965 ;
        RECT 173.225 109.225 173.505 112.685 ;
        RECT 177.660 112.385 177.940 176.290 ;
        RECT 175.525 112.105 177.940 112.385 ;
        RECT 175.525 109.225 175.805 112.105 ;
        RECT 178.580 111.805 178.860 176.290 ;
        RECT 177.825 111.525 178.860 111.805 ;
        RECT 179.500 111.805 179.780 176.290 ;
        RECT 180.420 112.385 180.700 176.290 ;
        RECT 181.340 112.965 181.620 176.290 ;
        RECT 181.810 176.000 182.070 176.320 ;
        RECT 182.330 176.290 182.470 177.700 ;
        RECT 183.710 177.590 183.850 179.885 ;
        RECT 184.170 178.270 184.310 181.440 ;
        RECT 184.630 179.380 184.770 185.520 ;
        RECT 185.090 181.760 185.230 188.920 ;
        RECT 185.030 181.440 185.290 181.760 ;
        RECT 185.030 180.760 185.290 181.080 ;
        RECT 185.090 179.380 185.230 180.760 ;
        RECT 184.570 179.060 184.830 179.380 ;
        RECT 185.030 179.060 185.290 179.380 ;
        RECT 184.570 178.270 184.830 178.360 ;
        RECT 184.170 178.130 184.830 178.270 ;
        RECT 184.570 178.040 184.830 178.130 ;
        RECT 185.550 177.930 185.690 188.920 ;
        RECT 185.950 188.580 186.210 188.900 ;
        RECT 186.010 182.100 186.150 188.580 ;
        RECT 186.410 188.240 186.670 188.560 ;
        RECT 186.470 186.520 186.610 188.240 ;
        RECT 187.390 188.160 187.530 188.920 ;
        RECT 186.930 188.020 187.530 188.160 ;
        RECT 186.410 186.200 186.670 186.520 ;
        RECT 186.410 185.520 186.670 185.840 ;
        RECT 186.470 182.100 186.610 185.520 ;
        RECT 185.950 181.780 186.210 182.100 ;
        RECT 186.410 181.780 186.670 182.100 ;
        RECT 186.410 181.100 186.670 181.420 ;
        RECT 185.940 179.885 186.220 180.255 ;
        RECT 185.090 177.790 185.690 177.930 ;
        RECT 183.710 177.450 184.770 177.590 ;
        RECT 182.890 176.825 184.430 177.195 ;
        RECT 183.650 176.570 183.910 176.660 ;
        RECT 184.630 176.570 184.770 177.450 ;
        RECT 183.250 176.430 183.910 176.570 ;
        RECT 183.250 176.290 183.390 176.430 ;
        RECT 183.650 176.340 183.910 176.430 ;
        RECT 184.170 176.430 184.770 176.570 ;
        RECT 184.170 176.290 184.310 176.430 ;
        RECT 185.090 176.290 185.230 177.790 ;
        RECT 186.010 176.290 186.150 179.885 ;
        RECT 186.470 178.700 186.610 181.100 ;
        RECT 186.410 178.380 186.670 178.700 ;
        RECT 186.410 177.700 186.670 178.020 ;
        RECT 186.470 176.660 186.610 177.700 ;
        RECT 186.410 176.340 186.670 176.660 ;
        RECT 186.930 176.290 187.070 188.020 ;
        RECT 187.850 187.200 187.990 192.070 ;
        RECT 188.710 190.960 188.970 191.280 ;
        RECT 188.770 190.260 188.910 190.960 ;
        RECT 188.710 189.940 188.970 190.260 ;
        RECT 190.150 189.240 190.290 192.320 ;
        RECT 191.010 191.980 191.270 192.300 ;
        RECT 189.630 189.150 189.890 189.240 ;
        RECT 188.770 189.010 189.890 189.150 ;
        RECT 188.250 188.240 188.510 188.560 ;
        RECT 187.330 186.880 187.590 187.200 ;
        RECT 187.790 186.880 188.050 187.200 ;
        RECT 187.390 183.540 187.530 186.880 ;
        RECT 188.310 185.015 188.450 188.240 ;
        RECT 188.240 184.645 188.520 185.015 ;
        RECT 187.780 183.965 188.060 184.335 ;
        RECT 187.790 183.820 188.050 183.965 ;
        RECT 187.390 183.400 188.450 183.540 ;
        RECT 187.330 183.030 187.590 183.120 ;
        RECT 187.330 182.890 187.990 183.030 ;
        RECT 187.330 182.800 187.590 182.890 ;
        RECT 187.850 176.290 187.990 182.890 ;
        RECT 188.310 177.590 188.450 183.400 ;
        RECT 188.770 178.215 188.910 189.010 ;
        RECT 189.630 188.920 189.890 189.010 ;
        RECT 190.090 188.920 190.350 189.240 ;
        RECT 189.170 186.880 189.430 187.200 ;
        RECT 189.230 182.100 189.370 186.880 ;
        RECT 190.150 186.860 190.290 188.920 ;
        RECT 191.070 188.560 191.210 191.980 ;
        RECT 191.530 189.240 191.670 192.320 ;
        RECT 192.450 192.300 192.590 194.700 ;
        RECT 195.150 194.420 195.410 194.680 ;
        RECT 195.150 194.360 196.270 194.420 ;
        RECT 195.210 194.280 196.270 194.360 ;
        RECT 196.130 194.000 196.270 194.280 ;
        RECT 194.690 193.680 194.950 194.000 ;
        RECT 196.070 193.680 196.330 194.000 ;
        RECT 194.750 192.300 194.890 193.680 ;
        RECT 192.390 191.980 192.650 192.300 ;
        RECT 194.690 191.980 194.950 192.300 ;
        RECT 196.130 191.960 196.270 193.680 ;
        RECT 199.350 192.980 199.490 199.800 ;
        RECT 201.400 198.585 202.940 198.955 ;
        RECT 207.570 194.020 207.830 194.340 ;
        RECT 201.400 193.145 202.940 193.515 ;
        RECT 199.290 192.660 199.550 192.980 ;
        RECT 200.670 192.320 200.930 192.640 ;
        RECT 196.070 191.640 196.330 191.960 ;
        RECT 192.145 190.425 193.685 190.795 ;
        RECT 196.130 190.030 197.190 190.170 ;
        RECT 191.470 188.920 191.730 189.240 ;
        RECT 191.930 188.920 192.190 189.240 ;
        RECT 193.310 188.920 193.570 189.240 ;
        RECT 191.010 188.240 191.270 188.560 ;
        RECT 190.540 187.365 190.820 187.735 ;
        RECT 190.550 187.220 190.810 187.365 ;
        RECT 191.070 186.860 191.210 188.240 ;
        RECT 191.530 187.200 191.670 188.920 ;
        RECT 191.990 188.415 192.130 188.920 ;
        RECT 193.370 188.560 193.510 188.920 ;
        RECT 195.150 188.580 195.410 188.900 ;
        RECT 195.610 188.580 195.870 188.900 ;
        RECT 191.920 188.045 192.200 188.415 ;
        RECT 193.310 188.240 193.570 188.560 ;
        RECT 193.770 188.300 194.030 188.560 ;
        RECT 193.770 188.240 194.890 188.300 ;
        RECT 191.930 187.220 192.190 187.540 ;
        RECT 191.470 186.880 191.730 187.200 ;
        RECT 190.090 186.540 190.350 186.860 ;
        RECT 191.010 186.540 191.270 186.860 ;
        RECT 189.630 186.200 189.890 186.520 ;
        RECT 189.690 182.860 189.830 186.200 ;
        RECT 190.150 183.800 190.290 186.540 ;
        RECT 190.550 186.200 190.810 186.520 ;
        RECT 190.610 185.695 190.750 186.200 ;
        RECT 191.990 185.750 192.130 187.220 ;
        RECT 193.370 186.180 193.510 188.240 ;
        RECT 193.830 188.160 194.890 188.240 ;
        RECT 193.830 186.860 194.430 186.940 ;
        RECT 193.770 186.800 194.430 186.860 ;
        RECT 193.770 186.540 194.030 186.800 ;
        RECT 193.310 185.860 193.570 186.180 ;
        RECT 190.540 185.325 190.820 185.695 ;
        RECT 191.070 185.610 192.130 185.750 ;
        RECT 191.070 184.900 191.210 185.610 ;
        RECT 190.610 184.760 191.210 184.900 ;
        RECT 190.610 184.480 190.750 184.760 ;
        RECT 191.460 184.645 191.740 185.015 ;
        RECT 192.145 184.985 193.685 185.355 ;
        RECT 191.470 184.500 191.730 184.645 ;
        RECT 190.550 184.160 190.810 184.480 ;
        RECT 192.390 183.820 192.650 184.140 ;
        RECT 190.090 183.480 190.350 183.800 ;
        RECT 191.930 183.140 192.190 183.460 ;
        RECT 189.690 182.720 190.750 182.860 ;
        RECT 191.010 182.800 191.270 183.120 ;
        RECT 191.470 182.800 191.730 183.120 ;
        RECT 189.170 181.780 189.430 182.100 ;
        RECT 190.080 181.925 190.360 182.295 ;
        RECT 189.170 180.760 189.430 181.080 ;
        RECT 190.150 180.820 190.290 181.925 ;
        RECT 189.230 179.380 189.370 180.760 ;
        RECT 189.690 180.680 190.290 180.820 ;
        RECT 189.690 179.380 189.830 180.680 ;
        RECT 190.090 180.080 190.350 180.400 ;
        RECT 189.170 179.060 189.430 179.380 ;
        RECT 189.630 179.060 189.890 179.380 ;
        RECT 190.150 178.700 190.290 180.080 ;
        RECT 190.090 178.380 190.350 178.700 ;
        RECT 188.700 177.845 188.980 178.215 ;
        RECT 189.630 178.040 189.890 178.360 ;
        RECT 188.310 177.450 189.370 177.590 ;
        RECT 189.690 177.535 189.830 178.040 ;
        RECT 188.700 176.485 188.980 176.855 ;
        RECT 189.230 176.740 189.370 177.450 ;
        RECT 189.620 177.165 189.900 177.535 ;
        RECT 190.090 177.360 190.350 177.680 ;
        RECT 189.230 176.600 189.830 176.740 ;
        RECT 190.150 176.660 190.290 177.360 ;
        RECT 188.770 176.290 188.910 176.485 ;
        RECT 189.690 176.290 189.830 176.600 ;
        RECT 190.090 176.340 190.350 176.660 ;
        RECT 190.610 176.290 190.750 182.720 ;
        RECT 191.070 178.215 191.210 182.800 ;
        RECT 191.530 179.380 191.670 182.800 ;
        RECT 191.990 180.400 192.130 183.140 ;
        RECT 192.450 180.740 192.590 183.820 ;
        RECT 193.770 181.440 194.030 181.760 ;
        RECT 192.390 180.420 192.650 180.740 ;
        RECT 191.930 180.080 192.190 180.400 ;
        RECT 192.145 179.545 193.685 179.915 ;
        RECT 193.830 179.380 193.970 181.440 ;
        RECT 194.290 179.380 194.430 186.800 ;
        RECT 194.750 182.100 194.890 188.160 ;
        RECT 195.210 187.200 195.350 188.580 ;
        RECT 195.150 186.880 195.410 187.200 ;
        RECT 195.140 184.645 195.420 185.015 ;
        RECT 195.670 184.820 195.810 188.580 ;
        RECT 195.210 183.800 195.350 184.645 ;
        RECT 195.610 184.500 195.870 184.820 ;
        RECT 195.150 183.480 195.410 183.800 ;
        RECT 194.690 181.780 194.950 182.100 ;
        RECT 196.130 182.010 196.270 190.030 ;
        RECT 196.520 189.405 196.800 189.775 ;
        RECT 196.590 187.540 196.730 189.405 ;
        RECT 197.050 189.150 197.190 190.030 ;
        RECT 197.450 189.150 197.710 189.240 ;
        RECT 197.050 189.010 197.710 189.150 ;
        RECT 197.450 188.920 197.710 189.010 ;
        RECT 199.750 188.240 200.010 188.560 ;
        RECT 196.530 187.220 196.790 187.540 ;
        RECT 197.050 187.310 198.570 187.450 ;
        RECT 197.050 184.730 197.190 187.310 ;
        RECT 198.430 186.860 198.570 187.310 ;
        RECT 197.450 186.540 197.710 186.860 ;
        RECT 197.910 186.540 198.170 186.860 ;
        RECT 198.370 186.540 198.630 186.860 ;
        RECT 196.590 184.590 197.190 184.730 ;
        RECT 196.590 184.140 196.730 184.590 ;
        RECT 196.530 183.820 196.790 184.140 ;
        RECT 196.520 183.285 196.800 183.655 ;
        RECT 196.990 183.480 197.250 183.800 ;
        RECT 196.530 183.140 196.790 183.285 ;
        RECT 195.210 181.870 196.270 182.010 ;
        RECT 194.690 180.420 194.950 180.740 ;
        RECT 191.470 179.060 191.730 179.380 ;
        RECT 193.770 179.060 194.030 179.380 ;
        RECT 194.230 179.060 194.490 179.380 ;
        RECT 194.750 179.040 194.890 180.420 ;
        RECT 194.690 178.720 194.950 179.040 ;
        RECT 193.310 178.380 193.570 178.700 ;
        RECT 191.000 177.845 191.280 178.215 ;
        RECT 191.930 178.040 192.190 178.360 ;
        RECT 191.070 176.600 191.670 176.740 ;
        RECT 182.260 113.545 182.540 176.290 ;
        RECT 183.180 114.125 183.460 176.290 ;
        RECT 184.100 114.705 184.380 176.290 ;
        RECT 185.020 115.285 185.300 176.290 ;
        RECT 185.940 115.865 186.220 176.290 ;
        RECT 186.860 116.445 187.140 176.290 ;
        RECT 187.780 117.025 188.060 176.290 ;
        RECT 188.700 117.605 188.980 176.290 ;
        RECT 189.620 118.185 189.900 176.290 ;
        RECT 190.540 118.765 190.820 176.290 ;
        RECT 191.070 175.640 191.210 176.600 ;
        RECT 191.530 176.290 191.670 176.600 ;
        RECT 191.010 175.320 191.270 175.640 ;
        RECT 191.460 119.345 191.740 176.290 ;
        RECT 191.990 175.980 192.130 178.040 ;
        RECT 192.450 176.430 193.050 176.570 ;
        RECT 192.450 176.290 192.590 176.430 ;
        RECT 191.930 175.660 192.190 175.980 ;
        RECT 192.380 119.925 192.660 176.290 ;
        RECT 192.910 175.495 193.050 176.430 ;
        RECT 193.370 176.290 193.510 178.380 ;
        RECT 194.230 178.270 194.490 178.360 ;
        RECT 194.230 178.130 194.890 178.270 ;
        RECT 194.230 178.040 194.490 178.130 ;
        RECT 193.830 176.600 194.430 176.740 ;
        RECT 193.830 176.320 193.970 176.600 ;
        RECT 192.840 175.125 193.120 175.495 ;
        RECT 193.300 120.505 193.580 176.290 ;
        RECT 193.770 176.000 194.030 176.320 ;
        RECT 194.290 176.290 194.430 176.600 ;
        RECT 194.750 176.320 194.890 178.130 ;
        RECT 194.220 121.085 194.500 176.290 ;
        RECT 194.690 176.000 194.950 176.320 ;
        RECT 195.210 176.290 195.350 181.870 ;
        RECT 197.050 181.080 197.190 183.480 ;
        RECT 197.510 182.100 197.650 186.540 ;
        RECT 197.970 184.820 198.110 186.540 ;
        RECT 198.830 185.860 199.090 186.180 ;
        RECT 199.280 186.005 199.560 186.375 ;
        RECT 199.290 185.860 199.550 186.005 ;
        RECT 198.370 185.520 198.630 185.840 ;
        RECT 197.910 184.500 198.170 184.820 ;
        RECT 197.910 182.800 198.170 183.120 ;
        RECT 197.450 181.780 197.710 182.100 ;
        RECT 197.440 181.500 197.720 181.615 ;
        RECT 197.970 181.500 198.110 182.800 ;
        RECT 198.430 182.100 198.570 185.520 ;
        RECT 198.370 181.780 198.630 182.100 ;
        RECT 197.440 181.360 198.110 181.500 ;
        RECT 198.890 181.420 199.030 185.860 ;
        RECT 199.810 184.335 199.950 188.240 ;
        RECT 200.200 187.365 200.480 187.735 ;
        RECT 200.270 186.180 200.410 187.365 ;
        RECT 200.210 185.860 200.470 186.180 ;
        RECT 199.740 183.965 200.020 184.335 ;
        RECT 200.210 183.710 200.470 183.800 ;
        RECT 199.810 183.570 200.470 183.710 ;
        RECT 199.290 183.140 199.550 183.460 ;
        RECT 197.440 181.245 197.720 181.360 ;
        RECT 198.370 181.100 198.630 181.420 ;
        RECT 198.830 181.100 199.090 181.420 ;
        RECT 196.990 180.760 197.250 181.080 ;
        RECT 198.430 180.935 198.570 181.100 ;
        RECT 199.350 181.080 199.490 183.140 ;
        RECT 198.360 180.565 198.640 180.935 ;
        RECT 199.290 180.760 199.550 181.080 ;
        RECT 199.350 179.380 199.490 180.760 ;
        RECT 199.290 179.060 199.550 179.380 ;
        RECT 195.610 178.720 195.870 179.040 ;
        RECT 197.450 178.720 197.710 179.040 ;
        RECT 195.670 178.360 195.810 178.720 ;
        RECT 195.610 178.040 195.870 178.360 ;
        RECT 196.990 177.360 197.250 177.680 ;
        RECT 195.670 176.660 196.270 176.740 ;
        RECT 195.610 176.600 196.270 176.660 ;
        RECT 195.610 176.340 195.870 176.600 ;
        RECT 196.130 176.290 196.270 176.600 ;
        RECT 197.050 176.290 197.190 177.360 ;
        RECT 195.140 121.665 195.420 176.290 ;
        RECT 196.060 122.245 196.340 176.290 ;
        RECT 196.980 122.825 197.260 176.290 ;
        RECT 197.510 175.640 197.650 178.720 ;
        RECT 199.280 177.845 199.560 178.215 ;
        RECT 199.290 177.700 199.550 177.845 ;
        RECT 197.900 177.165 198.180 177.535 ;
        RECT 199.810 177.420 199.950 183.570 ;
        RECT 200.210 183.480 200.470 183.570 ;
        RECT 200.210 182.800 200.470 183.120 ;
        RECT 200.270 182.100 200.410 182.800 ;
        RECT 200.730 182.100 200.870 192.320 ;
        RECT 204.350 190.960 204.610 191.280 ;
        RECT 201.400 187.705 202.940 188.075 ;
        RECT 202.050 186.540 202.310 186.860 ;
        RECT 202.110 185.015 202.250 186.540 ;
        RECT 202.040 184.645 202.320 185.015 ;
        RECT 203.890 183.820 204.150 184.140 ;
        RECT 203.430 183.480 203.690 183.800 ;
        RECT 201.400 182.265 202.940 182.635 ;
        RECT 200.210 181.780 200.470 182.100 ;
        RECT 200.670 181.780 200.930 182.100 ;
        RECT 202.960 180.565 203.240 180.935 ;
        RECT 203.030 179.380 203.170 180.565 ;
        RECT 202.970 179.060 203.230 179.380 ;
        RECT 203.490 179.290 203.630 183.480 ;
        RECT 203.950 181.080 204.090 183.820 ;
        RECT 203.890 180.760 204.150 181.080 ;
        RECT 204.410 179.380 204.550 190.960 ;
        RECT 207.630 184.820 207.770 194.020 ;
        RECT 209.010 190.260 209.150 199.800 ;
        RECT 217.230 199.460 217.490 199.780 ;
        RECT 210.655 195.865 212.195 196.235 ;
        RECT 209.870 190.960 210.130 191.280 ;
        RECT 208.950 189.940 209.210 190.260 ;
        RECT 209.930 189.580 210.070 190.960 ;
        RECT 210.655 190.425 212.195 190.795 ;
        RECT 209.870 189.260 210.130 189.580 ;
        RECT 210.330 189.095 210.590 189.240 ;
        RECT 210.320 188.725 210.600 189.095 ;
        RECT 217.290 187.540 217.430 199.460 ;
        RECT 219.910 198.585 221.450 198.955 ;
        RECT 219.910 193.145 221.450 193.515 ;
        RECT 226.950 190.260 227.090 199.800 ;
        RECT 229.165 195.865 230.705 196.235 ;
        RECT 229.165 190.425 230.705 190.795 ;
        RECT 226.890 189.940 227.150 190.260 ;
        RECT 225.970 189.600 226.230 189.920 ;
        RECT 221.830 188.240 222.090 188.560 ;
        RECT 219.910 187.705 221.450 188.075 ;
        RECT 216.770 187.220 217.030 187.540 ;
        RECT 217.230 187.220 217.490 187.540 ;
        RECT 219.070 187.220 219.330 187.540 ;
        RECT 208.020 186.685 208.300 187.055 ;
        RECT 209.870 186.770 210.130 186.860 ;
        RECT 208.090 186.520 208.230 186.685 ;
        RECT 209.470 186.630 210.130 186.770 ;
        RECT 212.160 186.685 212.440 187.055 ;
        RECT 213.550 186.770 213.810 186.860 ;
        RECT 214.930 186.770 215.190 186.860 ;
        RECT 208.030 186.200 208.290 186.520 ;
        RECT 207.570 184.500 207.830 184.820 ;
        RECT 206.190 183.480 206.450 183.800 ;
        RECT 206.250 182.100 206.390 183.480 ;
        RECT 206.650 183.030 206.910 183.120 ;
        RECT 206.650 182.890 207.770 183.030 ;
        RECT 206.650 182.800 206.910 182.890 ;
        RECT 206.190 181.780 206.450 182.100 ;
        RECT 205.730 181.330 205.990 181.420 ;
        RECT 205.330 181.190 205.990 181.330 ;
        RECT 203.490 179.150 204.090 179.290 ;
        RECT 200.670 178.040 200.930 178.360 ;
        RECT 202.510 178.270 202.770 178.360 ;
        RECT 202.510 178.130 203.630 178.270 ;
        RECT 202.510 178.040 202.770 178.130 ;
        RECT 199.810 177.280 200.410 177.420 ;
        RECT 197.970 176.290 198.110 177.165 ;
        RECT 198.430 176.600 199.030 176.740 ;
        RECT 197.450 175.320 197.710 175.640 ;
        RECT 197.900 123.405 198.180 176.290 ;
        RECT 198.430 175.980 198.570 176.600 ;
        RECT 198.890 176.290 199.030 176.600 ;
        RECT 199.350 176.600 199.950 176.740 ;
        RECT 200.270 176.660 200.410 177.280 ;
        RECT 199.350 176.320 199.490 176.600 ;
        RECT 198.370 175.660 198.630 175.980 ;
        RECT 198.820 123.985 199.100 176.290 ;
        RECT 199.290 176.000 199.550 176.320 ;
        RECT 199.810 176.290 199.950 176.600 ;
        RECT 200.210 176.340 200.470 176.660 ;
        RECT 200.730 176.290 200.870 178.040 ;
        RECT 201.400 176.825 202.940 177.195 ;
        RECT 201.130 176.570 201.390 176.660 ;
        RECT 202.970 176.570 203.230 176.660 ;
        RECT 201.130 176.430 201.790 176.570 ;
        RECT 201.130 176.340 201.390 176.430 ;
        RECT 201.650 176.290 201.790 176.430 ;
        RECT 202.570 176.430 203.230 176.570 ;
        RECT 202.570 176.290 202.710 176.430 ;
        RECT 202.970 176.340 203.230 176.430 ;
        RECT 203.490 176.290 203.630 178.130 ;
        RECT 203.950 176.660 204.090 179.150 ;
        RECT 204.350 179.060 204.610 179.380 ;
        RECT 204.810 178.270 205.070 178.360 ;
        RECT 204.410 178.130 205.070 178.270 ;
        RECT 203.890 176.340 204.150 176.660 ;
        RECT 204.410 176.290 204.550 178.130 ;
        RECT 204.810 178.040 205.070 178.130 ;
        RECT 205.330 176.290 205.470 181.190 ;
        RECT 205.730 181.100 205.990 181.190 ;
        RECT 207.630 180.400 207.770 182.890 ;
        RECT 206.650 180.080 206.910 180.400 ;
        RECT 207.110 180.080 207.370 180.400 ;
        RECT 207.570 180.080 207.830 180.400 ;
        RECT 206.710 178.700 206.850 180.080 ;
        RECT 206.650 178.380 206.910 178.700 ;
        RECT 207.170 178.215 207.310 180.080 ;
        RECT 208.090 179.460 208.230 186.200 ;
        RECT 208.950 181.780 209.210 182.100 ;
        RECT 208.480 179.460 208.760 179.575 ;
        RECT 208.090 179.320 208.760 179.460 ;
        RECT 208.480 179.205 208.760 179.320 ;
        RECT 206.190 177.700 206.450 178.020 ;
        RECT 207.100 177.845 207.380 178.215 ;
        RECT 206.250 176.290 206.390 177.700 ;
        RECT 208.020 177.165 208.300 177.535 ;
        RECT 207.100 176.485 207.380 176.855 ;
        RECT 207.170 176.290 207.310 176.485 ;
        RECT 208.090 176.290 208.230 177.165 ;
        RECT 209.010 176.290 209.150 181.780 ;
        RECT 209.470 178.950 209.610 186.630 ;
        RECT 209.870 186.540 210.130 186.630 ;
        RECT 212.170 186.540 212.430 186.685 ;
        RECT 213.550 186.630 214.210 186.770 ;
        RECT 213.550 186.540 213.810 186.630 ;
        RECT 213.090 186.200 213.350 186.520 ;
        RECT 209.870 185.860 210.130 186.180 ;
        RECT 209.930 184.140 210.070 185.860 ;
        RECT 210.655 184.985 212.195 185.355 ;
        RECT 209.870 184.050 210.130 184.140 ;
        RECT 209.870 183.910 210.530 184.050 ;
        RECT 209.870 183.820 210.130 183.910 ;
        RECT 210.390 181.420 210.530 183.910 ;
        RECT 211.710 183.655 211.970 183.800 ;
        RECT 211.700 183.285 211.980 183.655 ;
        RECT 213.150 183.370 213.290 186.200 ;
        RECT 213.540 184.645 213.820 185.015 ;
        RECT 213.610 184.480 213.750 184.645 ;
        RECT 213.550 184.160 213.810 184.480 ;
        RECT 213.150 183.230 213.750 183.370 ;
        RECT 213.610 182.295 213.750 183.230 ;
        RECT 210.790 181.780 211.050 182.100 ;
        RECT 213.540 181.925 213.820 182.295 ;
        RECT 210.850 181.420 210.990 181.780 ;
        RECT 210.330 181.100 210.590 181.420 ;
        RECT 210.790 181.100 211.050 181.420 ;
        RECT 211.710 181.100 211.970 181.420 ;
        RECT 211.770 180.935 211.910 181.100 ;
        RECT 213.550 180.990 213.810 181.080 ;
        RECT 211.700 180.565 211.980 180.935 ;
        RECT 212.690 180.850 213.810 180.990 ;
        RECT 211.710 180.310 211.970 180.400 ;
        RECT 212.690 180.310 212.830 180.850 ;
        RECT 213.550 180.760 213.810 180.850 ;
        RECT 211.710 180.170 212.830 180.310 ;
        RECT 211.710 180.080 211.970 180.170 ;
        RECT 213.550 180.080 213.810 180.400 ;
        RECT 209.860 179.460 210.140 179.575 ;
        RECT 210.655 179.545 212.195 179.915 ;
        RECT 209.860 179.320 210.530 179.460 ;
        RECT 209.860 179.205 210.140 179.320 ;
        RECT 209.470 178.810 210.070 178.950 ;
        RECT 209.930 176.290 210.070 178.810 ;
        RECT 210.390 178.360 210.530 179.320 ;
        RECT 212.620 179.290 212.900 179.575 ;
        RECT 210.850 179.205 212.900 179.290 ;
        RECT 210.850 179.150 212.830 179.205 ;
        RECT 210.330 178.040 210.590 178.360 ;
        RECT 210.330 177.360 210.590 177.680 ;
        RECT 210.390 176.660 210.530 177.360 ;
        RECT 210.330 176.340 210.590 176.660 ;
        RECT 210.850 176.290 210.990 179.150 ;
        RECT 211.700 178.525 211.980 178.895 ;
        RECT 213.610 178.700 213.750 180.080 ;
        RECT 211.770 178.360 211.910 178.525 ;
        RECT 213.550 178.380 213.810 178.700 ;
        RECT 211.250 178.040 211.510 178.360 ;
        RECT 211.710 178.040 211.970 178.360 ;
        RECT 211.310 176.660 211.450 178.040 ;
        RECT 214.070 177.680 214.210 186.630 ;
        RECT 214.930 186.630 215.590 186.770 ;
        RECT 214.930 186.540 215.190 186.630 ;
        RECT 214.930 185.520 215.190 185.840 ;
        RECT 214.990 184.820 215.130 185.520 ;
        RECT 214.930 184.500 215.190 184.820 ;
        RECT 214.470 184.220 214.730 184.480 ;
        RECT 214.920 184.220 215.200 184.335 ;
        RECT 214.470 184.160 215.200 184.220 ;
        RECT 214.530 184.080 215.200 184.160 ;
        RECT 214.920 183.965 215.200 184.080 ;
        RECT 214.930 183.710 215.190 183.800 ;
        RECT 214.530 183.570 215.190 183.710 ;
        RECT 211.710 177.360 211.970 177.680 ;
        RECT 214.010 177.360 214.270 177.680 ;
        RECT 211.250 176.340 211.510 176.660 ;
        RECT 211.770 176.290 211.910 177.360 ;
        RECT 214.010 176.570 214.270 176.660 ;
        RECT 212.230 176.430 212.830 176.570 ;
        RECT 199.740 124.565 200.020 176.290 ;
        RECT 200.660 125.145 200.940 176.290 ;
        RECT 201.580 125.725 201.860 176.290 ;
        RECT 202.500 126.305 202.780 176.290 ;
        RECT 203.420 126.885 203.700 176.290 ;
        RECT 204.340 127.465 204.620 176.290 ;
        RECT 205.260 128.045 205.540 176.290 ;
        RECT 206.180 128.625 206.460 176.290 ;
        RECT 207.100 129.205 207.380 176.290 ;
        RECT 208.020 129.785 208.300 176.290 ;
        RECT 208.940 130.365 209.220 176.290 ;
        RECT 209.860 130.945 210.140 176.290 ;
        RECT 210.780 131.525 211.060 176.290 ;
        RECT 211.700 132.105 211.980 176.290 ;
        RECT 212.230 176.175 212.370 176.430 ;
        RECT 212.690 176.290 212.830 176.430 ;
        RECT 213.610 176.430 214.270 176.570 ;
        RECT 213.610 176.290 213.750 176.430 ;
        RECT 214.010 176.340 214.270 176.430 ;
        RECT 214.530 176.290 214.670 183.570 ;
        RECT 214.930 183.480 215.190 183.570 ;
        RECT 214.930 180.760 215.190 181.080 ;
        RECT 214.990 180.400 215.130 180.760 ;
        RECT 214.930 180.080 215.190 180.400 ;
        RECT 215.450 178.610 215.590 186.630 ;
        RECT 215.850 185.695 216.110 185.840 ;
        RECT 215.840 185.325 216.120 185.695 ;
        RECT 215.850 183.480 216.110 183.800 ;
        RECT 215.910 181.615 216.050 183.480 ;
        RECT 216.310 182.800 216.570 183.120 ;
        RECT 215.840 181.245 216.120 181.615 ;
        RECT 215.850 180.935 216.110 181.080 ;
        RECT 215.840 180.565 216.120 180.935 ;
        RECT 215.840 179.885 216.120 180.255 ;
        RECT 215.910 179.380 216.050 179.885 ;
        RECT 215.850 179.060 216.110 179.380 ;
        RECT 214.990 178.470 215.590 178.610 ;
        RECT 214.990 176.660 215.130 178.470 ;
        RECT 216.370 178.360 216.510 182.800 ;
        RECT 216.830 182.100 216.970 187.220 ;
        RECT 217.230 185.860 217.490 186.180 ;
        RECT 217.290 182.100 217.430 185.860 ;
        RECT 218.610 184.160 218.870 184.480 ;
        RECT 218.150 183.480 218.410 183.800 ;
        RECT 217.690 182.800 217.950 183.120 ;
        RECT 218.210 182.975 218.350 183.480 ;
        RECT 216.770 181.780 217.030 182.100 ;
        RECT 217.230 181.780 217.490 182.100 ;
        RECT 217.750 181.330 217.890 182.800 ;
        RECT 218.140 182.605 218.420 182.975 ;
        RECT 218.670 182.180 218.810 184.160 ;
        RECT 216.830 181.190 217.890 181.330 ;
        RECT 218.210 182.040 218.810 182.180 ;
        RECT 216.310 178.040 216.570 178.360 ;
        RECT 215.390 177.700 215.650 178.020 ;
        RECT 215.450 177.535 215.590 177.700 ;
        RECT 215.380 177.165 215.660 177.535 ;
        RECT 216.830 177.420 216.970 181.190 ;
        RECT 217.690 180.080 217.950 180.400 ;
        RECT 217.230 178.040 217.490 178.360 ;
        RECT 217.750 178.215 217.890 180.080 ;
        RECT 217.290 177.535 217.430 178.040 ;
        RECT 217.680 177.845 217.960 178.215 ;
        RECT 218.210 177.590 218.350 182.040 ;
        RECT 218.610 181.440 218.870 181.760 ;
        RECT 218.670 179.040 218.810 181.440 ;
        RECT 219.130 180.935 219.270 187.220 ;
        RECT 221.890 186.860 222.030 188.240 ;
        RECT 226.030 188.160 226.170 189.600 ;
        RECT 226.890 189.260 227.150 189.580 ;
        RECT 227.340 189.405 227.620 189.775 ;
        RECT 230.630 189.520 232.610 189.660 ;
        RECT 235.170 189.600 235.430 189.920 ;
        RECT 226.430 188.580 226.690 188.900 ;
        RECT 225.570 188.020 226.170 188.160 ;
        RECT 225.050 187.220 225.310 187.540 ;
        RECT 219.990 186.540 220.250 186.860 ;
        RECT 221.830 186.540 222.090 186.860 ;
        RECT 222.290 186.540 222.550 186.860 ;
        RECT 219.530 185.520 219.790 185.840 ;
        RECT 219.060 180.565 219.340 180.935 ;
        RECT 218.610 178.720 218.870 179.040 ;
        RECT 219.590 178.360 219.730 185.520 ;
        RECT 220.050 183.120 220.190 186.540 ;
        RECT 222.350 184.480 222.490 186.540 ;
        RECT 222.750 186.200 223.010 186.520 ;
        RECT 223.210 186.200 223.470 186.520 ;
        RECT 222.810 184.820 222.950 186.200 ;
        RECT 222.750 184.500 223.010 184.820 ;
        RECT 222.290 184.160 222.550 184.480 ;
        RECT 221.370 184.050 221.630 184.140 ;
        RECT 221.370 183.910 222.030 184.050 ;
        RECT 221.370 183.820 221.630 183.910 ;
        RECT 219.990 182.800 220.250 183.120 ;
        RECT 219.910 182.265 221.450 182.635 ;
        RECT 221.370 181.615 221.630 181.760 ;
        RECT 221.360 181.245 221.640 181.615 ;
        RECT 219.070 178.215 219.330 178.360 ;
        RECT 219.060 177.845 219.340 178.215 ;
        RECT 219.530 178.040 219.790 178.360 ;
        RECT 220.900 177.845 221.180 178.215 ;
        RECT 220.970 177.590 221.110 177.845 ;
        RECT 221.890 177.680 222.030 183.910 ;
        RECT 223.270 183.370 223.410 186.200 ;
        RECT 225.110 186.090 225.250 187.220 ;
        RECT 224.650 185.950 225.250 186.090 ;
        RECT 223.670 185.520 223.930 185.840 ;
        RECT 223.730 185.015 223.870 185.520 ;
        RECT 223.660 184.645 223.940 185.015 ;
        RECT 223.730 184.140 223.870 184.645 ;
        RECT 224.650 184.140 224.790 185.950 ;
        RECT 225.040 185.325 225.320 185.695 ;
        RECT 223.670 183.820 223.930 184.140 ;
        RECT 224.590 183.820 224.850 184.140 ;
        RECT 222.350 183.230 223.410 183.370 ;
        RECT 222.350 178.895 222.490 183.230 ;
        RECT 223.200 182.860 223.480 182.975 ;
        RECT 222.810 182.720 223.480 182.860 ;
        RECT 222.280 178.525 222.560 178.895 ;
        RECT 215.910 177.280 216.970 177.420 ;
        RECT 215.910 176.740 216.050 177.280 ;
        RECT 217.220 177.165 217.500 177.535 ;
        RECT 217.750 177.450 218.350 177.590 ;
        RECT 219.130 177.450 221.110 177.590 ;
        RECT 217.750 176.740 217.890 177.450 ;
        RECT 214.930 176.340 215.190 176.660 ;
        RECT 215.450 176.600 216.050 176.740 ;
        RECT 216.370 176.600 216.970 176.740 ;
        RECT 215.450 176.290 215.590 176.600 ;
        RECT 216.370 176.290 216.510 176.600 ;
        RECT 216.830 176.320 216.970 176.600 ;
        RECT 217.290 176.600 217.890 176.740 ;
        RECT 218.210 176.600 218.810 176.740 ;
        RECT 212.160 175.805 212.440 176.175 ;
        RECT 212.620 132.685 212.900 176.290 ;
        RECT 213.540 133.265 213.820 176.290 ;
        RECT 214.460 133.845 214.740 176.290 ;
        RECT 215.380 134.425 215.660 176.290 ;
        RECT 216.300 135.005 216.580 176.290 ;
        RECT 216.770 176.000 217.030 176.320 ;
        RECT 217.290 176.290 217.430 176.600 ;
        RECT 218.210 176.290 218.350 176.600 ;
        RECT 217.220 135.585 217.500 176.290 ;
        RECT 218.140 136.165 218.420 176.290 ;
        RECT 218.670 176.175 218.810 176.600 ;
        RECT 219.130 176.290 219.270 177.450 ;
        RECT 221.830 177.360 222.090 177.680 ;
        RECT 219.910 176.825 221.450 177.195 ;
        RECT 221.370 176.570 221.630 176.660 ;
        RECT 220.050 176.430 220.650 176.570 ;
        RECT 220.050 176.290 220.190 176.430 ;
        RECT 218.600 175.805 218.880 176.175 ;
        RECT 219.060 136.745 219.340 176.290 ;
        RECT 219.980 137.325 220.260 176.290 ;
        RECT 220.510 174.960 220.650 176.430 ;
        RECT 220.970 176.430 221.630 176.570 ;
        RECT 220.970 176.290 221.110 176.430 ;
        RECT 221.370 176.340 221.630 176.430 ;
        RECT 221.890 176.600 222.490 176.740 ;
        RECT 221.890 176.290 222.030 176.600 ;
        RECT 220.450 174.640 220.710 174.960 ;
        RECT 220.900 137.905 221.180 176.290 ;
        RECT 221.820 138.485 222.100 176.290 ;
        RECT 222.350 175.640 222.490 176.600 ;
        RECT 222.810 176.290 222.950 182.720 ;
        RECT 223.200 182.605 223.480 182.720 ;
        RECT 223.730 180.310 223.870 183.820 ;
        RECT 225.110 183.655 225.250 185.325 ;
        RECT 225.040 183.285 225.320 183.655 ;
        RECT 224.590 182.800 224.850 183.120 ;
        RECT 224.130 181.615 224.390 181.760 ;
        RECT 224.120 181.245 224.400 181.615 ;
        RECT 224.130 180.310 224.390 180.400 ;
        RECT 223.730 180.170 224.390 180.310 ;
        RECT 223.200 179.205 223.480 179.575 ;
        RECT 223.270 176.660 223.410 179.205 ;
        RECT 223.730 179.040 223.870 180.170 ;
        RECT 224.130 180.080 224.390 180.170 ;
        RECT 224.650 179.575 224.790 182.800 ;
        RECT 225.050 180.080 225.310 180.400 ;
        RECT 224.580 179.205 224.860 179.575 ;
        RECT 223.670 178.720 223.930 179.040 ;
        RECT 225.110 178.780 225.250 180.080 ;
        RECT 224.190 178.640 225.250 178.780 ;
        RECT 224.190 177.590 224.330 178.640 ;
        RECT 224.590 178.100 224.850 178.360 ;
        RECT 224.590 178.040 225.250 178.100 ;
        RECT 224.650 177.960 225.250 178.040 ;
        RECT 224.190 177.450 224.790 177.590 ;
        RECT 224.120 176.740 224.400 176.855 ;
        RECT 223.210 176.340 223.470 176.660 ;
        RECT 223.730 176.600 224.400 176.740 ;
        RECT 223.730 176.290 223.870 176.600 ;
        RECT 224.120 176.485 224.400 176.600 ;
        RECT 224.650 176.290 224.790 177.450 ;
        RECT 225.110 176.660 225.250 177.960 ;
        RECT 225.050 176.340 225.310 176.660 ;
        RECT 225.570 176.290 225.710 188.020 ;
        RECT 226.490 187.450 226.630 188.580 ;
        RECT 226.030 187.310 226.630 187.450 ;
        RECT 226.030 183.800 226.170 187.310 ;
        RECT 226.950 186.770 227.090 189.260 ;
        RECT 227.410 189.240 227.550 189.405 ;
        RECT 230.630 189.240 230.770 189.520 ;
        RECT 227.350 188.920 227.610 189.240 ;
        RECT 228.730 188.920 228.990 189.240 ;
        RECT 227.810 188.580 228.070 188.900 ;
        RECT 227.340 187.365 227.620 187.735 ;
        RECT 227.870 187.450 228.010 188.580 ;
        RECT 228.790 188.560 228.930 188.920 ;
        RECT 229.190 188.580 229.450 188.900 ;
        RECT 230.100 188.725 230.380 189.095 ;
        RECT 230.570 188.920 230.830 189.240 ;
        RECT 231.950 189.150 232.210 189.240 ;
        RECT 231.090 189.010 232.210 189.150 ;
        RECT 228.730 188.240 228.990 188.560 ;
        RECT 227.410 186.860 227.550 187.365 ;
        RECT 227.870 187.310 228.930 187.450 ;
        RECT 226.490 186.630 227.090 186.770 ;
        RECT 226.490 186.260 226.630 186.630 ;
        RECT 227.350 186.540 227.610 186.860 ;
        RECT 227.800 186.685 228.080 187.055 ;
        RECT 228.790 186.860 228.930 187.310 ;
        RECT 227.810 186.540 228.070 186.685 ;
        RECT 228.730 186.540 228.990 186.860 ;
        RECT 226.490 186.120 227.550 186.260 ;
        RECT 225.970 183.480 226.230 183.800 ;
        RECT 226.030 181.760 226.170 183.480 ;
        RECT 226.420 183.285 226.700 183.655 ;
        RECT 225.970 181.440 226.230 181.760 ;
        RECT 226.030 180.935 226.170 181.440 ;
        RECT 226.490 181.420 226.630 183.285 ;
        RECT 226.430 181.100 226.690 181.420 ;
        RECT 225.960 180.565 226.240 180.935 ;
        RECT 226.030 178.360 226.170 180.565 ;
        RECT 226.430 180.420 226.690 180.740 ;
        RECT 225.970 178.040 226.230 178.360 ;
        RECT 226.490 178.270 226.630 180.420 ;
        RECT 226.490 178.130 227.090 178.270 ;
        RECT 226.950 177.420 227.090 178.130 ;
        RECT 226.030 177.280 227.090 177.420 ;
        RECT 222.290 175.320 222.550 175.640 ;
        RECT 222.740 139.065 223.020 176.290 ;
        RECT 223.660 139.645 223.940 176.290 ;
        RECT 224.580 140.225 224.860 176.290 ;
        RECT 225.500 140.805 225.780 176.290 ;
        RECT 226.030 175.300 226.170 177.280 ;
        RECT 226.490 176.430 227.090 176.570 ;
        RECT 226.490 176.290 226.630 176.430 ;
        RECT 225.970 174.980 226.230 175.300 ;
        RECT 226.420 141.385 226.700 176.290 ;
        RECT 226.950 175.300 227.090 176.430 ;
        RECT 227.410 176.290 227.550 186.120 ;
        RECT 229.250 185.750 229.390 188.580 ;
        RECT 230.170 188.560 230.310 188.725 ;
        RECT 230.110 188.240 230.370 188.560 ;
        RECT 228.330 185.610 229.390 185.750 ;
        RECT 227.800 182.605 228.080 182.975 ;
        RECT 227.870 178.270 228.010 182.605 ;
        RECT 228.330 179.040 228.470 185.610 ;
        RECT 229.165 184.985 230.705 185.355 ;
        RECT 231.090 184.050 231.230 189.010 ;
        RECT 231.950 188.920 232.210 189.010 ;
        RECT 231.490 188.240 231.750 188.560 ;
        RECT 230.170 183.910 231.230 184.050 ;
        RECT 228.720 180.565 229.000 180.935 ;
        RECT 228.730 180.420 228.990 180.565 ;
        RECT 230.170 180.310 230.310 183.910 ;
        RECT 231.550 181.420 231.690 188.240 ;
        RECT 232.470 186.860 232.610 189.520 ;
        RECT 232.870 189.260 233.130 189.580 ;
        RECT 231.950 186.540 232.210 186.860 ;
        RECT 232.410 186.540 232.670 186.860 ;
        RECT 232.010 186.375 232.150 186.540 ;
        RECT 231.940 186.005 232.220 186.375 ;
        RECT 232.410 185.520 232.670 185.840 ;
        RECT 232.470 184.820 232.610 185.520 ;
        RECT 232.410 184.500 232.670 184.820 ;
        RECT 231.950 184.160 232.210 184.480 ;
        RECT 232.010 181.420 232.150 184.160 ;
        RECT 232.410 183.655 232.670 183.800 ;
        RECT 232.400 183.285 232.680 183.655 ;
        RECT 232.410 182.800 232.670 183.120 ;
        RECT 232.930 182.975 233.070 189.260 ;
        RECT 233.330 188.240 233.590 188.560 ;
        RECT 231.490 181.100 231.750 181.420 ;
        RECT 231.950 181.100 232.210 181.420 ;
        RECT 231.940 180.820 232.220 180.935 ;
        RECT 231.550 180.680 232.220 180.820 ;
        RECT 230.170 180.170 231.230 180.310 ;
        RECT 229.165 179.545 230.705 179.915 ;
        RECT 231.090 179.290 231.230 180.170 ;
        RECT 230.170 179.150 231.230 179.290 ;
        RECT 228.270 178.720 228.530 179.040 ;
        RECT 229.190 178.270 229.450 178.360 ;
        RECT 227.870 178.130 228.470 178.270 ;
        RECT 228.330 176.290 228.470 178.130 ;
        RECT 228.790 178.130 229.450 178.270 ;
        RECT 228.790 177.535 228.930 178.130 ;
        RECT 229.190 178.040 229.450 178.130 ;
        RECT 228.720 177.165 229.000 177.535 ;
        RECT 229.640 177.420 229.920 177.535 ;
        RECT 229.250 177.280 229.920 177.420 ;
        RECT 229.250 176.290 229.390 177.280 ;
        RECT 229.640 177.165 229.920 177.280 ;
        RECT 230.170 176.290 230.310 179.150 ;
        RECT 231.550 178.780 231.690 180.680 ;
        RECT 231.940 180.565 232.220 180.680 ;
        RECT 232.470 179.040 232.610 182.800 ;
        RECT 232.860 182.605 233.140 182.975 ;
        RECT 232.860 181.245 233.140 181.615 ;
        RECT 231.090 178.640 231.690 178.780 ;
        RECT 232.410 178.720 232.670 179.040 ;
        RECT 232.930 178.700 233.070 181.245 ;
        RECT 231.090 176.290 231.230 178.640 ;
        RECT 232.870 178.380 233.130 178.700 ;
        RECT 231.490 178.040 231.750 178.360 ;
        RECT 232.410 178.040 232.670 178.360 ;
        RECT 231.550 176.320 231.690 178.040 ;
        RECT 226.890 174.980 227.150 175.300 ;
        RECT 227.340 141.965 227.620 176.290 ;
        RECT 228.260 142.545 228.540 176.290 ;
        RECT 229.180 143.125 229.460 176.290 ;
        RECT 230.100 143.705 230.380 176.290 ;
        RECT 231.020 144.285 231.300 176.290 ;
        RECT 231.490 176.000 231.750 176.320 ;
        RECT 232.470 176.175 232.610 178.040 ;
        RECT 233.390 176.660 233.530 188.240 ;
        RECT 234.240 187.365 234.520 187.735 ;
        RECT 233.780 186.685 234.060 187.055 ;
        RECT 233.850 179.040 233.990 186.685 ;
        RECT 234.310 186.180 234.450 187.365 ;
        RECT 234.250 185.860 234.510 186.180 ;
        RECT 234.250 184.335 234.510 184.480 ;
        RECT 234.240 183.965 234.520 184.335 ;
        RECT 235.230 183.800 235.370 189.600 ;
        RECT 236.150 187.540 236.290 199.800 ;
        RECT 238.420 198.585 239.960 198.955 ;
        RECT 238.420 193.145 239.960 193.515 ;
        RECT 238.420 187.705 239.960 188.075 ;
        RECT 236.090 187.220 236.350 187.540 ;
        RECT 236.090 186.540 236.350 186.860 ;
        RECT 237.470 186.540 237.730 186.860 ;
        RECT 234.710 183.480 234.970 183.800 ;
        RECT 235.170 183.480 235.430 183.800 ;
        RECT 233.790 178.720 234.050 179.040 ;
        RECT 233.790 178.215 234.050 178.360 ;
        RECT 233.780 177.845 234.060 178.215 ;
        RECT 234.250 177.360 234.510 177.680 ;
        RECT 234.310 176.660 234.450 177.360 ;
        RECT 234.770 176.855 234.910 183.480 ;
        RECT 235.630 182.800 235.890 183.120 ;
        RECT 235.690 182.100 235.830 182.800 ;
        RECT 235.630 181.780 235.890 182.100 ;
        RECT 236.150 181.500 236.290 186.540 ;
        RECT 235.690 181.360 236.290 181.500 ;
        RECT 235.170 178.040 235.430 178.360 ;
        RECT 233.330 176.340 233.590 176.660 ;
        RECT 234.250 176.340 234.510 176.660 ;
        RECT 234.700 176.485 234.980 176.855 ;
        RECT 232.400 175.805 232.680 176.175 ;
        RECT 235.230 174.960 235.370 178.040 ;
        RECT 235.690 177.535 235.830 181.360 ;
        RECT 237.530 180.935 237.670 186.540 ;
        RECT 237.930 183.480 238.190 183.800 ;
        RECT 237.460 180.565 237.740 180.935 ;
        RECT 236.090 180.080 236.350 180.400 ;
        RECT 236.550 180.080 236.810 180.400 ;
        RECT 235.620 177.165 235.900 177.535 ;
        RECT 235.170 174.640 235.430 174.960 ;
        RECT 236.150 174.815 236.290 180.080 ;
        RECT 236.610 179.380 236.750 180.080 ;
        RECT 236.550 179.060 236.810 179.380 ;
        RECT 236.550 178.040 236.810 178.360 ;
        RECT 236.610 175.640 236.750 178.040 ;
        RECT 236.550 175.320 236.810 175.640 ;
        RECT 237.990 175.300 238.130 183.480 ;
        RECT 238.420 182.265 239.960 182.635 ;
        RECT 238.420 176.825 239.960 177.195 ;
        RECT 237.930 174.980 238.190 175.300 ;
        RECT 236.080 174.445 236.360 174.815 ;
        RECT 231.020 144.005 309.205 144.285 ;
        RECT 230.100 143.425 306.905 143.705 ;
        RECT 229.180 142.845 304.605 143.125 ;
        RECT 228.260 142.265 302.305 142.545 ;
        RECT 227.340 141.685 300.005 141.965 ;
        RECT 226.420 141.105 297.705 141.385 ;
        RECT 225.500 140.525 295.405 140.805 ;
        RECT 224.580 139.945 293.105 140.225 ;
        RECT 223.660 139.365 290.805 139.645 ;
        RECT 222.740 138.785 288.505 139.065 ;
        RECT 221.820 138.205 286.205 138.485 ;
        RECT 220.900 137.625 283.905 137.905 ;
        RECT 219.980 137.045 281.605 137.325 ;
        RECT 219.060 136.465 279.305 136.745 ;
        RECT 218.140 135.885 277.005 136.165 ;
        RECT 217.220 135.305 274.705 135.585 ;
        RECT 216.300 134.725 272.405 135.005 ;
        RECT 215.380 134.145 270.105 134.425 ;
        RECT 214.460 133.565 267.805 133.845 ;
        RECT 213.540 132.985 265.505 133.265 ;
        RECT 212.620 132.405 263.205 132.685 ;
        RECT 211.700 131.825 260.905 132.105 ;
        RECT 210.780 131.245 258.605 131.525 ;
        RECT 209.860 130.665 256.305 130.945 ;
        RECT 208.940 130.085 254.005 130.365 ;
        RECT 208.020 129.505 251.705 129.785 ;
        RECT 207.100 128.925 249.405 129.205 ;
        RECT 206.180 128.345 247.105 128.625 ;
        RECT 205.260 127.765 244.805 128.045 ;
        RECT 204.340 127.185 242.505 127.465 ;
        RECT 203.420 126.605 240.205 126.885 ;
        RECT 202.500 126.025 237.905 126.305 ;
        RECT 201.580 125.445 235.605 125.725 ;
        RECT 200.660 124.865 233.305 125.145 ;
        RECT 199.740 124.285 231.005 124.565 ;
        RECT 198.820 123.705 228.705 123.985 ;
        RECT 197.900 123.125 226.405 123.405 ;
        RECT 196.980 122.545 224.105 122.825 ;
        RECT 196.060 121.965 221.805 122.245 ;
        RECT 195.140 121.385 219.505 121.665 ;
        RECT 194.220 120.805 217.205 121.085 ;
        RECT 193.300 120.225 214.905 120.505 ;
        RECT 192.380 119.645 212.605 119.925 ;
        RECT 191.460 119.065 210.305 119.345 ;
        RECT 190.540 118.485 208.005 118.765 ;
        RECT 189.620 117.905 205.705 118.185 ;
        RECT 188.700 117.325 203.405 117.605 ;
        RECT 187.780 116.745 201.105 117.025 ;
        RECT 186.860 116.165 198.805 116.445 ;
        RECT 185.940 115.585 196.505 115.865 ;
        RECT 185.020 115.005 194.205 115.285 ;
        RECT 184.100 114.425 191.905 114.705 ;
        RECT 183.180 113.845 189.605 114.125 ;
        RECT 182.260 113.265 187.305 113.545 ;
        RECT 181.340 112.685 185.005 112.965 ;
        RECT 180.420 112.105 182.705 112.385 ;
        RECT 179.500 111.525 180.405 111.805 ;
        RECT 177.825 109.225 178.105 111.525 ;
        RECT 180.125 109.225 180.405 111.525 ;
        RECT 182.425 109.225 182.705 112.105 ;
        RECT 184.725 109.225 185.005 112.685 ;
        RECT 187.025 109.225 187.305 113.265 ;
        RECT 189.325 109.225 189.605 113.845 ;
        RECT 191.625 109.225 191.905 114.425 ;
        RECT 193.925 109.225 194.205 115.005 ;
        RECT 196.225 109.225 196.505 115.585 ;
        RECT 198.525 109.225 198.805 116.165 ;
        RECT 200.825 109.225 201.105 116.745 ;
        RECT 203.125 109.225 203.405 117.325 ;
        RECT 205.425 109.225 205.705 117.905 ;
        RECT 207.725 109.225 208.005 118.485 ;
        RECT 210.025 109.225 210.305 119.065 ;
        RECT 212.325 109.225 212.605 119.645 ;
        RECT 214.625 109.225 214.905 120.225 ;
        RECT 216.925 109.225 217.205 120.805 ;
        RECT 219.225 109.225 219.505 121.385 ;
        RECT 221.525 109.225 221.805 121.965 ;
        RECT 223.825 109.225 224.105 122.545 ;
        RECT 226.125 109.225 226.405 123.125 ;
        RECT 228.425 109.225 228.705 123.705 ;
        RECT 230.725 109.225 231.005 124.285 ;
        RECT 233.025 109.225 233.305 124.865 ;
        RECT 235.325 109.225 235.605 125.445 ;
        RECT 237.625 109.225 237.905 126.025 ;
        RECT 239.925 109.225 240.205 126.605 ;
        RECT 242.225 109.225 242.505 127.185 ;
        RECT 244.525 109.225 244.805 127.765 ;
        RECT 246.825 109.225 247.105 128.345 ;
        RECT 249.125 109.225 249.405 128.925 ;
        RECT 251.425 109.225 251.705 129.505 ;
        RECT 253.725 109.225 254.005 130.085 ;
        RECT 256.025 109.225 256.305 130.665 ;
        RECT 258.325 109.225 258.605 131.245 ;
        RECT 260.625 109.225 260.905 131.825 ;
        RECT 262.925 109.225 263.205 132.405 ;
        RECT 265.225 109.225 265.505 132.985 ;
        RECT 267.525 109.225 267.805 133.565 ;
        RECT 269.825 109.225 270.105 134.145 ;
        RECT 272.125 109.225 272.405 134.725 ;
        RECT 274.425 109.225 274.705 135.305 ;
        RECT 276.725 109.225 277.005 135.885 ;
        RECT 279.025 109.225 279.305 136.465 ;
        RECT 281.325 109.225 281.605 137.045 ;
        RECT 283.625 109.225 283.905 137.625 ;
        RECT 285.925 109.225 286.205 138.205 ;
        RECT 288.225 109.225 288.505 138.785 ;
        RECT 290.525 109.225 290.805 139.365 ;
        RECT 292.825 109.225 293.105 139.945 ;
        RECT 295.125 109.225 295.405 140.525 ;
        RECT 297.425 109.225 297.705 141.105 ;
        RECT 299.725 109.225 300.005 141.685 ;
        RECT 302.025 109.225 302.305 142.265 ;
        RECT 304.325 109.225 304.605 142.845 ;
        RECT 306.625 109.225 306.905 143.425 ;
        RECT 308.925 109.225 309.205 144.005 ;
        RECT 164.095 106.075 164.235 109.225 ;
        RECT 166.395 106.075 166.535 109.225 ;
        RECT 164.035 105.755 164.295 106.075 ;
        RECT 166.335 105.755 166.595 106.075 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 165.875 103.035 166.135 103.355 ;
        RECT 165.415 102.015 165.675 102.335 ;
        RECT 163.575 94.195 163.835 94.515 ;
        RECT 163.635 93.350 163.775 94.195 ;
        RECT 165.475 93.835 165.615 102.015 ;
        RECT 165.935 99.955 166.075 103.035 ;
        RECT 166.795 101.675 167.055 101.995 ;
        RECT 166.855 100.635 166.995 101.675 ;
        RECT 168.695 100.715 168.835 109.225 ;
        RECT 170.995 106.075 171.135 109.225 ;
        RECT 173.295 106.075 173.435 109.225 ;
        RECT 170.935 105.755 171.195 106.075 ;
        RECT 173.235 105.755 173.495 106.075 ;
        RECT 174.155 105.075 174.415 105.395 ;
        RECT 174.615 105.075 174.875 105.395 ;
        RECT 173.695 104.055 173.955 104.375 ;
        RECT 172.775 102.355 173.035 102.675 ;
        RECT 168.235 100.635 168.835 100.715 ;
        RECT 166.795 100.315 167.055 100.635 ;
        RECT 168.175 100.575 168.835 100.635 ;
        RECT 168.175 100.315 168.435 100.575 ;
        RECT 172.835 100.295 172.975 102.355 ;
        RECT 172.775 99.975 173.035 100.295 ;
        RECT 165.875 99.635 166.135 99.955 ;
        RECT 168.175 99.635 168.435 99.955 ;
        RECT 165.875 94.195 166.135 94.515 ;
        RECT 165.415 93.515 165.675 93.835 ;
        RECT 163.565 92.980 163.845 93.350 ;
        RECT 146.290 88.455 148.395 92.555 ;
        RECT 165.475 91.795 165.615 93.515 ;
        RECT 165.935 92.475 166.075 94.195 ;
        RECT 165.875 92.155 166.135 92.475 ;
        RECT 165.415 91.475 165.675 91.795 ;
        RECT 165.475 89.075 165.615 91.475 ;
        RECT 164.955 88.755 165.215 89.075 ;
        RECT 165.415 88.755 165.675 89.075 ;
        RECT 146.290 83.775 148.395 87.875 ;
        RECT 165.015 87.035 165.155 88.755 ;
        RECT 168.235 88.735 168.375 99.635 ;
        RECT 170.015 99.295 170.275 99.615 ;
        RECT 170.075 97.915 170.215 99.295 ;
        RECT 170.015 97.595 170.275 97.915 ;
        RECT 172.835 97.315 172.975 99.975 ;
        RECT 172.835 97.175 173.435 97.315 ;
        RECT 170.015 95.895 170.275 96.215 ;
        RECT 171.395 95.895 171.655 96.215 ;
        RECT 170.075 91.795 170.215 95.895 ;
        RECT 171.455 94.855 171.595 95.895 ;
        RECT 173.295 94.855 173.435 97.175 ;
        RECT 171.395 94.535 171.655 94.855 ;
        RECT 173.235 94.535 173.495 94.855 ;
        RECT 170.015 91.475 170.275 91.795 ;
        RECT 173.295 91.455 173.435 94.535 ;
        RECT 173.235 91.135 173.495 91.455 ;
        RECT 173.295 89.075 173.435 91.135 ;
        RECT 173.755 90.775 173.895 104.055 ;
        RECT 174.215 101.510 174.355 105.075 ;
        RECT 174.145 101.140 174.425 101.510 ;
        RECT 174.155 96.235 174.415 96.555 ;
        RECT 174.215 92.475 174.355 96.235 ;
        RECT 174.155 92.155 174.415 92.475 ;
        RECT 173.695 90.455 173.955 90.775 ;
        RECT 173.235 88.755 173.495 89.075 ;
        RECT 168.175 88.415 168.435 88.735 ;
        RECT 172.775 88.415 173.035 88.735 ;
        RECT 164.955 86.715 165.215 87.035 ;
        RECT 172.835 86.015 172.975 88.415 ;
        RECT 172.775 85.695 173.035 86.015 ;
        RECT 146.290 77.925 148.395 83.195 ;
        RECT 174.155 80.935 174.415 81.255 ;
        RECT 173.235 80.255 173.495 80.575 ;
        RECT 169.555 79.575 169.815 79.895 ;
        RECT 170.935 79.575 171.195 79.895 ;
        RECT 146.290 73.245 148.395 77.345 ;
        RECT 169.615 75.475 169.755 79.575 ;
        RECT 170.995 78.535 171.135 79.575 ;
        RECT 170.935 78.215 171.195 78.535 ;
        RECT 172.775 78.215 173.035 78.535 ;
        RECT 172.835 76.155 172.975 78.215 ;
        RECT 173.295 76.155 173.435 80.255 ;
        RECT 172.775 75.835 173.035 76.155 ;
        RECT 173.235 75.835 173.495 76.155 ;
        RECT 169.555 75.155 169.815 75.475 ;
        RECT 165.415 74.815 165.675 75.135 ;
        RECT 146.290 68.565 148.395 72.665 ;
        RECT 165.475 69.695 165.615 74.815 ;
        RECT 172.835 73.395 172.975 75.835 ;
        RECT 174.215 73.435 174.355 80.935 ;
        RECT 172.375 73.255 172.975 73.395 ;
        RECT 170.015 71.415 170.275 71.735 ;
        RECT 170.075 70.035 170.215 71.415 ;
        RECT 170.015 69.715 170.275 70.035 ;
        RECT 172.375 69.695 172.515 73.255 ;
        RECT 174.155 73.115 174.415 73.435 ;
        RECT 165.415 69.375 165.675 69.695 ;
        RECT 172.315 69.375 172.575 69.695 ;
        RECT 146.290 63.885 148.395 67.985 ;
        RECT 165.475 66.635 165.615 69.375 ;
        RECT 171.395 68.695 171.655 69.015 ;
        RECT 171.455 67.315 171.595 68.695 ;
        RECT 172.375 67.995 172.515 69.375 ;
        RECT 172.315 67.675 172.575 67.995 ;
        RECT 170.015 66.995 170.275 67.315 ;
        RECT 171.395 66.995 171.655 67.315 ;
        RECT 165.415 66.315 165.675 66.635 ;
        RECT 165.475 64.255 165.615 66.315 ;
        RECT 169.095 65.975 169.355 66.295 ;
        RECT 169.155 64.595 169.295 65.975 ;
        RECT 170.075 65.275 170.215 66.995 ;
        RECT 170.015 64.955 170.275 65.275 ;
        RECT 169.095 64.275 169.355 64.595 ;
        RECT 172.375 64.255 172.515 67.675 ;
        RECT 165.415 63.935 165.675 64.255 ;
        RECT 172.315 63.935 172.575 64.255 ;
        RECT 146.290 58.035 148.395 63.305 ;
        RECT 174.145 62.380 174.425 62.750 ;
        RECT 174.215 61.535 174.355 62.380 ;
        RECT 174.155 61.215 174.415 61.535 ;
        RECT 164.035 60.710 164.295 60.855 ;
        RECT 164.025 60.340 164.305 60.710 ;
        RECT 168.635 60.535 168.895 60.855 ;
        RECT 168.695 59.155 168.835 60.535 ;
        RECT 168.635 58.835 168.895 59.155 ;
        RECT 165.415 58.495 165.675 58.815 ;
        RECT 174.215 58.670 174.355 61.215 ;
        RECT 174.675 59.155 174.815 105.075 ;
        RECT 175.595 103.435 175.735 109.225 ;
        RECT 177.895 106.075 178.035 109.225 ;
        RECT 180.195 106.075 180.335 109.225 ;
        RECT 177.835 105.755 178.095 106.075 ;
        RECT 180.135 105.755 180.395 106.075 ;
        RECT 181.975 105.415 182.235 105.735 ;
        RECT 177.375 105.075 177.635 105.395 ;
        RECT 181.515 105.075 181.775 105.395 ;
        RECT 175.595 103.355 176.195 103.435 ;
        RECT 175.595 103.295 176.255 103.355 ;
        RECT 175.995 103.035 176.255 103.295 ;
        RECT 177.435 96.895 177.575 105.075 ;
        RECT 181.575 104.910 181.715 105.075 ;
        RECT 181.505 104.540 181.785 104.910 ;
        RECT 178.295 104.055 178.555 104.375 ;
        RECT 177.835 98.615 178.095 98.935 ;
        RECT 177.895 97.915 178.035 98.615 ;
        RECT 177.835 97.595 178.095 97.915 ;
        RECT 177.375 96.750 177.635 96.895 ;
        RECT 177.365 96.380 177.645 96.750 ;
        RECT 177.435 95.195 177.575 96.380 ;
        RECT 177.835 95.895 178.095 96.215 ;
        RECT 177.375 94.875 177.635 95.195 ;
        RECT 177.895 94.515 178.035 95.895 ;
        RECT 177.835 94.195 178.095 94.515 ;
        RECT 177.365 91.620 177.645 91.990 ;
        RECT 177.895 91.795 178.035 94.195 ;
        RECT 177.435 91.115 177.575 91.620 ;
        RECT 177.835 91.475 178.095 91.795 ;
        RECT 177.375 90.795 177.635 91.115 ;
        RECT 175.065 88.220 175.345 88.590 ;
        RECT 177.375 88.415 177.635 88.735 ;
        RECT 175.075 88.075 175.335 88.220 ;
        RECT 175.995 86.715 176.255 87.035 ;
        RECT 175.075 72.435 175.335 72.755 ;
        RECT 175.525 72.580 175.805 72.950 ;
        RECT 175.535 72.435 175.795 72.580 ;
        RECT 175.135 62.555 175.275 72.435 ;
        RECT 175.595 70.715 175.735 72.435 ;
        RECT 175.535 70.395 175.795 70.715 ;
        RECT 175.075 62.235 175.335 62.555 ;
        RECT 176.055 61.535 176.195 86.715 ;
        RECT 177.435 86.695 177.575 88.415 ;
        RECT 177.375 86.375 177.635 86.695 ;
        RECT 178.355 84.315 178.495 104.055 ;
        RECT 179.955 103.520 181.495 103.890 ;
        RECT 178.755 102.355 179.015 102.675 ;
        RECT 178.815 98.935 178.955 102.355 ;
        RECT 179.215 98.955 179.475 99.275 ;
        RECT 178.755 98.615 179.015 98.935 ;
        RECT 178.815 97.235 178.955 98.615 ;
        RECT 178.755 96.915 179.015 97.235 ;
        RECT 178.755 91.475 179.015 91.795 ;
        RECT 178.815 86.355 178.955 91.475 ;
        RECT 179.275 91.115 179.415 98.955 ;
        RECT 179.955 98.080 181.495 98.450 ;
        RECT 179.955 92.640 181.495 93.010 ;
        RECT 179.215 90.795 179.475 91.115 ;
        RECT 178.755 86.035 179.015 86.355 ;
        RECT 179.275 85.335 179.415 90.795 ;
        RECT 182.035 89.755 182.175 105.415 ;
        RECT 182.495 104.715 182.635 109.225 ;
        RECT 184.795 106.075 184.935 109.225 ;
        RECT 187.095 106.075 187.235 109.225 ;
        RECT 184.735 105.755 184.995 106.075 ;
        RECT 187.035 105.755 187.295 106.075 ;
        RECT 185.195 105.075 185.455 105.395 ;
        RECT 185.655 105.075 185.915 105.395 ;
        RECT 186.115 105.305 186.375 105.395 ;
        RECT 186.115 105.165 186.775 105.305 ;
        RECT 186.115 105.075 186.375 105.165 ;
        RECT 182.435 104.395 182.695 104.715 ;
        RECT 183.355 102.355 183.615 102.675 ;
        RECT 182.435 101.675 182.695 101.995 ;
        RECT 182.895 101.675 183.155 101.995 ;
        RECT 181.975 89.435 182.235 89.755 ;
        RECT 179.955 87.200 181.495 87.570 ;
        RECT 182.035 86.015 182.175 89.435 ;
        RECT 182.495 87.035 182.635 101.675 ;
        RECT 182.955 99.275 183.095 101.675 ;
        RECT 182.895 98.955 183.155 99.275 ;
        RECT 183.415 96.895 183.555 102.355 ;
        RECT 185.255 99.955 185.395 105.075 ;
        RECT 185.715 102.675 185.855 105.075 ;
        RECT 185.655 102.355 185.915 102.675 ;
        RECT 185.715 100.295 185.855 102.355 ;
        RECT 185.655 99.975 185.915 100.295 ;
        RECT 185.195 99.635 185.455 99.955 ;
        RECT 185.255 97.235 185.395 99.635 ;
        RECT 186.115 99.295 186.375 99.615 ;
        RECT 186.175 97.430 186.315 99.295 ;
        RECT 185.195 96.915 185.455 97.235 ;
        RECT 186.105 97.060 186.385 97.430 ;
        RECT 183.355 96.575 183.615 96.895 ;
        RECT 184.735 96.235 184.995 96.555 ;
        RECT 184.275 95.895 184.535 96.215 ;
        RECT 184.335 94.175 184.475 95.895 ;
        RECT 184.795 95.195 184.935 96.235 ;
        RECT 184.735 94.875 184.995 95.195 ;
        RECT 184.275 93.855 184.535 94.175 ;
        RECT 182.895 91.135 183.155 91.455 ;
        RECT 182.955 88.395 183.095 91.135 ;
        RECT 182.895 88.075 183.155 88.395 ;
        RECT 182.435 86.715 182.695 87.035 ;
        RECT 181.975 85.695 182.235 86.015 ;
        RECT 179.215 85.015 179.475 85.335 ;
        RECT 178.295 83.995 178.555 84.315 ;
        RECT 182.955 83.975 183.095 88.075 ;
        RECT 184.335 88.055 184.475 93.855 ;
        RECT 186.175 91.795 186.315 97.060 ;
        RECT 186.115 91.475 186.375 91.795 ;
        RECT 186.635 91.195 186.775 105.165 ;
        RECT 189.395 105.055 189.535 109.225 ;
        RECT 190.255 105.075 190.515 105.395 ;
        RECT 189.335 104.735 189.595 105.055 ;
        RECT 190.315 103.355 190.455 105.075 ;
        RECT 191.695 105.055 191.835 109.225 ;
        RECT 193.995 106.075 194.135 109.225 ;
        RECT 196.295 106.075 196.435 109.225 ;
        RECT 198.595 107.515 198.735 109.225 ;
        RECT 198.135 107.375 198.735 107.515 ;
        RECT 198.135 106.075 198.275 107.375 ;
        RECT 198.585 106.240 200.125 106.610 ;
        RECT 200.895 106.075 201.035 109.225 ;
        RECT 193.935 105.755 194.195 106.075 ;
        RECT 196.235 105.755 196.495 106.075 ;
        RECT 198.075 105.755 198.335 106.075 ;
        RECT 200.835 105.755 201.095 106.075 ;
        RECT 196.695 105.415 196.955 105.735 ;
        RECT 197.155 105.415 197.415 105.735 ;
        RECT 199.915 105.415 200.175 105.735 ;
        RECT 195.315 105.075 195.575 105.395 ;
        RECT 195.775 105.075 196.035 105.395 ;
        RECT 191.635 104.735 191.895 105.055 ;
        RECT 190.255 103.035 190.515 103.355 ;
        RECT 190.245 102.500 190.525 102.870 ;
        RECT 190.255 102.355 190.515 102.500 ;
        RECT 192.555 101.675 192.815 101.995 ;
        RECT 194.855 101.675 195.115 101.995 ;
        RECT 190.255 101.335 190.515 101.655 ;
        RECT 191.635 101.335 191.895 101.655 ;
        RECT 187.035 100.315 187.295 100.635 ;
        RECT 184.795 91.055 186.775 91.195 ;
        RECT 184.275 87.735 184.535 88.055 ;
        RECT 184.335 86.355 184.475 87.735 ;
        RECT 184.275 86.035 184.535 86.355 ;
        RECT 184.275 85.355 184.535 85.675 ;
        RECT 182.895 83.655 183.155 83.975 ;
        RECT 179.955 81.760 181.495 82.130 ;
        RECT 178.755 80.595 179.015 80.915 ;
        RECT 177.375 80.430 177.635 80.575 ;
        RECT 176.455 79.915 176.715 80.235 ;
        RECT 177.365 80.060 177.645 80.430 ;
        RECT 176.515 77.515 176.655 79.915 ;
        RECT 176.915 79.575 177.175 79.895 ;
        RECT 176.975 78.535 177.115 79.575 ;
        RECT 176.915 78.215 177.175 78.535 ;
        RECT 176.455 77.195 176.715 77.515 ;
        RECT 177.435 72.415 177.575 80.060 ;
        RECT 177.835 79.575 178.095 79.895 ;
        RECT 177.895 78.390 178.035 79.575 ;
        RECT 177.825 78.020 178.105 78.390 ;
        RECT 177.835 77.535 178.095 77.855 ;
        RECT 177.895 75.475 178.035 77.535 ;
        RECT 178.295 76.855 178.555 77.175 ;
        RECT 178.355 75.475 178.495 76.855 ;
        RECT 178.815 75.475 178.955 80.595 ;
        RECT 179.675 78.445 179.935 78.535 ;
        RECT 179.275 78.305 179.935 78.445 ;
        RECT 179.275 75.815 179.415 78.305 ;
        RECT 179.675 78.215 179.935 78.305 ;
        RECT 179.955 76.320 181.495 76.690 ;
        RECT 179.215 75.495 179.475 75.815 ;
        RECT 177.835 75.155 178.095 75.475 ;
        RECT 178.295 75.155 178.555 75.475 ;
        RECT 178.755 75.155 179.015 75.475 ;
        RECT 177.835 74.135 178.095 74.455 ;
        RECT 177.895 73.095 178.035 74.135 ;
        RECT 177.835 72.775 178.095 73.095 ;
        RECT 178.815 72.835 178.955 75.155 ;
        RECT 179.205 74.620 179.485 74.990 ;
        RECT 181.975 74.815 182.235 75.135 ;
        RECT 179.215 74.475 179.475 74.620 ;
        RECT 179.275 73.435 179.415 74.475 ;
        RECT 179.215 73.115 179.475 73.435 ;
        RECT 176.455 72.095 176.715 72.415 ;
        RECT 177.375 72.095 177.635 72.415 ;
        RECT 176.515 70.035 176.655 72.095 ;
        RECT 176.455 69.715 176.715 70.035 ;
        RECT 177.375 69.035 177.635 69.355 ;
        RECT 177.435 65.275 177.575 69.035 ;
        RECT 177.375 64.955 177.635 65.275 ;
        RECT 175.995 61.215 176.255 61.535 ;
        RECT 175.075 60.535 175.335 60.855 ;
        RECT 174.615 58.835 174.875 59.155 ;
        RECT 146.290 53.355 148.395 57.455 ;
        RECT 165.475 57.115 165.615 58.495 ;
        RECT 174.145 58.300 174.425 58.670 ;
        RECT 174.215 58.135 174.355 58.300 ;
        RECT 174.155 57.815 174.415 58.135 ;
        RECT 174.615 57.815 174.875 58.135 ;
        RECT 165.415 56.795 165.675 57.115 ;
        RECT 165.475 54.395 165.615 56.795 ;
        RECT 174.675 56.435 174.815 57.815 ;
        RECT 174.615 56.115 174.875 56.435 ;
        RECT 169.095 55.775 169.355 56.095 ;
        RECT 166.795 55.095 167.055 55.415 ;
        RECT 165.415 54.075 165.675 54.395 ;
        RECT 166.855 53.715 166.995 55.095 ;
        RECT 169.155 54.395 169.295 55.775 ;
        RECT 169.095 54.075 169.355 54.395 ;
        RECT 174.675 54.055 174.815 56.115 ;
        RECT 175.135 55.415 175.275 60.535 ;
        RECT 176.455 58.835 176.715 59.155 ;
        RECT 175.995 57.815 176.255 58.135 ;
        RECT 175.075 55.095 175.335 55.415 ;
        RECT 176.055 54.395 176.195 57.815 ;
        RECT 176.515 56.095 176.655 58.835 ;
        RECT 177.375 58.495 177.635 58.815 ;
        RECT 177.435 56.435 177.575 58.495 ;
        RECT 177.895 58.475 178.035 72.775 ;
        RECT 178.815 72.695 179.415 72.835 ;
        RECT 178.295 72.095 178.555 72.415 ;
        RECT 178.355 62.555 178.495 72.095 ;
        RECT 178.755 71.415 179.015 71.735 ;
        RECT 178.815 69.265 178.955 71.415 ;
        RECT 179.275 70.035 179.415 72.695 ;
        RECT 179.955 70.880 181.495 71.250 ;
        RECT 179.215 69.715 179.475 70.035 ;
        RECT 179.215 69.265 179.475 69.355 ;
        RECT 178.815 69.125 179.475 69.265 ;
        RECT 178.815 64.595 178.955 69.125 ;
        RECT 179.215 69.035 179.475 69.125 ;
        RECT 180.595 68.695 180.855 69.015 ;
        RECT 180.655 66.830 180.795 68.695 ;
        RECT 182.035 66.975 182.175 74.815 ;
        RECT 183.345 70.540 183.625 70.910 ;
        RECT 183.415 70.035 183.555 70.540 ;
        RECT 183.355 69.715 183.615 70.035 ;
        RECT 180.585 66.460 180.865 66.830 ;
        RECT 181.975 66.655 182.235 66.975 ;
        RECT 180.595 66.315 180.855 66.460 ;
        RECT 179.955 65.440 181.495 65.810 ;
        RECT 181.975 64.615 182.235 64.935 ;
        RECT 178.755 64.275 179.015 64.595 ;
        RECT 178.295 62.235 178.555 62.555 ;
        RECT 178.755 61.215 179.015 61.535 ;
        RECT 179.215 61.215 179.475 61.535 ;
        RECT 178.815 58.555 178.955 61.215 ;
        RECT 179.275 59.155 179.415 61.215 ;
        RECT 179.955 60.000 181.495 60.370 ;
        RECT 179.215 58.835 179.475 59.155 ;
        RECT 177.835 58.155 178.095 58.475 ;
        RECT 178.815 58.415 179.415 58.555 ;
        RECT 177.375 56.115 177.635 56.435 ;
        RECT 176.455 55.775 176.715 56.095 ;
        RECT 175.995 54.075 176.255 54.395 ;
        RECT 174.615 53.735 174.875 54.055 ;
        RECT 166.795 53.395 167.055 53.715 ;
        RECT 174.155 53.230 174.415 53.375 ;
        RECT 174.145 52.860 174.425 53.230 ;
        RECT 146.290 48.675 148.395 52.775 ;
        RECT 177.435 48.275 177.575 56.115 ;
        RECT 178.755 55.775 179.015 56.095 ;
        RECT 178.815 54.395 178.955 55.775 ;
        RECT 178.755 54.075 179.015 54.395 ;
        RECT 178.745 53.115 179.025 53.230 ;
        RECT 179.275 53.115 179.415 58.415 ;
        RECT 182.035 58.135 182.175 64.615 ;
        RECT 184.335 62.555 184.475 85.355 ;
        RECT 184.795 74.990 184.935 91.055 ;
        RECT 186.575 90.455 186.835 90.775 ;
        RECT 185.655 87.735 185.915 88.055 ;
        RECT 185.715 85.675 185.855 87.735 ;
        RECT 186.635 86.550 186.775 90.455 ;
        RECT 186.115 86.035 186.375 86.355 ;
        RECT 186.565 86.180 186.845 86.550 ;
        RECT 185.655 85.355 185.915 85.675 ;
        RECT 186.175 80.915 186.315 86.035 ;
        RECT 186.635 84.315 186.775 86.180 ;
        RECT 186.575 83.995 186.835 84.315 ;
        RECT 186.115 80.595 186.375 80.915 ;
        RECT 187.095 78.875 187.235 100.315 ;
        RECT 190.315 99.615 190.455 101.335 ;
        RECT 189.795 99.295 190.055 99.615 ;
        RECT 190.255 99.295 190.515 99.615 ;
        RECT 189.855 97.915 189.995 99.295 ;
        RECT 189.795 97.595 190.055 97.915 ;
        RECT 190.315 91.795 190.455 99.295 ;
        RECT 191.695 96.555 191.835 101.335 ;
        RECT 192.095 97.255 192.355 97.575 ;
        RECT 191.635 96.235 191.895 96.555 ;
        RECT 190.255 91.475 190.515 91.795 ;
        RECT 189.335 90.795 189.595 91.115 ;
        RECT 188.875 90.455 189.135 90.775 ;
        RECT 188.935 89.755 189.075 90.455 ;
        RECT 189.395 89.755 189.535 90.795 ;
        RECT 188.875 89.435 189.135 89.755 ;
        RECT 189.335 89.435 189.595 89.755 ;
        RECT 188.875 88.415 189.135 88.735 ;
        RECT 188.415 87.735 188.675 88.055 ;
        RECT 188.475 83.975 188.615 87.735 ;
        RECT 188.935 87.035 189.075 88.415 ;
        RECT 188.875 86.715 189.135 87.035 ;
        RECT 188.415 83.655 188.675 83.975 ;
        RECT 188.935 83.635 189.075 86.715 ;
        RECT 190.315 85.335 190.455 91.475 ;
        RECT 191.695 89.755 191.835 96.235 ;
        RECT 192.155 95.195 192.295 97.255 ;
        RECT 192.095 94.875 192.355 95.195 ;
        RECT 192.615 94.515 192.755 101.675 ;
        RECT 194.915 100.295 195.055 101.675 ;
        RECT 194.855 100.205 195.115 100.295 ;
        RECT 194.455 100.065 195.115 100.205 ;
        RECT 193.475 98.615 193.735 98.935 ;
        RECT 193.535 97.915 193.675 98.615 ;
        RECT 193.475 97.595 193.735 97.915 ;
        RECT 192.555 94.195 192.815 94.515 ;
        RECT 192.095 93.855 192.355 94.175 ;
        RECT 192.155 91.795 192.295 93.855 ;
        RECT 192.555 93.175 192.815 93.495 ;
        RECT 192.095 91.475 192.355 91.795 ;
        RECT 191.635 89.435 191.895 89.755 ;
        RECT 191.695 88.735 191.835 89.435 ;
        RECT 192.615 89.415 192.755 93.175 ;
        RECT 193.475 91.875 193.735 92.135 ;
        RECT 193.475 91.815 194.135 91.875 ;
        RECT 193.535 91.735 194.135 91.815 ;
        RECT 193.015 90.795 193.275 91.115 ;
        RECT 192.555 89.095 192.815 89.415 ;
        RECT 191.635 88.415 191.895 88.735 ;
        RECT 193.075 85.335 193.215 90.795 ;
        RECT 193.995 86.695 194.135 91.735 ;
        RECT 194.455 91.455 194.595 100.065 ;
        RECT 194.855 99.975 195.115 100.065 ;
        RECT 194.855 94.195 195.115 94.515 ;
        RECT 194.915 92.135 195.055 94.195 ;
        RECT 194.855 91.815 195.115 92.135 ;
        RECT 194.395 91.135 194.655 91.455 ;
        RECT 193.935 86.375 194.195 86.695 ;
        RECT 194.455 86.015 194.595 91.135 ;
        RECT 194.855 90.455 195.115 90.775 ;
        RECT 194.395 85.695 194.655 86.015 ;
        RECT 190.255 85.015 190.515 85.335 ;
        RECT 193.015 85.015 193.275 85.335 ;
        RECT 188.875 83.315 189.135 83.635 ;
        RECT 193.075 83.150 193.215 85.015 ;
        RECT 194.915 84.315 195.055 90.455 ;
        RECT 194.855 83.995 195.115 84.315 ;
        RECT 193.475 83.315 193.735 83.635 ;
        RECT 193.005 82.780 193.285 83.150 ;
        RECT 189.335 82.295 189.595 82.615 ;
        RECT 189.395 81.595 189.535 82.295 ;
        RECT 189.335 81.275 189.595 81.595 ;
        RECT 188.875 79.915 189.135 80.235 ;
        RECT 187.955 79.575 188.215 79.895 ;
        RECT 188.415 79.575 188.675 79.895 ;
        RECT 187.035 78.555 187.295 78.875 ;
        RECT 188.015 78.535 188.155 79.575 ;
        RECT 187.955 78.215 188.215 78.535 ;
        RECT 187.495 77.875 187.755 78.195 ;
        RECT 187.555 76.065 187.695 77.875 ;
        RECT 188.475 77.175 188.615 79.575 ;
        RECT 188.935 78.875 189.075 79.915 ;
        RECT 188.875 78.555 189.135 78.875 ;
        RECT 188.415 76.855 188.675 77.175 ;
        RECT 186.175 75.925 187.695 76.065 ;
        RECT 186.175 75.555 186.315 75.925 ;
        RECT 185.715 75.475 186.315 75.555 ;
        RECT 185.655 75.415 186.315 75.475 ;
        RECT 185.655 75.155 185.915 75.415 ;
        RECT 187.035 75.155 187.295 75.475 ;
        RECT 184.725 74.620 185.005 74.990 ;
        RECT 184.795 73.435 184.935 74.620 ;
        RECT 184.735 73.115 184.995 73.435 ;
        RECT 187.095 72.155 187.235 75.155 ;
        RECT 187.555 73.095 187.695 75.925 ;
        RECT 188.475 74.795 188.615 76.855 ;
        RECT 192.095 75.155 192.355 75.475 ;
        RECT 188.415 74.475 188.675 74.795 ;
        RECT 192.155 73.435 192.295 75.155 ;
        RECT 193.535 74.455 193.675 83.315 ;
        RECT 193.935 82.975 194.195 83.295 ;
        RECT 193.995 81.255 194.135 82.975 ;
        RECT 194.395 82.635 194.655 82.955 ;
        RECT 193.935 80.935 194.195 81.255 ;
        RECT 193.475 74.135 193.735 74.455 ;
        RECT 192.095 73.115 192.355 73.435 ;
        RECT 187.495 72.775 187.755 73.095 ;
        RECT 187.095 72.015 188.155 72.155 ;
        RECT 187.495 71.415 187.755 71.735 ;
        RECT 187.555 69.695 187.695 71.415 ;
        RECT 188.015 70.375 188.155 72.015 ;
        RECT 187.955 70.055 188.215 70.375 ;
        RECT 192.155 69.695 192.295 73.115 ;
        RECT 193.535 73.095 193.675 74.135 ;
        RECT 193.475 72.775 193.735 73.095 ;
        RECT 193.995 72.755 194.135 80.935 ;
        RECT 194.455 76.155 194.595 82.635 ;
        RECT 195.375 81.595 195.515 105.075 ;
        RECT 195.315 81.275 195.575 81.595 ;
        RECT 194.855 79.575 195.115 79.895 ;
        RECT 194.915 78.195 195.055 79.575 ;
        RECT 194.855 77.875 195.115 78.195 ;
        RECT 194.395 75.835 194.655 76.155 ;
        RECT 195.375 75.475 195.515 81.275 ;
        RECT 195.315 75.155 195.575 75.475 ;
        RECT 194.385 74.620 194.665 74.990 ;
        RECT 194.455 74.455 194.595 74.620 ;
        RECT 194.395 74.135 194.655 74.455 ;
        RECT 194.855 72.775 195.115 73.095 ;
        RECT 192.555 72.435 192.815 72.755 ;
        RECT 193.935 72.435 194.195 72.755 ;
        RECT 187.495 69.375 187.755 69.695 ;
        RECT 192.095 69.375 192.355 69.695 ;
        RECT 189.795 68.695 190.055 69.015 ;
        RECT 189.855 67.655 189.995 68.695 ;
        RECT 189.795 67.335 190.055 67.655 ;
        RECT 186.115 66.655 186.375 66.975 ;
        RECT 186.175 64.595 186.315 66.655 ;
        RECT 187.495 65.975 187.755 66.295 ;
        RECT 187.555 64.595 187.695 65.975 ;
        RECT 192.615 64.935 192.755 72.435 ;
        RECT 193.475 72.095 193.735 72.415 ;
        RECT 193.535 70.035 193.675 72.095 ;
        RECT 193.475 69.715 193.735 70.035 ;
        RECT 192.555 64.615 192.815 64.935 ;
        RECT 186.115 64.275 186.375 64.595 ;
        RECT 187.495 64.275 187.755 64.595 ;
        RECT 184.275 62.235 184.535 62.555 ;
        RECT 192.095 60.535 192.355 60.855 ;
        RECT 192.555 60.535 192.815 60.855 ;
        RECT 192.155 59.155 192.295 60.535 ;
        RECT 192.615 59.835 192.755 60.535 ;
        RECT 192.555 59.515 192.815 59.835 ;
        RECT 192.095 58.835 192.355 59.155 ;
        RECT 187.955 58.495 188.215 58.815 ;
        RECT 194.395 58.495 194.655 58.815 ;
        RECT 181.515 57.815 181.775 58.135 ;
        RECT 181.975 57.815 182.235 58.135 ;
        RECT 186.115 57.875 186.375 58.135 ;
        RECT 186.115 57.815 186.775 57.875 ;
        RECT 181.575 56.515 181.715 57.815 ;
        RECT 186.175 57.735 186.775 57.815 ;
        RECT 181.575 56.375 182.175 56.515 ;
        RECT 179.955 54.560 181.495 54.930 ;
        RECT 182.035 54.395 182.175 56.375 ;
        RECT 186.635 56.095 186.775 57.735 ;
        RECT 188.015 56.095 188.155 58.495 ;
        RECT 194.455 58.135 194.595 58.495 ;
        RECT 194.395 57.815 194.655 58.135 ;
        RECT 186.575 55.950 186.835 56.095 ;
        RECT 186.565 55.580 186.845 55.950 ;
        RECT 187.955 55.775 188.215 56.095 ;
        RECT 181.975 54.075 182.235 54.395 ;
        RECT 178.745 52.975 179.415 53.115 ;
        RECT 178.745 52.860 179.025 52.975 ;
        RECT 188.015 51.335 188.155 55.775 ;
        RECT 194.915 53.035 195.055 72.775 ;
        RECT 195.835 71.735 195.975 105.075 ;
        RECT 196.755 78.535 196.895 105.415 ;
        RECT 197.215 93.495 197.355 105.415 ;
        RECT 199.975 103.355 200.115 105.415 ;
        RECT 203.195 104.715 203.335 109.225 ;
        RECT 203.595 105.075 203.855 105.395 ;
        RECT 204.515 105.075 204.775 105.395 ;
        RECT 203.135 104.395 203.395 104.715 ;
        RECT 202.675 104.055 202.935 104.375 ;
        RECT 199.915 103.035 200.175 103.355 ;
        RECT 199.975 102.075 200.115 103.035 ;
        RECT 202.735 102.335 202.875 104.055 ;
        RECT 199.975 101.935 200.575 102.075 ;
        RECT 200.835 102.015 201.095 102.335 ;
        RECT 202.675 102.015 202.935 102.335 ;
        RECT 203.135 102.015 203.395 102.335 ;
        RECT 198.585 100.800 200.125 101.170 ;
        RECT 200.435 100.635 200.575 101.935 ;
        RECT 200.375 100.315 200.635 100.635 ;
        RECT 198.985 99.780 199.265 100.150 ;
        RECT 198.995 99.635 199.255 99.780 ;
        RECT 197.615 98.615 197.875 98.935 ;
        RECT 198.995 98.615 199.255 98.935 ;
        RECT 197.675 96.555 197.815 98.615 ;
        RECT 198.065 97.060 198.345 97.430 ;
        RECT 199.055 97.235 199.195 98.615 ;
        RECT 198.075 96.915 198.335 97.060 ;
        RECT 198.995 96.915 199.255 97.235 ;
        RECT 197.615 96.235 197.875 96.555 ;
        RECT 197.155 93.175 197.415 93.495 ;
        RECT 197.215 90.775 197.355 93.175 ;
        RECT 198.135 91.705 198.275 96.915 ;
        RECT 200.375 95.895 200.635 96.215 ;
        RECT 198.585 95.360 200.125 95.730 ;
        RECT 200.435 94.855 200.575 95.895 ;
        RECT 200.375 94.535 200.635 94.855 ;
        RECT 198.135 91.565 198.735 91.705 ;
        RECT 198.595 91.115 198.735 91.565 ;
        RECT 198.075 90.795 198.335 91.115 ;
        RECT 198.535 90.795 198.795 91.115 ;
        RECT 197.155 90.455 197.415 90.775 ;
        RECT 197.215 88.735 197.355 90.455 ;
        RECT 198.135 89.755 198.275 90.795 ;
        RECT 198.585 89.920 200.125 90.290 ;
        RECT 198.075 89.435 198.335 89.755 ;
        RECT 200.895 88.735 201.035 102.015 ;
        RECT 201.295 98.615 201.555 98.935 ;
        RECT 201.355 95.195 201.495 98.615 ;
        RECT 202.215 97.595 202.475 97.915 ;
        RECT 202.275 96.895 202.415 97.595 ;
        RECT 203.195 97.315 203.335 102.015 ;
        RECT 203.655 97.575 203.795 105.075 ;
        RECT 202.735 97.175 203.335 97.315 ;
        RECT 203.595 97.255 203.855 97.575 ;
        RECT 201.755 96.575 202.015 96.895 ;
        RECT 202.215 96.575 202.475 96.895 ;
        RECT 201.295 94.875 201.555 95.195 ;
        RECT 201.815 94.855 201.955 96.575 ;
        RECT 202.735 96.125 202.875 97.175 ;
        RECT 203.135 96.575 203.395 96.895 ;
        RECT 202.275 95.985 202.875 96.125 ;
        RECT 201.755 94.535 202.015 94.855 ;
        RECT 201.295 91.135 201.555 91.455 ;
        RECT 197.155 88.415 197.415 88.735 ;
        RECT 200.835 88.415 201.095 88.735 ;
        RECT 200.895 87.035 201.035 88.415 ;
        RECT 200.835 86.715 201.095 87.035 ;
        RECT 198.585 84.480 200.125 84.850 ;
        RECT 200.895 83.975 201.035 86.715 ;
        RECT 200.835 83.655 201.095 83.975 ;
        RECT 200.825 80.060 201.105 80.430 ;
        RECT 198.585 79.040 200.125 79.410 ;
        RECT 200.895 78.875 201.035 80.060 ;
        RECT 200.835 78.555 201.095 78.875 ;
        RECT 196.695 78.215 196.955 78.535 ;
        RECT 196.755 77.175 196.895 78.215 ;
        RECT 197.155 77.535 197.415 77.855 ;
        RECT 196.695 76.855 196.955 77.175 ;
        RECT 197.215 76.235 197.355 77.535 ;
        RECT 200.835 76.855 201.095 77.175 ;
        RECT 196.235 75.835 196.495 76.155 ;
        RECT 196.755 76.095 197.355 76.235 ;
        RECT 200.895 76.155 201.035 76.855 ;
        RECT 195.305 71.220 195.585 71.590 ;
        RECT 195.775 71.415 196.035 71.735 ;
        RECT 195.375 69.695 195.515 71.220 ;
        RECT 196.295 70.715 196.435 75.835 ;
        RECT 196.755 75.815 196.895 76.095 ;
        RECT 200.835 75.835 201.095 76.155 ;
        RECT 196.695 75.495 196.955 75.815 ;
        RECT 196.235 70.395 196.495 70.715 ;
        RECT 195.315 69.375 195.575 69.695 ;
        RECT 196.295 67.655 196.435 70.395 ;
        RECT 196.755 70.035 196.895 75.495 ;
        RECT 200.375 74.815 200.635 75.135 ;
        RECT 197.155 74.135 197.415 74.455 ;
        RECT 198.075 74.135 198.335 74.455 ;
        RECT 197.215 73.435 197.355 74.135 ;
        RECT 197.155 73.115 197.415 73.435 ;
        RECT 198.135 72.415 198.275 74.135 ;
        RECT 198.585 73.600 200.125 73.970 ;
        RECT 198.075 72.095 198.335 72.415 ;
        RECT 197.615 71.415 197.875 71.735 ;
        RECT 197.675 70.035 197.815 71.415 ;
        RECT 200.435 70.625 200.575 74.815 ;
        RECT 200.895 72.755 201.035 75.835 ;
        RECT 201.355 75.135 201.495 91.135 ;
        RECT 202.275 83.035 202.415 95.985 ;
        RECT 203.195 94.515 203.335 96.575 ;
        RECT 203.655 96.070 203.795 97.255 ;
        RECT 203.585 95.700 203.865 96.070 ;
        RECT 203.135 94.195 203.395 94.515 ;
        RECT 202.675 90.455 202.935 90.775 ;
        RECT 202.735 89.755 202.875 90.455 ;
        RECT 202.675 89.435 202.935 89.755 ;
        RECT 203.195 86.015 203.335 94.195 ;
        RECT 204.575 92.135 204.715 105.075 ;
        RECT 205.495 103.355 205.635 109.225 ;
        RECT 207.795 106.075 207.935 109.225 ;
        RECT 207.735 105.755 207.995 106.075 ;
        RECT 209.575 104.735 209.835 105.055 ;
        RECT 205.435 103.035 205.695 103.355 ;
        RECT 205.435 102.355 205.695 102.675 ;
        RECT 205.495 100.635 205.635 102.355 ;
        RECT 209.115 101.675 209.375 101.995 ;
        RECT 205.435 100.315 205.695 100.635 ;
        RECT 209.175 100.295 209.315 101.675 ;
        RECT 209.115 99.975 209.375 100.295 ;
        RECT 205.425 99.100 205.705 99.470 ;
        RECT 205.495 96.555 205.635 99.100 ;
        RECT 206.355 98.615 206.615 98.935 ;
        RECT 206.415 96.555 206.555 98.615 ;
        RECT 207.735 97.595 207.995 97.915 ;
        RECT 207.795 96.895 207.935 97.595 ;
        RECT 207.735 96.575 207.995 96.895 ;
        RECT 205.435 96.235 205.695 96.555 ;
        RECT 206.355 96.235 206.615 96.555 ;
        RECT 204.965 93.660 205.245 94.030 ;
        RECT 204.515 91.815 204.775 92.135 ;
        RECT 204.575 91.455 204.715 91.815 ;
        RECT 204.515 91.135 204.775 91.455 ;
        RECT 204.575 89.755 204.715 91.135 ;
        RECT 205.035 91.115 205.175 93.660 ;
        RECT 207.795 91.455 207.935 96.575 ;
        RECT 208.195 95.895 208.455 96.215 ;
        RECT 208.655 95.895 208.915 96.215 ;
        RECT 208.255 95.390 208.395 95.895 ;
        RECT 208.185 95.020 208.465 95.390 ;
        RECT 208.715 94.515 208.855 95.895 ;
        RECT 208.655 94.195 208.915 94.515 ;
        RECT 208.195 93.515 208.455 93.835 ;
        RECT 207.735 91.135 207.995 91.455 ;
        RECT 204.975 90.795 205.235 91.115 ;
        RECT 204.515 89.435 204.775 89.755 ;
        RECT 206.355 88.415 206.615 88.735 ;
        RECT 206.415 86.015 206.555 88.415 ;
        RECT 207.795 87.035 207.935 91.135 ;
        RECT 208.255 89.075 208.395 93.515 ;
        RECT 208.715 91.795 208.855 94.195 ;
        RECT 209.175 93.835 209.315 99.975 ;
        RECT 209.635 97.575 209.775 104.735 ;
        RECT 210.095 103.355 210.235 109.225 ;
        RECT 212.395 106.075 212.535 109.225 ;
        RECT 214.695 106.075 214.835 109.225 ;
        RECT 211.415 105.755 211.675 106.075 ;
        RECT 212.335 105.755 212.595 106.075 ;
        RECT 214.635 105.755 214.895 106.075 ;
        RECT 210.035 103.035 210.295 103.355 ;
        RECT 211.475 99.955 211.615 105.755 ;
        RECT 212.795 105.075 213.055 105.395 ;
        RECT 213.255 105.075 213.515 105.395 ;
        RECT 214.175 105.075 214.435 105.395 ;
        RECT 212.855 103.015 212.995 105.075 ;
        RECT 212.795 102.695 213.055 103.015 ;
        RECT 211.415 99.635 211.675 99.955 ;
        RECT 211.875 99.635 212.135 99.955 ;
        RECT 209.575 97.255 209.835 97.575 ;
        RECT 211.475 97.315 211.615 99.635 ;
        RECT 211.935 97.915 212.075 99.635 ;
        RECT 211.875 97.595 212.135 97.915 ;
        RECT 210.035 96.915 210.295 97.235 ;
        RECT 211.475 97.175 212.075 97.315 ;
        RECT 209.115 93.515 209.375 93.835 ;
        RECT 209.115 92.155 209.375 92.475 ;
        RECT 208.655 91.475 208.915 91.795 ;
        RECT 208.715 89.270 208.855 91.475 ;
        RECT 208.195 88.755 208.455 89.075 ;
        RECT 208.645 88.900 208.925 89.270 ;
        RECT 209.175 89.075 209.315 92.155 ;
        RECT 209.575 91.475 209.835 91.795 ;
        RECT 209.115 88.755 209.375 89.075 ;
        RECT 207.735 86.715 207.995 87.035 ;
        RECT 203.135 85.695 203.395 86.015 ;
        RECT 206.355 85.695 206.615 86.015 ;
        RECT 206.815 85.695 207.075 86.015 ;
        RECT 202.665 83.035 202.945 83.150 ;
        RECT 202.275 82.895 202.945 83.035 ;
        RECT 202.665 82.780 202.945 82.895 ;
        RECT 202.215 77.535 202.475 77.855 ;
        RECT 201.295 74.815 201.555 75.135 ;
        RECT 200.835 72.435 201.095 72.755 ;
        RECT 200.835 71.415 201.095 71.735 ;
        RECT 199.515 70.485 200.575 70.625 ;
        RECT 196.695 69.715 196.955 70.035 ;
        RECT 197.615 69.715 197.875 70.035 ;
        RECT 197.155 69.035 197.415 69.355 ;
        RECT 196.695 68.695 196.955 69.015 ;
        RECT 196.235 67.335 196.495 67.655 ;
        RECT 196.295 64.255 196.435 67.335 ;
        RECT 196.755 66.635 196.895 68.695 ;
        RECT 197.215 67.655 197.355 69.035 ;
        RECT 199.515 68.925 199.655 70.485 ;
        RECT 199.905 70.115 200.185 70.230 ;
        RECT 199.905 69.975 200.575 70.115 ;
        RECT 199.905 69.860 200.185 69.975 ;
        RECT 199.915 68.925 200.175 69.015 ;
        RECT 199.515 68.785 200.175 68.925 ;
        RECT 199.915 68.695 200.175 68.785 ;
        RECT 198.585 68.160 200.125 68.530 ;
        RECT 200.435 67.995 200.575 69.975 ;
        RECT 200.375 67.675 200.635 67.995 ;
        RECT 197.155 67.335 197.415 67.655 ;
        RECT 200.435 67.395 200.575 67.675 ;
        RECT 200.895 67.655 201.035 71.415 ;
        RECT 201.285 71.220 201.565 71.590 ;
        RECT 201.355 70.375 201.495 71.220 ;
        RECT 201.755 70.395 202.015 70.715 ;
        RECT 201.295 70.055 201.555 70.375 ;
        RECT 201.815 69.695 201.955 70.395 ;
        RECT 202.275 70.035 202.415 77.535 ;
        RECT 202.675 72.270 202.935 72.415 ;
        RECT 202.665 71.900 202.945 72.270 ;
        RECT 202.215 69.715 202.475 70.035 ;
        RECT 201.755 69.375 202.015 69.695 ;
        RECT 202.675 67.675 202.935 67.995 ;
        RECT 199.975 67.255 200.575 67.395 ;
        RECT 200.835 67.335 201.095 67.655 ;
        RECT 201.295 67.335 201.555 67.655 ;
        RECT 199.975 66.975 200.115 67.255 ;
        RECT 199.915 66.655 200.175 66.975 ;
        RECT 200.375 66.715 200.635 66.975 ;
        RECT 201.355 66.715 201.495 67.335 ;
        RECT 200.375 66.655 201.495 66.715 ;
        RECT 196.695 66.315 196.955 66.635 ;
        RECT 200.435 66.575 201.495 66.655 ;
        RECT 196.755 64.935 196.895 66.315 ;
        RECT 197.615 65.975 197.875 66.295 ;
        RECT 197.675 65.275 197.815 65.975 ;
        RECT 197.615 64.955 197.875 65.275 ;
        RECT 196.695 64.615 196.955 64.935 ;
        RECT 200.435 64.595 200.575 66.575 ;
        RECT 200.375 64.275 200.635 64.595 ;
        RECT 196.235 63.935 196.495 64.255 ;
        RECT 197.615 63.255 197.875 63.575 ;
        RECT 197.675 61.535 197.815 63.255 ;
        RECT 198.585 62.720 200.125 63.090 ;
        RECT 198.075 61.555 198.335 61.875 ;
        RECT 197.615 61.215 197.875 61.535 ;
        RECT 195.775 57.815 196.035 58.135 ;
        RECT 195.835 57.115 195.975 57.815 ;
        RECT 197.675 57.115 197.815 61.215 ;
        RECT 198.135 59.835 198.275 61.555 ;
        RECT 202.735 61.195 202.875 67.675 ;
        RECT 202.675 60.875 202.935 61.195 ;
        RECT 198.075 59.515 198.335 59.835 ;
        RECT 202.675 58.495 202.935 58.815 ;
        RECT 198.075 58.155 198.335 58.475 ;
        RECT 195.775 56.795 196.035 57.115 ;
        RECT 197.615 56.795 197.875 57.115 ;
        RECT 198.135 56.435 198.275 58.155 ;
        RECT 198.585 57.280 200.125 57.650 ;
        RECT 202.735 57.115 202.875 58.495 ;
        RECT 202.675 56.795 202.935 57.115 ;
        RECT 198.075 56.115 198.335 56.435 ;
        RECT 200.375 56.115 200.635 56.435 ;
        RECT 190.255 52.715 190.515 53.035 ;
        RECT 194.855 52.715 195.115 53.035 ;
        RECT 187.955 51.015 188.215 51.335 ;
        RECT 179.955 49.120 181.495 49.490 ;
        RECT 146.290 43.995 148.395 48.095 ;
        RECT 177.375 47.955 177.635 48.275 ;
        RECT 186.115 47.275 186.375 47.595 ;
        RECT 189.795 47.275 190.055 47.595 ;
        RECT 181.975 46.935 182.235 47.255 ;
        RECT 176.455 44.895 176.715 45.215 ;
        RECT 178.755 44.895 179.015 45.215 ;
        RECT 179.215 44.895 179.475 45.215 ;
        RECT 173.695 44.215 173.955 44.535 ;
        RECT 173.755 43.515 173.895 44.215 ;
        RECT 176.515 43.515 176.655 44.895 ;
        RECT 177.375 44.215 177.635 44.535 ;
        RECT 143.435 41.655 145.540 42.245 ;
        RECT 143.835 41.605 145.135 41.655 ;
        RECT 7.065 36.430 8.665 39.630 ;
        RECT 10.170 37.965 74.550 38.965 ;
        RECT 79.810 38.185 127.975 39.285 ;
        RECT 10.170 35.440 74.550 36.940 ;
        RECT 79.810 36.685 127.975 37.785 ;
        RECT 79.810 35.185 127.975 36.285 ;
        RECT 136.295 35.805 138.400 39.905 ;
        RECT 146.290 38.145 148.395 43.415 ;
        RECT 173.695 43.195 173.955 43.515 ;
        RECT 176.455 43.195 176.715 43.515 ;
        RECT 176.915 42.515 177.175 42.835 ;
        RECT 173.695 42.175 173.955 42.495 ;
        RECT 170.015 41.495 170.275 41.815 ;
        RECT 170.075 40.795 170.215 41.495 ;
        RECT 173.755 40.795 173.895 42.175 ;
        RECT 170.015 40.475 170.275 40.795 ;
        RECT 173.695 40.475 173.955 40.795 ;
        RECT 165.875 38.775 166.135 39.095 ;
        RECT 10.170 33.440 74.550 34.940 ;
        RECT 79.810 33.685 127.975 34.785 ;
        RECT 10.170 31.440 74.550 32.940 ;
        RECT 79.810 32.185 127.975 33.285 ;
        RECT 79.810 30.685 127.975 31.785 ;
        RECT 136.295 31.125 138.400 35.225 ;
        RECT 146.290 33.465 148.395 37.565 ;
        RECT 165.935 37.055 166.075 38.775 ;
        RECT 176.975 37.395 177.115 42.515 ;
        RECT 176.915 37.075 177.175 37.395 ;
        RECT 165.875 36.735 166.135 37.055 ;
        RECT 165.935 35.355 166.075 36.735 ;
        RECT 167.255 36.395 167.515 36.715 ;
        RECT 165.875 35.035 166.135 35.355 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 167.315 32.635 167.455 36.395 ;
        RECT 177.435 35.355 177.575 44.215 ;
        RECT 178.815 43.515 178.955 44.895 ;
        RECT 178.755 43.195 179.015 43.515 ;
        RECT 179.275 42.915 179.415 44.895 ;
        RECT 179.955 43.680 181.495 44.050 ;
        RECT 182.035 43.515 182.175 46.935 ;
        RECT 186.175 45.555 186.315 47.275 ;
        RECT 186.115 45.235 186.375 45.555 ;
        RECT 184.275 44.275 184.535 44.535 ;
        RECT 183.875 44.215 184.535 44.275 ;
        RECT 183.875 44.135 184.475 44.215 ;
        RECT 181.975 43.195 182.235 43.515 ;
        RECT 178.355 42.775 179.415 42.915 ;
        RECT 177.835 41.495 178.095 41.815 ;
        RECT 177.895 40.795 178.035 41.495 ;
        RECT 177.835 40.475 178.095 40.795 ;
        RECT 178.355 39.775 178.495 42.775 ;
        RECT 178.755 42.175 179.015 42.495 ;
        RECT 178.295 39.455 178.555 39.775 ;
        RECT 178.355 37.475 178.495 39.455 ;
        RECT 177.895 37.335 178.495 37.475 ;
        RECT 178.815 37.395 178.955 42.175 ;
        RECT 179.275 40.795 179.415 42.775 ;
        RECT 183.875 42.495 184.015 44.135 ;
        RECT 183.815 42.175 184.075 42.495 ;
        RECT 179.675 41.835 179.935 42.155 ;
        RECT 179.735 40.795 179.875 41.835 ;
        RECT 189.855 41.815 189.995 47.275 ;
        RECT 190.315 44.535 190.455 52.715 ;
        RECT 194.915 51.335 195.055 52.715 ;
        RECT 198.585 51.840 200.125 52.210 ;
        RECT 190.715 51.015 190.975 51.335 ;
        RECT 194.855 51.015 195.115 51.335 ;
        RECT 190.775 47.935 190.915 51.015 ;
        RECT 193.015 49.995 193.275 50.315 ;
        RECT 190.715 47.615 190.975 47.935 ;
        RECT 193.075 45.895 193.215 49.995 ;
        RECT 193.475 47.955 193.735 48.275 ;
        RECT 193.535 46.235 193.675 47.955 ;
        RECT 200.435 47.595 200.575 56.115 ;
        RECT 202.215 53.735 202.475 54.055 ;
        RECT 201.295 53.055 201.555 53.375 ;
        RECT 200.835 52.375 201.095 52.695 ;
        RECT 200.895 50.315 201.035 52.375 ;
        RECT 201.355 50.655 201.495 53.055 ;
        RECT 202.275 52.435 202.415 53.735 ;
        RECT 202.675 52.435 202.935 52.695 ;
        RECT 202.275 52.375 202.935 52.435 ;
        RECT 202.275 52.295 202.875 52.375 ;
        RECT 201.295 50.395 201.555 50.655 ;
        RECT 201.295 50.335 201.955 50.395 ;
        RECT 200.835 49.995 201.095 50.315 ;
        RECT 201.355 50.255 201.955 50.335 ;
        RECT 200.375 47.275 200.635 47.595 ;
        RECT 198.585 46.400 200.125 46.770 ;
        RECT 193.475 45.915 193.735 46.235 ;
        RECT 193.015 45.575 193.275 45.895 ;
        RECT 195.315 45.235 195.575 45.555 ;
        RECT 190.715 44.895 190.975 45.215 ;
        RECT 195.375 44.955 195.515 45.235 ;
        RECT 190.255 44.215 190.515 44.535 ;
        RECT 190.315 42.495 190.455 44.215 ;
        RECT 190.775 43.515 190.915 44.895 ;
        RECT 195.375 44.815 196.895 44.955 ;
        RECT 198.075 44.895 198.335 45.215 ;
        RECT 190.715 43.195 190.975 43.515 ;
        RECT 190.255 42.175 190.515 42.495 ;
        RECT 189.795 41.495 190.055 41.815 ;
        RECT 179.215 40.475 179.475 40.795 ;
        RECT 179.675 40.475 179.935 40.795 ;
        RECT 179.735 39.515 179.875 40.475 ;
        RECT 187.495 39.795 187.755 40.115 ;
        RECT 179.275 39.375 179.875 39.515 ;
        RECT 185.655 39.455 185.915 39.775 ;
        RECT 177.895 36.715 178.035 37.335 ;
        RECT 178.755 37.075 179.015 37.395 ;
        RECT 177.835 36.395 178.095 36.715 ;
        RECT 178.295 36.395 178.555 36.715 ;
        RECT 177.375 35.035 177.635 35.355 ;
        RECT 177.895 35.015 178.035 36.395 ;
        RECT 178.355 35.355 178.495 36.395 ;
        RECT 179.275 35.355 179.415 39.375 ;
        RECT 179.955 38.240 181.495 38.610 ;
        RECT 185.715 37.735 185.855 39.455 ;
        RECT 187.555 38.075 187.695 39.795 ;
        RECT 190.315 39.775 190.455 42.175 ;
        RECT 196.755 42.155 196.895 44.815 ;
        RECT 197.155 44.555 197.415 44.875 ;
        RECT 197.215 43.515 197.355 44.555 ;
        RECT 197.155 43.195 197.415 43.515 ;
        RECT 191.635 41.835 191.895 42.155 ;
        RECT 196.695 41.835 196.955 42.155 ;
        RECT 191.695 40.795 191.835 41.835 ;
        RECT 191.635 40.475 191.895 40.795 ;
        RECT 192.095 39.795 192.355 40.115 ;
        RECT 190.255 39.455 190.515 39.775 ;
        RECT 189.795 38.775 190.055 39.095 ;
        RECT 187.495 37.755 187.755 38.075 ;
        RECT 185.655 37.415 185.915 37.735 ;
        RECT 179.675 37.075 179.935 37.395 ;
        RECT 178.295 35.035 178.555 35.355 ;
        RECT 179.215 35.035 179.475 35.355 ;
        RECT 177.835 34.695 178.095 35.015 ;
        RECT 168.635 34.015 168.895 34.335 ;
        RECT 168.695 32.635 168.835 34.015 ;
        RECT 176.455 33.335 176.715 33.655 ;
        RECT 167.255 32.315 167.515 32.635 ;
        RECT 168.635 32.315 168.895 32.635 ;
        RECT 176.515 31.955 176.655 33.335 ;
        RECT 176.455 31.635 176.715 31.955 ;
        RECT 178.355 31.275 178.495 35.035 ;
        RECT 179.735 34.245 179.875 37.075 ;
        RECT 183.355 36.735 183.615 37.055 ;
        RECT 183.415 35.355 183.555 36.735 ;
        RECT 189.855 36.715 189.995 38.775 ;
        RECT 190.315 37.395 190.455 39.455 ;
        RECT 190.255 37.075 190.515 37.395 ;
        RECT 189.795 36.395 190.055 36.715 ;
        RECT 183.355 35.035 183.615 35.355 ;
        RECT 180.135 34.245 180.395 34.335 ;
        RECT 179.735 34.105 180.395 34.245 ;
        RECT 180.135 34.015 180.395 34.105 ;
        RECT 178.755 33.675 179.015 33.995 ;
        RECT 178.815 32.635 178.955 33.675 ;
        RECT 179.955 32.800 181.495 33.170 ;
        RECT 178.755 32.315 179.015 32.635 ;
        RECT 190.315 31.955 190.455 37.075 ;
        RECT 192.155 35.355 192.295 39.795 ;
        RECT 194.855 39.455 195.115 39.775 ;
        RECT 194.915 36.375 195.055 39.455 ;
        RECT 194.855 36.115 195.115 36.375 ;
        RECT 194.455 36.055 195.115 36.115 ;
        RECT 194.455 35.975 195.055 36.055 ;
        RECT 192.095 35.035 192.355 35.355 ;
        RECT 190.715 34.355 190.975 34.675 ;
        RECT 187.035 31.635 187.295 31.955 ;
        RECT 190.255 31.635 190.515 31.955 ;
        RECT 178.295 30.955 178.555 31.275 ;
        RECT 10.170 28.035 74.550 30.415 ;
        RECT 79.810 28.165 127.975 30.285 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 187.095 29.915 187.235 31.635 ;
        RECT 187.035 29.595 187.295 29.915 ;
        RECT 190.315 29.575 190.455 31.635 ;
        RECT 190.775 30.935 190.915 34.355 ;
        RECT 191.635 33.675 191.895 33.995 ;
        RECT 190.715 30.615 190.975 30.935 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 190.255 29.255 190.515 29.575 ;
        RECT 186.115 28.915 186.375 29.235 ;
        RECT 164.035 28.070 164.295 28.215 ;
        RECT 10.170 25.510 74.550 27.010 ;
        RECT 79.810 26.665 127.975 27.765 ;
        RECT 164.025 27.700 164.305 28.070 ;
        RECT 179.955 27.360 181.495 27.730 ;
        RECT 186.175 27.195 186.315 28.915 ;
        RECT 190.255 27.895 190.515 28.215 ;
        RECT 186.115 26.875 186.375 27.195 ;
        RECT 79.810 25.165 127.975 26.265 ;
        RECT 190.315 26.175 190.455 27.895 ;
        RECT 190.775 26.515 190.915 30.615 ;
        RECT 191.695 26.515 191.835 33.675 ;
        RECT 193.935 33.335 194.195 33.655 ;
        RECT 193.995 32.635 194.135 33.335 ;
        RECT 193.935 32.315 194.195 32.635 ;
        RECT 193.015 31.635 193.275 31.955 ;
        RECT 193.075 29.915 193.215 31.635 ;
        RECT 194.455 29.915 194.595 35.975 ;
        RECT 194.855 34.355 195.115 34.675 ;
        RECT 194.915 29.915 195.055 34.355 ;
        RECT 195.315 34.015 195.575 34.335 ;
        RECT 193.015 29.595 193.275 29.915 ;
        RECT 194.395 29.595 194.655 29.915 ;
        RECT 194.855 29.595 195.115 29.915 ;
        RECT 195.375 28.895 195.515 34.015 ;
        RECT 196.755 31.275 196.895 41.835 ;
        RECT 198.135 39.095 198.275 44.895 ;
        RECT 198.585 40.960 200.125 41.330 ;
        RECT 198.075 38.775 198.335 39.095 ;
        RECT 197.615 36.735 197.875 37.055 ;
        RECT 197.675 32.635 197.815 36.735 ;
        RECT 198.135 35.015 198.275 38.775 ;
        RECT 200.435 36.715 200.575 47.275 ;
        RECT 200.895 42.155 201.035 49.995 ;
        RECT 201.295 49.655 201.555 49.975 ;
        RECT 201.355 45.215 201.495 49.655 ;
        RECT 201.815 48.955 201.955 50.255 ;
        RECT 202.275 49.975 202.415 52.295 ;
        RECT 203.195 51.675 203.335 85.695 ;
        RECT 204.515 85.355 204.775 85.675 ;
        RECT 204.055 72.095 204.315 72.415 ;
        RECT 203.585 70.540 203.865 70.910 ;
        RECT 203.655 69.695 203.795 70.540 ;
        RECT 204.115 69.695 204.255 72.095 ;
        RECT 203.595 69.375 203.855 69.695 ;
        RECT 204.055 69.375 204.315 69.695 ;
        RECT 204.115 67.995 204.255 69.375 ;
        RECT 204.055 67.675 204.315 67.995 ;
        RECT 204.055 66.995 204.315 67.315 ;
        RECT 203.595 63.935 203.855 64.255 ;
        RECT 203.655 62.215 203.795 63.935 ;
        RECT 204.115 63.575 204.255 66.995 ;
        RECT 204.055 63.255 204.315 63.575 ;
        RECT 203.595 61.895 203.855 62.215 ;
        RECT 203.655 59.155 203.795 61.895 ;
        RECT 204.575 61.875 204.715 85.355 ;
        RECT 206.415 78.535 206.555 85.695 ;
        RECT 206.355 78.215 206.615 78.535 ;
        RECT 206.875 78.195 207.015 85.695 ;
        RECT 207.795 83.830 207.935 86.715 ;
        RECT 207.725 83.460 208.005 83.830 ;
        RECT 206.815 77.875 207.075 78.195 ;
        RECT 205.895 77.195 206.155 77.515 ;
        RECT 205.435 72.435 205.695 72.755 ;
        RECT 205.495 69.015 205.635 72.435 ;
        RECT 205.435 68.695 205.695 69.015 ;
        RECT 204.975 66.655 205.235 66.975 ;
        RECT 204.515 61.555 204.775 61.875 ;
        RECT 204.055 60.875 204.315 61.195 ;
        RECT 203.595 58.835 203.855 59.155 ;
        RECT 204.115 53.375 204.255 60.875 ;
        RECT 205.035 58.815 205.175 66.655 ;
        RECT 205.495 61.535 205.635 68.695 ;
        RECT 205.955 66.975 206.095 77.195 ;
        RECT 207.275 72.435 207.535 72.755 ;
        RECT 207.335 69.695 207.475 72.435 ;
        RECT 208.255 70.375 208.395 88.755 ;
        RECT 208.645 86.860 208.925 87.230 ;
        RECT 208.655 86.715 208.915 86.860 ;
        RECT 208.655 85.925 208.915 86.015 ;
        RECT 209.175 85.925 209.315 88.755 ;
        RECT 208.655 85.785 209.315 85.925 ;
        RECT 208.655 85.695 208.915 85.785 ;
        RECT 209.115 85.015 209.375 85.335 ;
        RECT 209.175 83.635 209.315 85.015 ;
        RECT 209.115 83.315 209.375 83.635 ;
        RECT 209.635 78.785 209.775 91.475 ;
        RECT 209.175 78.645 209.775 78.785 ;
        RECT 208.655 77.875 208.915 78.195 ;
        RECT 208.715 76.155 208.855 77.875 ;
        RECT 208.655 75.835 208.915 76.155 ;
        RECT 209.175 75.135 209.315 78.645 ;
        RECT 210.095 78.195 210.235 96.915 ;
        RECT 210.485 95.020 210.765 95.390 ;
        RECT 210.555 81.595 210.695 95.020 ;
        RECT 210.945 93.660 211.225 94.030 ;
        RECT 211.015 84.315 211.155 93.660 ;
        RECT 211.415 88.755 211.675 89.075 ;
        RECT 210.955 83.995 211.215 84.315 ;
        RECT 210.495 81.275 210.755 81.595 ;
        RECT 211.475 80.995 211.615 88.755 ;
        RECT 211.935 84.315 212.075 97.175 ;
        RECT 211.875 83.995 212.135 84.315 ;
        RECT 213.315 83.715 213.455 105.075 ;
        RECT 213.715 93.515 213.975 93.835 ;
        RECT 213.775 91.115 213.915 93.515 ;
        RECT 213.715 90.795 213.975 91.115 ;
        RECT 213.775 89.755 213.915 90.795 ;
        RECT 213.715 89.435 213.975 89.755 ;
        RECT 213.315 83.575 213.915 83.715 ;
        RECT 212.795 82.975 213.055 83.295 ;
        RECT 213.255 82.975 213.515 83.295 ;
        RECT 210.555 80.855 211.615 80.995 ;
        RECT 209.575 77.875 209.835 78.195 ;
        RECT 210.035 77.875 210.295 78.195 ;
        RECT 209.115 74.815 209.375 75.135 ;
        RECT 208.195 70.055 208.455 70.375 ;
        RECT 208.655 70.055 208.915 70.375 ;
        RECT 207.275 69.375 207.535 69.695 ;
        RECT 207.735 69.035 207.995 69.355 ;
        RECT 207.275 66.995 207.535 67.315 ;
        RECT 205.895 66.655 206.155 66.975 ;
        RECT 206.815 64.615 207.075 64.935 ;
        RECT 206.875 63.915 207.015 64.615 ;
        RECT 206.815 63.595 207.075 63.915 ;
        RECT 206.875 62.555 207.015 63.595 ;
        RECT 205.895 62.235 206.155 62.555 ;
        RECT 206.815 62.235 207.075 62.555 ;
        RECT 205.435 61.215 205.695 61.535 ;
        RECT 205.955 61.195 206.095 62.235 ;
        RECT 205.895 60.875 206.155 61.195 ;
        RECT 207.335 59.495 207.475 66.995 ;
        RECT 207.795 65.275 207.935 69.035 ;
        RECT 208.195 67.225 208.455 67.315 ;
        RECT 208.715 67.225 208.855 70.055 ;
        RECT 209.175 70.035 209.315 74.815 ;
        RECT 209.115 69.715 209.375 70.035 ;
        RECT 209.175 67.995 209.315 69.715 ;
        RECT 209.635 69.695 209.775 77.875 ;
        RECT 210.095 74.455 210.235 77.875 ;
        RECT 210.035 74.135 210.295 74.455 ;
        RECT 210.555 70.375 210.695 80.855 ;
        RECT 211.875 80.255 212.135 80.575 ;
        RECT 210.955 77.535 211.215 77.855 ;
        RECT 210.495 70.055 210.755 70.375 ;
        RECT 209.575 69.375 209.835 69.695 ;
        RECT 209.635 67.995 209.775 69.375 ;
        RECT 209.115 67.675 209.375 67.995 ;
        RECT 209.575 67.675 209.835 67.995 ;
        RECT 210.035 67.565 210.295 67.655 ;
        RECT 210.035 67.425 210.695 67.565 ;
        RECT 210.035 67.335 210.295 67.425 ;
        RECT 208.195 67.085 208.855 67.225 ;
        RECT 208.195 66.995 208.455 67.085 ;
        RECT 209.115 66.995 209.375 67.315 ;
        RECT 207.735 64.955 207.995 65.275 ;
        RECT 208.255 64.255 208.395 66.995 ;
        RECT 209.175 66.715 209.315 66.995 ;
        RECT 208.715 66.575 209.315 66.715 ;
        RECT 208.715 65.275 208.855 66.575 ;
        RECT 208.655 64.955 208.915 65.275 ;
        RECT 208.715 64.595 208.855 64.955 ;
        RECT 208.655 64.275 208.915 64.595 ;
        RECT 208.195 63.935 208.455 64.255 ;
        RECT 208.715 63.915 208.855 64.275 ;
        RECT 208.655 63.595 208.915 63.915 ;
        RECT 208.715 60.855 208.855 63.595 ;
        RECT 210.555 63.430 210.695 67.425 ;
        RECT 211.015 67.315 211.155 77.535 ;
        RECT 211.935 75.475 212.075 80.255 ;
        RECT 211.875 75.155 212.135 75.475 ;
        RECT 211.875 71.415 212.135 71.735 ;
        RECT 211.935 69.355 212.075 71.415 ;
        RECT 211.875 69.035 212.135 69.355 ;
        RECT 210.955 66.995 211.215 67.315 ;
        RECT 212.335 66.995 212.595 67.315 ;
        RECT 210.485 63.060 210.765 63.430 ;
        RECT 211.015 60.855 211.155 66.995 ;
        RECT 211.875 64.615 212.135 64.935 ;
        RECT 212.395 64.790 212.535 66.995 ;
        RECT 208.655 60.535 208.915 60.855 ;
        RECT 210.955 60.535 211.215 60.855 ;
        RECT 207.275 59.175 207.535 59.495 ;
        RECT 206.815 58.835 207.075 59.155 ;
        RECT 204.975 58.495 205.235 58.815 ;
        RECT 204.975 57.815 205.235 58.135 ;
        RECT 205.035 56.775 205.175 57.815 ;
        RECT 204.975 56.455 205.235 56.775 ;
        RECT 206.355 56.115 206.615 56.435 ;
        RECT 204.515 53.395 204.775 53.715 ;
        RECT 204.055 53.055 204.315 53.375 ;
        RECT 203.135 51.355 203.395 51.675 ;
        RECT 204.575 50.655 204.715 53.395 ;
        RECT 206.415 53.035 206.555 56.115 ;
        RECT 206.875 55.415 207.015 58.835 ;
        RECT 206.815 55.095 207.075 55.415 ;
        RECT 206.355 52.715 206.615 53.035 ;
        RECT 203.135 50.335 203.395 50.655 ;
        RECT 204.515 50.335 204.775 50.655 ;
        RECT 202.215 49.655 202.475 49.975 ;
        RECT 201.755 48.635 202.015 48.955 ;
        RECT 202.275 48.615 202.415 49.655 ;
        RECT 202.215 48.295 202.475 48.615 ;
        RECT 202.275 47.935 202.415 48.295 ;
        RECT 202.215 47.615 202.475 47.935 ;
        RECT 203.195 47.255 203.335 50.335 ;
        RECT 206.875 50.315 207.015 55.095 ;
        RECT 207.335 51.675 207.475 59.175 ;
        RECT 208.715 58.475 208.855 60.535 ;
        RECT 211.015 59.595 211.155 60.535 ;
        RECT 211.015 59.455 211.615 59.595 ;
        RECT 208.655 58.155 208.915 58.475 ;
        RECT 207.735 55.775 207.995 56.095 ;
        RECT 207.275 51.355 207.535 51.675 ;
        RECT 206.815 49.995 207.075 50.315 ;
        RECT 207.795 48.955 207.935 55.775 ;
        RECT 208.195 51.355 208.455 51.675 ;
        RECT 204.975 48.635 205.235 48.955 ;
        RECT 207.735 48.635 207.995 48.955 ;
        RECT 205.035 47.935 205.175 48.635 ;
        RECT 208.255 47.935 208.395 51.355 ;
        RECT 204.975 47.615 205.235 47.935 ;
        RECT 208.195 47.615 208.455 47.935 ;
        RECT 208.255 47.255 208.395 47.615 ;
        RECT 203.135 46.935 203.395 47.255 ;
        RECT 204.515 46.935 204.775 47.255 ;
        RECT 208.195 46.935 208.455 47.255 ;
        RECT 203.195 46.235 203.335 46.935 ;
        RECT 203.135 45.915 203.395 46.235 ;
        RECT 201.295 44.895 201.555 45.215 ;
        RECT 201.755 43.195 202.015 43.515 ;
        RECT 200.835 41.835 201.095 42.155 ;
        RECT 200.895 40.795 201.035 41.835 ;
        RECT 201.815 40.795 201.955 43.195 ;
        RECT 204.575 42.835 204.715 46.935 ;
        RECT 208.715 45.215 208.855 58.155 ;
        RECT 211.475 57.115 211.615 59.455 ;
        RECT 211.415 56.795 211.675 57.115 ;
        RECT 210.955 56.515 211.215 56.775 ;
        RECT 211.935 56.515 212.075 64.615 ;
        RECT 212.325 64.420 212.605 64.790 ;
        RECT 212.855 61.875 212.995 82.975 ;
        RECT 213.315 80.235 213.455 82.975 ;
        RECT 213.775 81.110 213.915 83.575 ;
        RECT 213.705 80.740 213.985 81.110 ;
        RECT 213.255 79.915 213.515 80.235 ;
        RECT 213.315 64.110 213.455 79.915 ;
        RECT 213.775 78.390 213.915 80.740 ;
        RECT 214.235 79.895 214.375 105.075 ;
        RECT 216.995 104.795 217.135 109.225 ;
        RECT 218.775 107.115 219.035 107.435 ;
        RECT 218.835 106.075 218.975 107.115 ;
        RECT 218.775 105.755 219.035 106.075 ;
        RECT 216.535 104.655 217.135 104.795 ;
        RECT 214.635 101.675 214.895 101.995 ;
        RECT 214.175 79.575 214.435 79.895 ;
        RECT 213.705 78.020 213.985 78.390 ;
        RECT 214.235 78.195 214.375 79.575 ;
        RECT 214.175 77.875 214.435 78.195 ;
        RECT 213.715 77.195 213.975 77.515 ;
        RECT 213.775 76.155 213.915 77.195 ;
        RECT 213.715 75.835 213.975 76.155 ;
        RECT 213.245 63.740 213.525 64.110 ;
        RECT 212.795 61.555 213.055 61.875 ;
        RECT 210.955 56.455 212.075 56.515 ;
        RECT 211.015 56.375 212.075 56.455 ;
        RECT 212.335 56.115 212.595 56.435 ;
        RECT 210.495 55.435 210.755 55.755 ;
        RECT 210.555 53.375 210.695 55.435 ;
        RECT 209.575 53.055 209.835 53.375 ;
        RECT 210.495 53.055 210.755 53.375 ;
        RECT 209.635 50.655 209.775 53.055 ;
        RECT 210.035 52.715 210.295 53.035 ;
        RECT 210.095 50.995 210.235 52.715 ;
        RECT 210.955 52.375 211.215 52.695 ;
        RECT 211.415 52.375 211.675 52.695 ;
        RECT 211.015 50.995 211.155 52.375 ;
        RECT 211.475 51.675 211.615 52.375 ;
        RECT 212.395 51.675 212.535 56.115 ;
        RECT 211.415 51.355 211.675 51.675 ;
        RECT 212.335 51.355 212.595 51.675 ;
        RECT 210.035 50.675 210.295 50.995 ;
        RECT 210.955 50.675 211.215 50.995 ;
        RECT 209.575 50.335 209.835 50.655 ;
        RECT 209.635 47.935 209.775 50.335 ;
        RECT 210.095 50.315 210.235 50.675 ;
        RECT 210.035 49.995 210.295 50.315 ;
        RECT 210.095 48.955 210.235 49.995 ;
        RECT 211.015 48.955 211.155 50.675 ;
        RECT 210.035 48.635 210.295 48.955 ;
        RECT 210.955 48.635 211.215 48.955 ;
        RECT 209.575 47.615 209.835 47.935 ;
        RECT 209.115 45.235 209.375 45.555 ;
        RECT 207.735 44.895 207.995 45.215 ;
        RECT 208.655 44.895 208.915 45.215 ;
        RECT 204.515 42.515 204.775 42.835 ;
        RECT 200.835 40.475 201.095 40.795 ;
        RECT 201.755 40.475 202.015 40.795 ;
        RECT 203.135 39.795 203.395 40.115 ;
        RECT 200.835 39.455 201.095 39.775 ;
        RECT 200.895 38.075 201.035 39.455 ;
        RECT 200.835 37.755 201.095 38.075 ;
        RECT 200.375 36.395 200.635 36.715 ;
        RECT 198.585 35.520 200.125 35.890 ;
        RECT 198.075 34.695 198.335 35.015 ;
        RECT 197.615 32.315 197.875 32.635 ;
        RECT 196.695 30.955 196.955 31.275 ;
        RECT 200.435 30.935 200.575 36.395 ;
        RECT 200.835 34.015 201.095 34.335 ;
        RECT 200.895 32.635 201.035 34.015 ;
        RECT 200.835 32.315 201.095 32.635 ;
        RECT 200.375 30.615 200.635 30.935 ;
        RECT 198.585 30.080 200.125 30.450 ;
        RECT 200.435 29.825 200.575 30.615 ;
        RECT 199.975 29.685 200.575 29.825 ;
        RECT 195.315 28.575 195.575 28.895 ;
        RECT 190.715 26.195 190.975 26.515 ;
        RECT 191.635 26.195 191.895 26.515 ;
        RECT 190.255 25.855 190.515 26.175 ;
        RECT 199.975 25.835 200.115 29.685 ;
        RECT 201.755 29.255 202.015 29.575 ;
        RECT 201.815 27.195 201.955 29.255 ;
        RECT 203.195 28.895 203.335 39.795 ;
        RECT 204.575 39.775 204.715 42.515 ;
        RECT 204.515 39.455 204.775 39.775 ;
        RECT 205.895 38.775 206.155 39.095 ;
        RECT 205.955 37.395 206.095 38.775 ;
        RECT 205.895 37.075 206.155 37.395 ;
        RECT 204.055 35.035 204.315 35.355 ;
        RECT 203.135 28.575 203.395 28.895 ;
        RECT 201.755 26.875 202.015 27.195 ;
        RECT 204.115 26.175 204.255 35.035 ;
        RECT 205.955 30.935 206.095 37.075 ;
        RECT 207.275 36.395 207.535 36.715 ;
        RECT 207.335 35.355 207.475 36.395 ;
        RECT 207.275 35.035 207.535 35.355 ;
        RECT 206.355 34.015 206.615 34.335 ;
        RECT 205.435 30.615 205.695 30.935 ;
        RECT 205.895 30.615 206.155 30.935 ;
        RECT 205.495 29.235 205.635 30.615 ;
        RECT 205.435 28.915 205.695 29.235 ;
        RECT 205.495 27.195 205.635 28.915 ;
        RECT 206.415 28.215 206.555 34.015 ;
        RECT 207.795 32.295 207.935 44.895 ;
        RECT 209.175 42.155 209.315 45.235 ;
        RECT 209.115 41.835 209.375 42.155 ;
        RECT 211.415 41.835 211.675 42.155 ;
        RECT 211.475 40.115 211.615 41.835 ;
        RECT 211.415 39.795 211.675 40.115 ;
        RECT 212.855 38.075 212.995 61.555 ;
        RECT 213.315 55.755 213.455 63.740 ;
        RECT 213.775 59.495 213.915 75.835 ;
        RECT 214.235 75.135 214.375 77.875 ;
        RECT 214.175 74.815 214.435 75.135 ;
        RECT 214.695 72.950 214.835 101.675 ;
        RECT 216.535 100.635 216.675 104.655 ;
        RECT 217.215 103.520 218.755 103.890 ;
        RECT 219.295 102.585 219.435 109.225 ;
        RECT 221.075 106.775 221.335 107.095 ;
        RECT 221.135 106.075 221.275 106.775 ;
        RECT 221.595 106.075 221.735 109.225 ;
        RECT 223.895 107.095 224.035 109.225 ;
        RECT 224.295 107.455 224.555 107.775 ;
        RECT 223.835 106.775 224.095 107.095 ;
        RECT 221.075 105.755 221.335 106.075 ;
        RECT 221.535 105.755 221.795 106.075 ;
        RECT 219.695 104.735 219.955 105.055 ;
        RECT 221.995 104.735 222.255 105.055 ;
        RECT 218.835 102.445 219.435 102.585 ;
        RECT 218.835 100.635 218.975 102.445 ;
        RECT 219.235 101.675 219.495 101.995 ;
        RECT 216.475 100.315 216.735 100.635 ;
        RECT 218.775 100.315 219.035 100.635 ;
        RECT 215.095 99.635 215.355 99.955 ;
        RECT 215.155 95.195 215.295 99.635 ;
        RECT 216.475 99.295 216.735 99.615 ;
        RECT 216.015 98.615 216.275 98.935 ;
        RECT 216.075 96.895 216.215 98.615 ;
        RECT 216.535 97.235 216.675 99.295 ;
        RECT 217.215 98.080 218.755 98.450 ;
        RECT 219.295 97.915 219.435 101.675 ;
        RECT 219.755 100.635 219.895 104.735 ;
        RECT 220.615 104.395 220.875 104.715 ;
        RECT 219.695 100.315 219.955 100.635 ;
        RECT 219.755 97.915 219.895 100.315 ;
        RECT 220.675 99.470 220.815 104.395 ;
        RECT 220.605 99.100 220.885 99.470 ;
        RECT 220.675 98.110 220.815 99.100 ;
        RECT 219.235 97.595 219.495 97.915 ;
        RECT 219.695 97.595 219.955 97.915 ;
        RECT 220.605 97.740 220.885 98.110 ;
        RECT 218.315 97.255 218.575 97.575 ;
        RECT 216.475 96.915 216.735 97.235 ;
        RECT 216.015 96.575 216.275 96.895 ;
        RECT 216.015 95.895 216.275 96.215 ;
        RECT 215.095 94.875 215.355 95.195 ;
        RECT 215.555 93.175 215.815 93.495 ;
        RECT 215.095 90.455 215.355 90.775 ;
        RECT 215.155 85.335 215.295 90.455 ;
        RECT 215.615 89.755 215.755 93.175 ;
        RECT 215.555 89.435 215.815 89.755 ;
        RECT 215.095 85.015 215.355 85.335 ;
        RECT 215.155 76.155 215.295 85.015 ;
        RECT 215.555 81.275 215.815 81.595 ;
        RECT 215.095 75.835 215.355 76.155 ;
        RECT 215.095 74.135 215.355 74.455 ;
        RECT 214.625 72.580 214.905 72.950 ;
        RECT 214.635 66.995 214.895 67.315 ;
        RECT 214.695 65.275 214.835 66.995 ;
        RECT 214.635 64.955 214.895 65.275 ;
        RECT 215.155 61.390 215.295 74.135 ;
        RECT 215.615 62.555 215.755 81.275 ;
        RECT 216.075 80.915 216.215 95.895 ;
        RECT 218.375 94.710 218.515 97.255 ;
        RECT 219.685 97.060 219.965 97.430 ;
        RECT 221.075 97.255 221.335 97.575 ;
        RECT 219.755 96.895 219.895 97.060 ;
        RECT 219.695 96.575 219.955 96.895 ;
        RECT 220.155 96.805 220.415 96.895 ;
        RECT 220.155 96.665 220.815 96.805 ;
        RECT 220.155 96.575 220.415 96.665 ;
        RECT 219.695 95.895 219.955 96.215 ;
        RECT 219.755 95.195 219.895 95.895 ;
        RECT 219.235 94.875 219.495 95.195 ;
        RECT 219.695 94.875 219.955 95.195 ;
        RECT 216.475 94.195 216.735 94.515 ;
        RECT 218.305 94.340 218.585 94.710 ;
        RECT 218.315 94.195 218.575 94.340 ;
        RECT 218.775 94.195 219.035 94.515 ;
        RECT 216.535 92.475 216.675 94.195 ;
        RECT 218.835 93.495 218.975 94.195 ;
        RECT 218.775 93.175 219.035 93.495 ;
        RECT 217.215 92.640 218.755 93.010 ;
        RECT 216.475 92.155 216.735 92.475 ;
        RECT 216.935 90.795 217.195 91.115 ;
        RECT 216.995 88.735 217.135 90.795 ;
        RECT 216.935 88.415 217.195 88.735 ;
        RECT 217.215 87.200 218.755 87.570 ;
        RECT 219.295 86.605 219.435 94.875 ;
        RECT 219.695 94.195 219.955 94.515 ;
        RECT 220.155 94.195 220.415 94.515 ;
        RECT 219.755 91.795 219.895 94.195 ;
        RECT 219.695 91.475 219.955 91.795 ;
        RECT 219.695 90.455 219.955 90.775 ;
        RECT 219.755 89.755 219.895 90.455 ;
        RECT 220.215 89.755 220.355 94.195 ;
        RECT 220.675 92.475 220.815 96.665 ;
        RECT 221.135 95.195 221.275 97.255 ;
        RECT 221.535 95.895 221.795 96.215 ;
        RECT 221.075 94.875 221.335 95.195 ;
        RECT 221.595 94.425 221.735 95.895 ;
        RECT 221.135 94.285 221.735 94.425 ;
        RECT 221.135 93.495 221.275 94.285 ;
        RECT 221.075 93.175 221.335 93.495 ;
        RECT 220.615 92.155 220.875 92.475 ;
        RECT 220.615 91.310 220.875 91.455 ;
        RECT 220.605 90.940 220.885 91.310 ;
        RECT 221.535 91.025 221.795 91.115 ;
        RECT 221.135 90.885 221.795 91.025 ;
        RECT 219.695 89.435 219.955 89.755 ;
        RECT 220.155 89.435 220.415 89.755 ;
        RECT 221.135 89.415 221.275 90.885 ;
        RECT 221.535 90.795 221.795 90.885 ;
        RECT 222.055 89.665 222.195 104.735 ;
        RECT 223.365 99.780 223.645 100.150 ;
        RECT 223.375 99.635 223.635 99.780 ;
        RECT 224.355 96.895 224.495 107.455 ;
        RECT 226.195 106.075 226.335 109.225 ;
        RECT 228.495 106.075 228.635 109.225 ;
        RECT 226.135 105.755 226.395 106.075 ;
        RECT 228.435 105.755 228.695 106.075 ;
        RECT 229.355 105.075 229.615 105.395 ;
        RECT 226.135 103.035 226.395 103.355 ;
        RECT 226.195 100.635 226.335 103.035 ;
        RECT 228.435 101.675 228.695 101.995 ;
        RECT 228.495 100.635 228.635 101.675 ;
        RECT 229.415 101.510 229.555 105.075 ;
        RECT 230.795 104.375 230.935 109.225 ;
        RECT 233.095 106.075 233.235 109.225 ;
        RECT 235.395 106.075 235.535 109.225 ;
        RECT 235.845 106.240 237.385 106.610 ;
        RECT 233.035 105.755 233.295 106.075 ;
        RECT 235.335 105.755 235.595 106.075 ;
        RECT 231.655 105.305 231.915 105.395 ;
        RECT 231.655 105.165 232.315 105.305 ;
        RECT 231.655 105.075 231.915 105.165 ;
        RECT 230.735 104.055 230.995 104.375 ;
        RECT 229.345 101.140 229.625 101.510 ;
        RECT 224.755 100.315 225.015 100.635 ;
        RECT 226.135 100.315 226.395 100.635 ;
        RECT 228.435 100.315 228.695 100.635 ;
        RECT 222.455 96.575 222.715 96.895 ;
        RECT 224.295 96.805 224.555 96.895 ;
        RECT 222.975 96.665 224.555 96.805 ;
        RECT 222.515 96.215 222.655 96.575 ;
        RECT 222.455 95.895 222.715 96.215 ;
        RECT 222.455 94.875 222.715 95.195 ;
        RECT 222.515 94.710 222.655 94.875 ;
        RECT 222.445 94.340 222.725 94.710 ;
        RECT 222.975 94.175 223.115 96.665 ;
        RECT 224.295 96.575 224.555 96.665 ;
        RECT 224.815 95.275 224.955 100.315 ;
        RECT 227.055 99.975 227.315 100.295 ;
        RECT 225.675 99.295 225.935 99.615 ;
        RECT 225.215 97.595 225.475 97.915 ;
        RECT 225.275 96.215 225.415 97.595 ;
        RECT 225.215 95.895 225.475 96.215 ;
        RECT 223.435 95.135 224.955 95.275 ;
        RECT 222.455 93.855 222.715 94.175 ;
        RECT 222.915 93.855 223.175 94.175 ;
        RECT 221.595 89.525 222.195 89.665 ;
        RECT 221.075 89.095 221.335 89.415 ;
        RECT 221.075 88.415 221.335 88.735 ;
        RECT 219.295 86.465 220.815 86.605 ;
        RECT 220.155 85.870 220.415 86.015 ;
        RECT 220.145 85.500 220.425 85.870 ;
        RECT 216.475 82.635 216.735 82.955 ;
        RECT 216.015 80.595 216.275 80.915 ;
        RECT 216.535 80.430 216.675 82.635 ;
        RECT 217.215 81.760 218.755 82.130 ;
        RECT 216.465 80.060 216.745 80.430 ;
        RECT 220.155 80.255 220.415 80.575 ;
        RECT 216.015 78.555 216.275 78.875 ;
        RECT 216.075 74.455 216.215 78.555 ;
        RECT 216.535 75.135 216.675 80.060 ;
        RECT 219.695 78.555 219.955 78.875 ;
        RECT 219.755 78.195 219.895 78.555 ;
        RECT 220.215 78.195 220.355 80.255 ;
        RECT 218.775 77.875 219.035 78.195 ;
        RECT 219.695 77.875 219.955 78.195 ;
        RECT 220.155 77.875 220.415 78.195 ;
        RECT 218.835 77.425 218.975 77.875 ;
        RECT 218.835 77.285 219.435 77.425 ;
        RECT 219.685 77.340 219.965 77.710 ;
        RECT 217.215 76.320 218.755 76.690 ;
        RECT 219.295 76.155 219.435 77.285 ;
        RECT 219.235 75.835 219.495 76.155 ;
        RECT 216.475 74.815 216.735 75.135 ;
        RECT 216.015 74.135 216.275 74.455 ;
        RECT 216.015 70.395 216.275 70.715 ;
        RECT 215.555 62.235 215.815 62.555 ;
        RECT 216.075 61.535 216.215 70.395 ;
        RECT 214.635 60.875 214.895 61.195 ;
        RECT 215.085 61.020 215.365 61.390 ;
        RECT 215.555 61.215 215.815 61.535 ;
        RECT 216.015 61.215 216.275 61.535 ;
        RECT 214.695 59.835 214.835 60.875 ;
        RECT 214.635 59.515 214.895 59.835 ;
        RECT 215.155 59.495 215.295 61.020 ;
        RECT 213.715 59.175 213.975 59.495 ;
        RECT 215.095 59.175 215.355 59.495 ;
        RECT 215.615 58.475 215.755 61.215 ;
        RECT 216.535 58.475 216.675 74.815 ;
        RECT 219.235 74.475 219.495 74.795 ;
        RECT 219.295 73.630 219.435 74.475 ;
        RECT 219.225 73.260 219.505 73.630 ;
        RECT 219.755 73.435 219.895 77.340 ;
        RECT 220.215 77.030 220.355 77.875 ;
        RECT 220.145 76.660 220.425 77.030 ;
        RECT 220.155 75.155 220.415 75.475 ;
        RECT 220.215 74.310 220.355 75.155 ;
        RECT 220.145 73.940 220.425 74.310 ;
        RECT 219.695 73.115 219.955 73.435 ;
        RECT 220.675 73.395 220.815 86.465 ;
        RECT 221.135 82.470 221.275 88.415 ;
        RECT 221.065 82.100 221.345 82.470 ;
        RECT 221.135 78.195 221.275 82.100 ;
        RECT 221.595 78.875 221.735 89.525 ;
        RECT 222.515 87.230 222.655 93.855 ;
        RECT 223.435 89.755 223.575 95.135 ;
        RECT 223.835 94.535 224.095 94.855 ;
        RECT 223.895 93.235 224.035 94.535 ;
        RECT 224.815 94.515 224.955 95.135 ;
        RECT 224.755 94.195 225.015 94.515 ;
        RECT 224.745 93.235 225.025 93.350 ;
        RECT 223.895 93.095 225.025 93.235 ;
        RECT 224.745 92.980 225.025 93.095 ;
        RECT 224.285 90.940 224.565 91.310 ;
        RECT 224.355 90.775 224.495 90.940 ;
        RECT 223.835 90.455 224.095 90.775 ;
        RECT 224.295 90.455 224.555 90.775 ;
        RECT 223.375 89.435 223.635 89.755 ;
        RECT 223.375 88.755 223.635 89.075 ;
        RECT 223.435 88.055 223.575 88.755 ;
        RECT 223.375 87.965 223.635 88.055 ;
        RECT 222.975 87.825 223.635 87.965 ;
        RECT 222.445 86.860 222.725 87.230 ;
        RECT 222.455 86.375 222.715 86.695 ;
        RECT 222.515 84.315 222.655 86.375 ;
        RECT 222.455 83.995 222.715 84.315 ;
        RECT 222.455 82.295 222.715 82.615 ;
        RECT 222.515 80.235 222.655 82.295 ;
        RECT 222.455 80.145 222.715 80.235 ;
        RECT 222.055 80.005 222.715 80.145 ;
        RECT 221.535 78.555 221.795 78.875 ;
        RECT 221.075 77.875 221.335 78.195 ;
        RECT 221.065 73.940 221.345 74.310 ;
        RECT 220.215 73.255 220.815 73.395 ;
        RECT 219.235 71.755 219.495 72.075 ;
        RECT 217.215 70.880 218.755 71.250 ;
        RECT 219.295 66.635 219.435 71.755 ;
        RECT 219.235 66.315 219.495 66.635 ;
        RECT 217.215 65.440 218.755 65.810 ;
        RECT 216.935 64.615 217.195 64.935 ;
        RECT 216.995 61.535 217.135 64.615 ;
        RECT 219.235 63.595 219.495 63.915 ;
        RECT 219.295 62.635 219.435 63.595 ;
        RECT 218.375 62.555 219.435 62.635 ;
        RECT 219.755 62.555 219.895 73.115 ;
        RECT 220.215 66.830 220.355 73.255 ;
        RECT 221.135 67.225 221.275 73.940 ;
        RECT 221.595 72.075 221.735 78.555 ;
        RECT 222.055 75.135 222.195 80.005 ;
        RECT 222.455 79.915 222.715 80.005 ;
        RECT 222.455 78.555 222.715 78.875 ;
        RECT 221.995 74.815 222.255 75.135 ;
        RECT 222.055 73.435 222.195 74.815 ;
        RECT 222.515 74.795 222.655 78.555 ;
        RECT 222.975 78.195 223.115 87.825 ;
        RECT 223.375 87.735 223.635 87.825 ;
        RECT 223.375 85.695 223.635 86.015 ;
        RECT 223.435 83.635 223.575 85.695 ;
        RECT 223.895 83.635 224.035 90.455 ;
        RECT 224.815 88.395 224.955 92.980 ;
        RECT 224.755 88.075 225.015 88.395 ;
        RECT 225.275 87.795 225.415 95.895 ;
        RECT 224.815 87.655 225.415 87.795 ;
        RECT 224.295 85.355 224.555 85.675 ;
        RECT 223.375 83.315 223.635 83.635 ;
        RECT 223.835 83.315 224.095 83.635 ;
        RECT 223.435 80.235 223.575 83.315 ;
        RECT 223.895 80.915 224.035 83.315 ;
        RECT 223.835 80.595 224.095 80.915 ;
        RECT 223.375 79.915 223.635 80.235 ;
        RECT 223.435 78.875 223.575 79.915 ;
        RECT 223.375 78.555 223.635 78.875 ;
        RECT 222.915 77.875 223.175 78.195 ;
        RECT 223.365 78.020 223.645 78.390 ;
        RECT 223.375 77.875 223.635 78.020 ;
        RECT 223.375 77.195 223.635 77.515 ;
        RECT 223.435 75.815 223.575 77.195 ;
        RECT 223.375 75.495 223.635 75.815 ;
        RECT 223.895 75.135 224.035 80.595 ;
        RECT 223.835 74.815 224.095 75.135 ;
        RECT 222.455 74.475 222.715 74.795 ;
        RECT 221.995 73.115 222.255 73.435 ;
        RECT 222.515 73.095 222.655 74.475 ;
        RECT 222.455 72.775 222.715 73.095 ;
        RECT 221.535 71.755 221.795 72.075 ;
        RECT 221.595 70.625 221.735 71.755 ;
        RECT 221.595 70.485 222.195 70.625 ;
        RECT 222.055 70.035 222.195 70.485 ;
        RECT 221.995 69.715 222.255 70.035 ;
        RECT 220.675 67.085 221.275 67.225 ;
        RECT 220.145 66.460 220.425 66.830 ;
        RECT 220.675 66.205 220.815 67.085 ;
        RECT 221.995 66.995 222.255 67.315 ;
        RECT 221.535 66.655 221.795 66.975 ;
        RECT 220.215 66.065 220.815 66.205 ;
        RECT 218.315 62.495 219.435 62.555 ;
        RECT 218.315 62.235 218.575 62.495 ;
        RECT 216.935 61.215 217.195 61.535 ;
        RECT 217.215 60.000 218.755 60.370 ;
        RECT 215.555 58.155 215.815 58.475 ;
        RECT 216.475 58.155 216.735 58.475 ;
        RECT 214.175 56.795 214.435 57.115 ;
        RECT 214.235 55.755 214.375 56.795 ;
        RECT 214.635 56.455 214.895 56.775 ;
        RECT 213.255 55.435 213.515 55.755 ;
        RECT 214.175 55.435 214.435 55.755 ;
        RECT 214.235 54.055 214.375 55.435 ;
        RECT 214.175 53.735 214.435 54.055 ;
        RECT 214.175 52.375 214.435 52.695 ;
        RECT 214.235 50.995 214.375 52.375 ;
        RECT 214.175 50.675 214.435 50.995 ;
        RECT 214.695 48.275 214.835 56.455 ;
        RECT 215.615 55.755 215.755 58.155 ;
        RECT 219.295 56.095 219.435 62.495 ;
        RECT 219.695 62.235 219.955 62.555 ;
        RECT 220.215 61.535 220.355 66.065 ;
        RECT 221.595 65.275 221.735 66.655 ;
        RECT 221.535 64.955 221.795 65.275 ;
        RECT 220.615 63.935 220.875 64.255 ;
        RECT 222.055 64.110 222.195 66.995 ;
        RECT 220.675 61.875 220.815 63.935 ;
        RECT 221.985 63.740 222.265 64.110 ;
        RECT 221.525 63.060 221.805 63.430 ;
        RECT 220.615 61.555 220.875 61.875 ;
        RECT 220.155 61.215 220.415 61.535 ;
        RECT 219.235 55.775 219.495 56.095 ;
        RECT 215.555 55.435 215.815 55.755 ;
        RECT 215.615 51.675 215.755 55.435 ;
        RECT 216.475 55.095 216.735 55.415 ;
        RECT 216.535 53.375 216.675 55.095 ;
        RECT 217.215 54.560 218.755 54.930 ;
        RECT 216.015 53.055 216.275 53.375 ;
        RECT 216.475 53.055 216.735 53.375 ;
        RECT 215.555 51.355 215.815 51.675 ;
        RECT 216.075 50.655 216.215 53.055 ;
        RECT 216.015 50.335 216.275 50.655 ;
        RECT 215.095 49.995 215.355 50.315 ;
        RECT 214.635 47.955 214.895 48.275 ;
        RECT 214.695 46.315 214.835 47.955 ;
        RECT 215.155 47.255 215.295 49.995 ;
        RECT 215.555 48.635 215.815 48.955 ;
        RECT 215.095 46.935 215.355 47.255 ;
        RECT 214.235 46.175 214.835 46.315 ;
        RECT 213.715 43.195 213.975 43.515 ;
        RECT 213.255 42.855 213.515 43.175 ;
        RECT 213.315 40.795 213.455 42.855 ;
        RECT 213.255 40.475 213.515 40.795 ;
        RECT 212.795 37.755 213.055 38.075 ;
        RECT 212.335 36.055 212.595 36.375 ;
        RECT 209.575 35.035 209.835 35.355 ;
        RECT 209.635 34.675 209.775 35.035 ;
        RECT 210.495 34.695 210.755 35.015 ;
        RECT 209.575 34.355 209.835 34.675 ;
        RECT 207.735 31.975 207.995 32.295 ;
        RECT 210.555 29.915 210.695 34.695 ;
        RECT 212.395 31.275 212.535 36.055 ;
        RECT 212.855 35.355 212.995 37.755 ;
        RECT 212.795 35.035 213.055 35.355 ;
        RECT 213.255 34.355 213.515 34.675 ;
        RECT 213.315 33.655 213.455 34.355 ;
        RECT 213.775 34.335 213.915 43.195 ;
        RECT 214.235 42.835 214.375 46.175 ;
        RECT 215.615 45.215 215.755 48.635 ;
        RECT 216.075 46.235 216.215 50.335 ;
        RECT 216.535 48.865 216.675 53.055 ;
        RECT 216.935 52.375 217.195 52.695 ;
        RECT 219.695 52.435 219.955 52.695 ;
        RECT 219.295 52.375 219.955 52.435 ;
        RECT 216.995 50.315 217.135 52.375 ;
        RECT 219.295 52.295 219.895 52.375 ;
        RECT 216.935 49.995 217.195 50.315 ;
        RECT 217.215 49.120 218.755 49.490 ;
        RECT 216.535 48.725 217.135 48.865 ;
        RECT 216.475 46.935 216.735 47.255 ;
        RECT 216.015 45.915 216.275 46.235 ;
        RECT 216.535 45.895 216.675 46.935 ;
        RECT 216.475 45.575 216.735 45.895 ;
        RECT 215.555 44.895 215.815 45.215 ;
        RECT 216.475 44.895 216.735 45.215 ;
        RECT 214.175 42.515 214.435 42.835 ;
        RECT 216.535 42.495 216.675 44.895 ;
        RECT 216.995 44.535 217.135 48.725 ;
        RECT 219.295 47.935 219.435 52.295 ;
        RECT 220.215 51.755 220.355 61.215 ;
        RECT 221.595 60.855 221.735 63.060 ;
        RECT 221.535 60.535 221.795 60.855 ;
        RECT 221.535 57.815 221.795 58.135 ;
        RECT 221.075 56.115 221.335 56.435 ;
        RECT 221.135 53.375 221.275 56.115 ;
        RECT 221.075 53.055 221.335 53.375 ;
        RECT 220.215 51.615 220.815 51.755 ;
        RECT 220.155 50.675 220.415 50.995 ;
        RECT 219.695 50.335 219.955 50.655 ;
        RECT 219.755 48.275 219.895 50.335 ;
        RECT 219.695 47.955 219.955 48.275 ;
        RECT 219.235 47.615 219.495 47.935 ;
        RECT 219.755 45.215 219.895 47.955 ;
        RECT 220.215 47.935 220.355 50.675 ;
        RECT 220.675 50.315 220.815 51.615 ;
        RECT 220.615 49.995 220.875 50.315 ;
        RECT 220.675 48.615 220.815 49.995 ;
        RECT 221.595 49.975 221.735 57.815 ;
        RECT 221.535 49.655 221.795 49.975 ;
        RECT 220.615 48.295 220.875 48.615 ;
        RECT 222.515 47.935 222.655 72.775 ;
        RECT 223.895 71.735 224.035 74.815 ;
        RECT 223.835 71.415 224.095 71.735 ;
        RECT 223.835 70.055 224.095 70.375 ;
        RECT 223.895 68.075 224.035 70.055 ;
        RECT 224.355 69.695 224.495 85.355 ;
        RECT 224.815 80.575 224.955 87.655 ;
        RECT 225.215 82.635 225.475 82.955 ;
        RECT 224.755 80.255 225.015 80.575 ;
        RECT 225.275 78.535 225.415 82.635 ;
        RECT 225.215 78.215 225.475 78.535 ;
        RECT 225.735 77.765 225.875 99.295 ;
        RECT 227.115 96.895 227.255 99.975 ;
        RECT 227.975 99.635 228.235 99.955 ;
        RECT 231.655 99.635 231.915 99.955 ;
        RECT 227.055 96.575 227.315 96.895 ;
        RECT 228.035 96.555 228.175 99.635 ;
        RECT 231.715 98.935 231.855 99.635 ;
        RECT 231.655 98.615 231.915 98.935 ;
        RECT 228.425 97.060 228.705 97.430 ;
        RECT 228.495 96.555 228.635 97.060 ;
        RECT 229.355 96.915 229.615 97.235 ;
        RECT 227.975 96.235 228.235 96.555 ;
        RECT 228.435 96.235 228.695 96.555 ;
        RECT 228.035 95.195 228.175 96.235 ;
        RECT 227.975 94.875 228.235 95.195 ;
        RECT 228.895 93.175 229.155 93.495 ;
        RECT 226.595 92.155 226.855 92.475 ;
        RECT 227.975 92.155 228.235 92.475 ;
        RECT 226.655 90.775 226.795 92.155 ;
        RECT 227.055 91.135 227.315 91.455 ;
        RECT 226.595 90.455 226.855 90.775 ;
        RECT 226.135 88.985 226.395 89.075 ;
        RECT 226.135 88.845 226.795 88.985 ;
        RECT 226.135 88.755 226.395 88.845 ;
        RECT 226.135 87.735 226.395 88.055 ;
        RECT 225.275 77.625 225.875 77.765 ;
        RECT 224.755 77.195 225.015 77.515 ;
        RECT 224.815 75.475 224.955 77.195 ;
        RECT 224.755 75.155 225.015 75.475 ;
        RECT 224.755 71.755 225.015 72.075 ;
        RECT 224.295 69.375 224.555 69.695 ;
        RECT 222.975 67.935 224.035 68.075 ;
        RECT 222.975 66.975 223.115 67.935 ;
        RECT 224.815 67.905 224.955 71.755 ;
        RECT 225.275 67.995 225.415 77.625 ;
        RECT 225.665 73.260 225.945 73.630 ;
        RECT 224.355 67.765 224.955 67.905 ;
        RECT 223.375 67.565 223.635 67.655 ;
        RECT 224.355 67.565 224.495 67.765 ;
        RECT 225.215 67.675 225.475 67.995 ;
        RECT 223.375 67.425 224.495 67.565 ;
        RECT 223.375 67.335 223.635 67.425 ;
        RECT 222.915 66.655 223.175 66.975 ;
        RECT 223.835 66.315 224.095 66.635 ;
        RECT 222.915 64.955 223.175 65.275 ;
        RECT 222.975 63.575 223.115 64.955 ;
        RECT 223.895 64.595 224.035 66.315 ;
        RECT 223.835 64.275 224.095 64.595 ;
        RECT 224.355 64.255 224.495 67.425 ;
        RECT 225.735 67.315 225.875 73.260 ;
        RECT 226.195 67.995 226.335 87.735 ;
        RECT 226.655 87.035 226.795 88.845 ;
        RECT 227.115 88.395 227.255 91.135 ;
        RECT 228.035 89.075 228.175 92.155 ;
        RECT 227.975 88.755 228.235 89.075 ;
        RECT 227.055 88.075 227.315 88.395 ;
        RECT 226.595 86.715 226.855 87.035 ;
        RECT 227.115 83.975 227.255 88.075 ;
        RECT 227.515 86.265 227.775 86.355 ;
        RECT 228.035 86.265 228.175 88.755 ;
        RECT 227.515 86.125 228.175 86.265 ;
        RECT 227.515 86.035 227.775 86.125 ;
        RECT 226.585 83.460 226.865 83.830 ;
        RECT 227.055 83.655 227.315 83.975 ;
        RECT 226.655 70.375 226.795 83.460 ;
        RECT 227.055 82.975 227.315 83.295 ;
        RECT 227.115 82.470 227.255 82.975 ;
        RECT 227.575 82.615 227.715 86.035 ;
        RECT 228.435 85.870 228.695 86.015 ;
        RECT 228.425 85.500 228.705 85.870 ;
        RECT 227.045 82.100 227.325 82.470 ;
        RECT 227.515 82.295 227.775 82.615 ;
        RECT 227.515 80.255 227.775 80.575 ;
        RECT 227.055 79.575 227.315 79.895 ;
        RECT 227.115 76.155 227.255 79.575 ;
        RECT 227.575 76.155 227.715 80.255 ;
        RECT 228.435 79.575 228.695 79.895 ;
        RECT 227.975 77.875 228.235 78.195 ;
        RECT 227.055 75.835 227.315 76.155 ;
        RECT 227.515 75.835 227.775 76.155 ;
        RECT 228.035 75.135 228.175 77.875 ;
        RECT 227.975 74.815 228.235 75.135 ;
        RECT 227.505 74.195 227.785 74.310 ;
        RECT 228.035 74.195 228.175 74.815 ;
        RECT 227.505 74.055 228.175 74.195 ;
        RECT 227.505 73.940 227.785 74.055 ;
        RECT 227.055 72.775 227.315 73.095 ;
        RECT 226.595 70.055 226.855 70.375 ;
        RECT 226.595 69.375 226.855 69.695 ;
        RECT 226.135 67.675 226.395 67.995 ;
        RECT 224.755 66.995 225.015 67.315 ;
        RECT 225.675 67.225 225.935 67.315 ;
        RECT 226.125 67.225 226.405 67.510 ;
        RECT 225.675 67.140 226.405 67.225 ;
        RECT 225.675 67.085 226.335 67.140 ;
        RECT 225.675 66.995 225.935 67.085 ;
        RECT 224.815 65.275 224.955 66.995 ;
        RECT 226.655 66.150 226.795 69.375 ;
        RECT 226.585 65.780 226.865 66.150 ;
        RECT 224.755 64.955 225.015 65.275 ;
        RECT 224.295 63.935 224.555 64.255 ;
        RECT 222.915 63.255 223.175 63.575 ;
        RECT 223.835 63.255 224.095 63.575 ;
        RECT 223.895 62.555 224.035 63.255 ;
        RECT 223.835 62.235 224.095 62.555 ;
        RECT 226.595 60.875 226.855 61.195 ;
        RECT 226.655 59.595 226.795 60.875 ;
        RECT 226.195 59.455 226.795 59.595 ;
        RECT 226.195 58.815 226.335 59.455 ;
        RECT 226.135 58.495 226.395 58.815 ;
        RECT 224.755 57.815 225.015 58.135 ;
        RECT 223.835 56.115 224.095 56.435 ;
        RECT 223.895 48.955 224.035 56.115 ;
        RECT 224.815 55.270 224.955 57.815 ;
        RECT 225.675 56.115 225.935 56.435 ;
        RECT 224.745 54.900 225.025 55.270 ;
        RECT 224.815 54.395 224.955 54.900 ;
        RECT 225.735 54.395 225.875 56.115 ;
        RECT 224.755 54.075 225.015 54.395 ;
        RECT 225.675 54.075 225.935 54.395 ;
        RECT 226.595 52.375 226.855 52.695 ;
        RECT 226.655 51.335 226.795 52.375 ;
        RECT 226.595 51.015 226.855 51.335 ;
        RECT 223.835 48.635 224.095 48.955 ;
        RECT 227.115 47.935 227.255 72.775 ;
        RECT 228.495 69.550 228.635 79.575 ;
        RECT 228.425 69.180 228.705 69.550 ;
        RECT 228.495 67.315 228.635 69.180 ;
        RECT 228.435 66.995 228.695 67.315 ;
        RECT 228.435 66.315 228.695 66.635 ;
        RECT 228.495 59.235 228.635 66.315 ;
        RECT 228.955 61.445 229.095 93.175 ;
        RECT 229.415 80.575 229.555 96.915 ;
        RECT 231.195 96.575 231.455 96.895 ;
        RECT 229.815 95.895 230.075 96.215 ;
        RECT 229.875 94.855 230.015 95.895 ;
        RECT 229.815 94.535 230.075 94.855 ;
        RECT 229.815 91.815 230.075 92.135 ;
        RECT 229.875 88.395 230.015 91.815 ;
        RECT 230.275 88.415 230.535 88.735 ;
        RECT 229.815 88.075 230.075 88.395 ;
        RECT 229.815 86.375 230.075 86.695 ;
        RECT 229.875 83.035 230.015 86.375 ;
        RECT 230.335 83.635 230.475 88.415 ;
        RECT 230.735 85.355 230.995 85.675 ;
        RECT 230.275 83.315 230.535 83.635 ;
        RECT 229.875 82.895 230.475 83.035 ;
        RECT 230.795 82.955 230.935 85.355 ;
        RECT 229.355 80.255 229.615 80.575 ;
        RECT 229.415 77.595 229.555 80.255 ;
        RECT 229.805 80.060 230.085 80.430 ;
        RECT 229.875 78.195 230.015 80.060 ;
        RECT 229.815 77.875 230.075 78.195 ;
        RECT 229.415 77.455 230.015 77.595 ;
        RECT 229.355 74.135 229.615 74.455 ;
        RECT 229.415 67.315 229.555 74.135 ;
        RECT 229.875 72.755 230.015 77.455 ;
        RECT 230.335 73.095 230.475 82.895 ;
        RECT 230.735 82.635 230.995 82.955 ;
        RECT 230.735 80.935 230.995 81.255 ;
        RECT 230.275 72.775 230.535 73.095 ;
        RECT 229.815 72.435 230.075 72.755 ;
        RECT 230.795 69.695 230.935 80.935 ;
        RECT 230.735 69.375 230.995 69.695 ;
        RECT 229.815 68.695 230.075 69.015 ;
        RECT 230.275 68.695 230.535 69.015 ;
        RECT 229.875 67.995 230.015 68.695 ;
        RECT 229.815 67.675 230.075 67.995 ;
        RECT 229.355 66.995 229.615 67.315 ;
        RECT 230.335 66.295 230.475 68.695 ;
        RECT 230.275 65.975 230.535 66.295 ;
        RECT 230.275 64.615 230.535 64.935 ;
        RECT 229.355 61.445 229.615 61.535 ;
        RECT 228.955 61.305 229.615 61.445 ;
        RECT 229.355 61.215 229.615 61.305 ;
        RECT 227.575 59.095 228.635 59.235 ;
        RECT 230.335 59.155 230.475 64.615 ;
        RECT 230.795 64.255 230.935 69.375 ;
        RECT 231.255 65.275 231.395 96.575 ;
        RECT 231.715 95.390 231.855 98.615 ;
        RECT 231.645 95.020 231.925 95.390 ;
        RECT 232.175 94.765 232.315 105.165 ;
        RECT 233.035 105.075 233.295 105.395 ;
        RECT 235.795 105.075 236.055 105.395 ;
        RECT 236.255 105.075 236.515 105.395 ;
        RECT 232.575 104.055 232.835 104.375 ;
        RECT 232.635 99.615 232.775 104.055 ;
        RECT 232.575 99.295 232.835 99.615 ;
        RECT 231.715 94.625 232.315 94.765 ;
        RECT 231.715 80.575 231.855 94.625 ;
        RECT 232.575 94.195 232.835 94.515 ;
        RECT 232.115 90.795 232.375 91.115 ;
        RECT 232.175 88.395 232.315 90.795 ;
        RECT 232.115 88.075 232.375 88.395 ;
        RECT 232.635 84.315 232.775 94.195 ;
        RECT 233.095 86.695 233.235 105.075 ;
        RECT 235.855 102.675 235.995 105.075 ;
        RECT 236.315 103.355 236.455 105.075 ;
        RECT 236.715 104.735 236.975 105.055 ;
        RECT 236.775 103.355 236.915 104.735 ;
        RECT 237.695 104.715 237.835 109.225 ;
        RECT 239.995 106.075 240.135 109.225 ;
        RECT 241.775 106.775 242.035 107.095 ;
        RECT 239.935 105.755 240.195 106.075 ;
        RECT 241.315 105.075 241.575 105.395 ;
        RECT 237.635 104.395 237.895 104.715 ;
        RECT 240.395 104.055 240.655 104.375 ;
        RECT 236.255 103.035 236.515 103.355 ;
        RECT 236.715 103.035 236.975 103.355 ;
        RECT 235.795 102.355 236.055 102.675 ;
        RECT 237.635 102.190 237.895 102.335 ;
        RECT 237.625 101.820 237.905 102.190 ;
        RECT 239.935 101.675 240.195 101.995 ;
        RECT 237.635 101.335 237.895 101.655 ;
        RECT 235.845 100.800 237.385 101.170 ;
        RECT 236.715 100.315 236.975 100.635 ;
        RECT 235.795 99.295 236.055 99.615 ;
        RECT 234.875 98.955 235.135 99.275 ;
        RECT 235.335 98.955 235.595 99.275 ;
        RECT 234.405 97.060 234.685 97.430 ;
        RECT 234.415 96.915 234.675 97.060 ;
        RECT 234.935 96.895 235.075 98.955 ;
        RECT 234.875 96.575 235.135 96.895 ;
        RECT 234.415 96.235 234.675 96.555 ;
        RECT 234.475 91.455 234.615 96.235 ;
        RECT 234.935 94.855 235.075 96.575 ;
        RECT 235.395 95.105 235.535 98.955 ;
        RECT 235.855 96.895 235.995 99.295 ;
        RECT 236.775 97.575 236.915 100.315 ;
        RECT 237.695 99.955 237.835 101.335 ;
        RECT 239.465 100.460 239.745 100.830 ;
        RECT 239.995 100.635 240.135 101.675 ;
        RECT 237.635 99.635 237.895 99.955 ;
        RECT 236.715 97.255 236.975 97.575 ;
        RECT 237.165 97.060 237.445 97.430 ;
        RECT 237.235 96.895 237.375 97.060 ;
        RECT 235.795 96.575 236.055 96.895 ;
        RECT 237.175 96.575 237.435 96.895 ;
        RECT 235.845 95.360 237.385 95.730 ;
        RECT 235.395 94.965 235.995 95.105 ;
        RECT 234.875 94.535 235.135 94.855 ;
        RECT 235.325 94.340 235.605 94.710 ;
        RECT 235.855 94.515 235.995 94.965 ;
        RECT 237.695 94.515 237.835 99.635 ;
        RECT 239.535 97.915 239.675 100.460 ;
        RECT 239.935 100.315 240.195 100.635 ;
        RECT 240.455 99.955 240.595 104.055 ;
        RECT 240.395 99.635 240.655 99.955 ;
        RECT 241.375 98.790 241.515 105.075 ;
        RECT 241.835 99.955 241.975 106.775 ;
        RECT 242.295 106.075 242.435 109.225 ;
        RECT 242.235 105.755 242.495 106.075 ;
        RECT 244.595 105.735 244.735 109.225 ;
        RECT 246.375 108.135 246.635 108.455 ;
        RECT 244.535 105.415 244.795 105.735 ;
        RECT 246.435 105.395 246.575 108.135 ;
        RECT 246.375 105.075 246.635 105.395 ;
        RECT 244.995 104.735 245.255 105.055 ;
        RECT 244.075 104.395 244.335 104.715 ;
        RECT 244.135 100.635 244.275 104.395 ;
        RECT 245.055 101.655 245.195 104.735 ;
        RECT 244.995 101.335 245.255 101.655 ;
        RECT 244.075 100.315 244.335 100.635 ;
        RECT 241.775 99.635 242.035 99.955 ;
        RECT 241.305 98.420 241.585 98.790 ;
        RECT 239.475 97.595 239.735 97.915 ;
        RECT 238.555 96.805 238.815 96.895 ;
        RECT 238.155 96.750 238.815 96.805 ;
        RECT 238.085 96.665 238.815 96.750 ;
        RECT 238.085 96.380 238.365 96.665 ;
        RECT 238.555 96.575 238.815 96.665 ;
        RECT 239.935 96.805 240.195 96.895 ;
        RECT 239.935 96.665 240.595 96.805 ;
        RECT 241.375 96.750 241.515 98.420 ;
        RECT 239.935 96.575 240.195 96.665 ;
        RECT 238.615 95.195 238.755 96.575 ;
        RECT 238.555 94.875 238.815 95.195 ;
        RECT 235.395 94.175 235.535 94.340 ;
        RECT 235.795 94.195 236.055 94.515 ;
        RECT 237.635 94.195 237.895 94.515 ;
        RECT 238.085 94.340 238.365 94.710 ;
        RECT 238.095 94.195 238.355 94.340 ;
        RECT 239.475 94.195 239.735 94.515 ;
        RECT 239.935 94.195 240.195 94.515 ;
        RECT 235.335 93.855 235.595 94.175 ;
        RECT 234.415 91.135 234.675 91.455 ;
        RECT 234.875 91.135 235.135 91.455 ;
        RECT 233.955 88.415 234.215 88.735 ;
        RECT 234.015 86.695 234.155 88.415 ;
        RECT 233.035 86.375 233.295 86.695 ;
        RECT 233.955 86.375 234.215 86.695 ;
        RECT 233.495 85.015 233.755 85.335 ;
        RECT 232.575 83.995 232.835 84.315 ;
        RECT 233.035 83.315 233.295 83.635 ;
        RECT 231.655 80.255 231.915 80.575 ;
        RECT 231.715 78.535 231.855 80.255 ;
        RECT 231.655 78.215 231.915 78.535 ;
        RECT 231.715 75.670 231.855 78.215 ;
        RECT 232.575 77.875 232.835 78.195 ;
        RECT 232.115 77.195 232.375 77.515 ;
        RECT 231.645 75.300 231.925 75.670 ;
        RECT 232.175 73.435 232.315 77.195 ;
        RECT 232.635 75.135 232.775 77.875 ;
        RECT 232.575 74.815 232.835 75.135 ;
        RECT 232.115 73.115 232.375 73.435 ;
        RECT 232.105 71.900 232.385 72.270 ;
        RECT 232.175 70.910 232.315 71.900 ;
        RECT 232.105 70.540 232.385 70.910 ;
        RECT 232.115 69.375 232.375 69.695 ;
        RECT 231.195 64.955 231.455 65.275 ;
        RECT 230.735 63.935 230.995 64.255 ;
        RECT 231.255 64.110 231.395 64.955 ;
        RECT 231.185 63.740 231.465 64.110 ;
        RECT 232.175 63.575 232.315 69.375 ;
        RECT 232.635 69.355 232.775 74.815 ;
        RECT 232.575 69.035 232.835 69.355 ;
        RECT 232.115 63.255 232.375 63.575 ;
        RECT 231.655 61.555 231.915 61.875 ;
        RECT 231.715 59.835 231.855 61.555 ;
        RECT 231.655 59.515 231.915 59.835 ;
        RECT 227.575 58.815 227.715 59.095 ;
        RECT 227.515 58.495 227.775 58.815 ;
        RECT 228.495 57.115 228.635 59.095 ;
        RECT 230.275 58.835 230.535 59.155 ;
        RECT 231.185 58.980 231.465 59.350 ;
        RECT 231.255 58.815 231.395 58.980 ;
        RECT 231.655 58.835 231.915 59.155 ;
        RECT 229.355 58.495 229.615 58.815 ;
        RECT 231.195 58.495 231.455 58.815 ;
        RECT 228.895 57.815 229.155 58.135 ;
        RECT 228.435 56.795 228.695 57.115 ;
        RECT 228.955 56.095 229.095 57.815 ;
        RECT 229.415 56.095 229.555 58.495 ;
        RECT 230.275 57.815 230.535 58.135 ;
        RECT 230.335 56.630 230.475 57.815 ;
        RECT 230.265 56.260 230.545 56.630 ;
        RECT 228.895 55.775 229.155 56.095 ;
        RECT 229.355 55.775 229.615 56.095 ;
        RECT 229.355 55.095 229.615 55.415 ;
        RECT 229.415 54.395 229.555 55.095 ;
        RECT 229.355 54.075 229.615 54.395 ;
        RECT 227.515 51.015 227.775 51.335 ;
        RECT 220.155 47.615 220.415 47.935 ;
        RECT 222.455 47.615 222.715 47.935 ;
        RECT 227.055 47.615 227.315 47.935 ;
        RECT 224.755 46.935 225.015 47.255 ;
        RECT 226.135 46.935 226.395 47.255 ;
        RECT 224.815 45.215 224.955 46.935 ;
        RECT 226.195 45.215 226.335 46.935 ;
        RECT 226.595 45.235 226.855 45.555 ;
        RECT 219.695 44.895 219.955 45.215 ;
        RECT 224.755 44.895 225.015 45.215 ;
        RECT 226.135 44.895 226.395 45.215 ;
        RECT 216.935 44.215 217.195 44.535 ;
        RECT 224.295 44.215 224.555 44.535 ;
        RECT 217.215 43.680 218.755 44.050 ;
        RECT 216.475 42.175 216.735 42.495 ;
        RECT 214.175 39.795 214.435 40.115 ;
        RECT 214.235 36.715 214.375 39.795 ;
        RECT 214.175 36.395 214.435 36.715 ;
        RECT 213.715 34.015 213.975 34.335 ;
        RECT 213.255 33.335 213.515 33.655 ;
        RECT 216.015 33.335 216.275 33.655 ;
        RECT 212.335 30.955 212.595 31.275 ;
        RECT 210.495 29.595 210.755 29.915 ;
        RECT 213.315 29.575 213.455 33.335 ;
        RECT 216.075 31.615 216.215 33.335 ;
        RECT 216.535 31.955 216.675 42.175 ;
        RECT 218.775 41.835 219.035 42.155 ;
        RECT 218.835 40.795 218.975 41.835 ;
        RECT 224.355 40.795 224.495 44.215 ;
        RECT 225.215 43.195 225.475 43.515 ;
        RECT 225.275 40.795 225.415 43.195 ;
        RECT 226.655 42.835 226.795 45.235 ;
        RECT 226.595 42.515 226.855 42.835 ;
        RECT 227.115 42.495 227.255 47.615 ;
        RECT 227.055 42.175 227.315 42.495 ;
        RECT 218.775 40.475 219.035 40.795 ;
        RECT 224.295 40.475 224.555 40.795 ;
        RECT 225.215 40.475 225.475 40.795 ;
        RECT 224.755 39.455 225.015 39.775 ;
        RECT 217.215 38.240 218.755 38.610 ;
        RECT 224.815 38.075 224.955 39.455 ;
        RECT 224.755 37.755 225.015 38.075 ;
        RECT 221.535 36.735 221.795 37.055 ;
        RECT 222.915 36.735 223.175 37.055 ;
        RECT 220.155 36.395 220.415 36.715 ;
        RECT 217.215 32.800 218.755 33.170 ;
        RECT 216.475 31.635 216.735 31.955 ;
        RECT 215.555 31.295 215.815 31.615 ;
        RECT 216.015 31.295 216.275 31.615 ;
        RECT 214.175 30.615 214.435 30.935 ;
        RECT 213.255 29.255 213.515 29.575 ;
        RECT 214.235 29.235 214.375 30.615 ;
        RECT 215.095 29.825 215.355 29.915 ;
        RECT 215.615 29.825 215.755 31.295 ;
        RECT 216.015 30.615 216.275 30.935 ;
        RECT 216.075 29.915 216.215 30.615 ;
        RECT 215.095 29.685 215.755 29.825 ;
        RECT 215.095 29.595 215.355 29.685 ;
        RECT 216.015 29.595 216.275 29.915 ;
        RECT 214.175 28.915 214.435 29.235 ;
        RECT 220.215 29.145 220.355 36.395 ;
        RECT 220.615 36.055 220.875 36.375 ;
        RECT 221.075 36.055 221.335 36.375 ;
        RECT 220.675 32.635 220.815 36.055 ;
        RECT 221.135 35.355 221.275 36.055 ;
        RECT 221.595 35.355 221.735 36.735 ;
        RECT 221.075 35.035 221.335 35.355 ;
        RECT 221.535 35.035 221.795 35.355 ;
        RECT 222.975 35.015 223.115 36.735 ;
        RECT 224.815 35.355 224.955 37.755 ;
        RECT 225.675 37.075 225.935 37.395 ;
        RECT 225.735 35.355 225.875 37.075 ;
        RECT 224.755 35.035 225.015 35.355 ;
        RECT 225.675 35.035 225.935 35.355 ;
        RECT 227.575 35.015 227.715 51.015 ;
        RECT 227.975 49.655 228.235 49.975 ;
        RECT 228.035 47.255 228.175 49.655 ;
        RECT 230.275 48.635 230.535 48.955 ;
        RECT 228.435 47.275 228.695 47.595 ;
        RECT 227.975 46.935 228.235 47.255 ;
        RECT 227.975 41.495 228.235 41.815 ;
        RECT 228.035 39.095 228.175 41.495 ;
        RECT 228.495 39.095 228.635 47.275 ;
        RECT 230.335 40.795 230.475 48.635 ;
        RECT 230.735 45.235 230.995 45.555 ;
        RECT 230.795 43.515 230.935 45.235 ;
        RECT 231.715 45.215 231.855 58.835 ;
        RECT 232.175 58.815 232.315 63.255 ;
        RECT 232.575 61.555 232.835 61.875 ;
        RECT 232.115 58.495 232.375 58.815 ;
        RECT 232.635 58.475 232.775 61.555 ;
        RECT 232.575 58.155 232.835 58.475 ;
        RECT 233.095 45.555 233.235 83.315 ;
        RECT 233.555 81.790 233.695 85.015 ;
        RECT 234.015 83.635 234.155 86.375 ;
        RECT 234.935 85.925 235.075 91.135 ;
        RECT 235.395 89.665 235.535 93.855 ;
        RECT 235.845 89.920 237.385 90.290 ;
        RECT 235.395 89.525 237.375 89.665 ;
        RECT 237.235 89.075 237.375 89.525 ;
        RECT 236.715 88.755 236.975 89.075 ;
        RECT 237.175 88.755 237.435 89.075 ;
        RECT 236.775 87.035 236.915 88.755 ;
        RECT 237.175 88.075 237.435 88.395 ;
        RECT 236.715 86.715 236.975 87.035 ;
        RECT 237.235 86.265 237.375 88.075 ;
        RECT 237.695 87.910 237.835 94.195 ;
        RECT 238.155 93.835 238.295 94.195 ;
        RECT 238.095 93.515 238.355 93.835 ;
        RECT 237.625 87.540 237.905 87.910 ;
        RECT 237.635 86.265 237.895 86.355 ;
        RECT 237.235 86.125 237.895 86.265 ;
        RECT 237.635 86.035 237.895 86.125 ;
        RECT 235.335 85.925 235.595 86.015 ;
        RECT 234.935 85.785 235.595 85.925 ;
        RECT 235.335 85.695 235.595 85.785 ;
        RECT 234.875 83.995 235.135 84.315 ;
        RECT 233.955 83.315 234.215 83.635 ;
        RECT 234.415 82.975 234.675 83.295 ;
        RECT 233.955 82.295 234.215 82.615 ;
        RECT 233.485 81.420 233.765 81.790 ;
        RECT 233.555 81.255 233.695 81.420 ;
        RECT 233.495 80.935 233.755 81.255 ;
        RECT 234.015 78.275 234.155 82.295 ;
        RECT 233.555 78.135 234.155 78.275 ;
        RECT 233.555 74.795 233.695 78.135 ;
        RECT 233.955 77.535 234.215 77.855 ;
        RECT 234.015 77.030 234.155 77.535 ;
        RECT 233.945 76.660 234.225 77.030 ;
        RECT 233.955 75.155 234.215 75.475 ;
        RECT 233.495 74.475 233.755 74.795 ;
        RECT 233.495 72.435 233.755 72.755 ;
        RECT 233.555 66.975 233.695 72.435 ;
        RECT 234.015 69.695 234.155 75.155 ;
        RECT 233.955 69.375 234.215 69.695 ;
        RECT 233.495 66.655 233.755 66.975 ;
        RECT 233.955 61.895 234.215 62.215 ;
        RECT 234.015 61.195 234.155 61.895 ;
        RECT 233.495 60.875 233.755 61.195 ;
        RECT 233.955 60.875 234.215 61.195 ;
        RECT 233.555 60.595 233.695 60.875 ;
        RECT 234.475 60.595 234.615 82.975 ;
        RECT 234.935 78.875 235.075 83.995 ;
        RECT 234.875 78.555 235.135 78.875 ;
        RECT 234.875 77.875 235.135 78.195 ;
        RECT 234.935 72.950 235.075 77.875 ;
        RECT 235.395 77.855 235.535 85.695 ;
        RECT 235.845 84.480 237.385 84.850 ;
        RECT 236.715 82.635 236.975 82.955 ;
        RECT 236.775 81.255 236.915 82.635 ;
        RECT 237.175 82.295 237.435 82.615 ;
        RECT 237.235 81.595 237.375 82.295 ;
        RECT 237.175 81.275 237.435 81.595 ;
        RECT 236.715 80.935 236.975 81.255 ;
        RECT 235.845 79.040 237.385 79.410 ;
        RECT 237.175 78.215 237.435 78.535 ;
        RECT 235.335 77.535 235.595 77.855 ;
        RECT 236.715 77.535 236.975 77.855 ;
        RECT 236.255 76.855 236.515 77.175 ;
        RECT 236.315 76.350 236.455 76.855 ;
        RECT 236.245 75.980 236.525 76.350 ;
        RECT 235.335 75.495 235.595 75.815 ;
        RECT 235.395 73.345 235.535 75.495 ;
        RECT 236.775 74.455 236.915 77.535 ;
        RECT 237.235 76.915 237.375 78.215 ;
        RECT 237.695 77.425 237.835 86.035 ;
        RECT 238.155 85.335 238.295 93.515 ;
        RECT 239.015 93.175 239.275 93.495 ;
        RECT 239.075 92.135 239.215 93.175 ;
        RECT 239.015 91.815 239.275 92.135 ;
        RECT 239.535 91.875 239.675 94.195 ;
        RECT 239.995 92.475 240.135 94.195 ;
        RECT 239.935 92.155 240.195 92.475 ;
        RECT 240.455 92.135 240.595 96.665 ;
        RECT 241.305 96.380 241.585 96.750 ;
        RECT 241.315 95.895 241.575 96.215 ;
        RECT 240.855 93.515 241.115 93.835 ;
        RECT 239.535 91.735 240.135 91.875 ;
        RECT 240.395 91.815 240.655 92.135 ;
        RECT 238.555 90.795 238.815 91.115 ;
        RECT 238.615 87.230 238.755 90.795 ;
        RECT 239.475 90.455 239.735 90.775 ;
        RECT 239.535 88.395 239.675 90.455 ;
        RECT 239.475 88.075 239.735 88.395 ;
        RECT 239.465 87.540 239.745 87.910 ;
        RECT 238.545 86.860 238.825 87.230 ;
        RECT 238.095 85.015 238.355 85.335 ;
        RECT 238.615 77.855 238.755 86.860 ;
        RECT 239.535 86.695 239.675 87.540 ;
        RECT 239.475 86.375 239.735 86.695 ;
        RECT 239.475 85.355 239.735 85.675 ;
        RECT 239.535 84.315 239.675 85.355 ;
        RECT 239.475 83.995 239.735 84.315 ;
        RECT 239.015 83.655 239.275 83.975 ;
        RECT 239.075 81.595 239.215 83.655 ;
        RECT 239.015 81.275 239.275 81.595 ;
        RECT 239.995 81.255 240.135 91.735 ;
        RECT 240.395 88.755 240.655 89.075 ;
        RECT 240.455 86.605 240.595 88.755 ;
        RECT 240.915 88.645 241.055 93.515 ;
        RECT 241.375 88.985 241.515 95.895 ;
        RECT 241.835 94.855 241.975 99.635 ;
        RECT 244.535 98.615 244.795 98.935 ;
        RECT 242.235 96.235 242.495 96.555 ;
        RECT 241.775 94.535 242.035 94.855 ;
        RECT 242.295 94.515 242.435 96.235 ;
        RECT 242.695 95.105 242.955 95.195 ;
        RECT 243.615 95.105 243.875 95.195 ;
        RECT 242.695 94.965 243.875 95.105 ;
        RECT 244.065 95.020 244.345 95.390 ;
        RECT 242.695 94.875 242.955 94.965 ;
        RECT 243.615 94.875 243.875 94.965 ;
        RECT 244.135 94.515 244.275 95.020 ;
        RECT 242.235 94.195 242.495 94.515 ;
        RECT 243.615 94.195 243.875 94.515 ;
        RECT 244.075 94.195 244.335 94.515 ;
        RECT 241.775 93.515 242.035 93.835 ;
        RECT 241.835 92.475 241.975 93.515 ;
        RECT 242.295 93.350 242.435 94.195 ;
        RECT 243.675 93.915 243.815 94.195 ;
        RECT 243.215 93.775 243.815 93.915 ;
        RECT 242.225 93.235 242.505 93.350 ;
        RECT 242.225 93.095 242.895 93.235 ;
        RECT 242.225 92.980 242.505 93.095 ;
        RECT 241.775 92.155 242.035 92.475 ;
        RECT 242.225 91.620 242.505 91.990 ;
        RECT 242.295 89.415 242.435 91.620 ;
        RECT 242.755 91.455 242.895 93.095 ;
        RECT 243.215 91.795 243.355 93.775 ;
        RECT 243.155 91.475 243.415 91.795 ;
        RECT 242.695 91.135 242.955 91.455 ;
        RECT 242.695 89.435 242.955 89.755 ;
        RECT 242.235 89.095 242.495 89.415 ;
        RECT 241.375 88.845 241.975 88.985 ;
        RECT 240.915 88.505 241.515 88.645 ;
        RECT 240.855 86.605 241.115 86.695 ;
        RECT 240.455 86.465 241.115 86.605 ;
        RECT 240.855 86.375 241.115 86.465 ;
        RECT 240.385 85.500 240.665 85.870 ;
        RECT 240.395 85.355 240.655 85.500 ;
        RECT 239.005 80.995 239.285 81.110 ;
        RECT 239.005 80.915 239.675 80.995 ;
        RECT 239.935 80.935 240.195 81.255 ;
        RECT 239.005 80.855 239.735 80.915 ;
        RECT 239.005 80.740 239.285 80.855 ;
        RECT 239.475 80.595 239.735 80.855 ;
        RECT 240.455 80.315 240.595 85.355 ;
        RECT 240.845 84.820 241.125 85.190 ;
        RECT 240.915 83.635 241.055 84.820 ;
        RECT 240.855 83.315 241.115 83.635 ;
        RECT 240.455 80.175 241.055 80.315 ;
        RECT 241.375 80.235 241.515 88.505 ;
        RECT 241.835 88.395 241.975 88.845 ;
        RECT 241.775 88.075 242.035 88.395 ;
        RECT 242.235 88.075 242.495 88.395 ;
        RECT 242.295 86.945 242.435 88.075 ;
        RECT 241.835 86.805 242.435 86.945 ;
        RECT 241.835 83.295 241.975 86.805 ;
        RECT 242.755 86.435 242.895 89.435 ;
        RECT 243.155 88.755 243.415 89.075 ;
        RECT 242.295 86.295 242.895 86.435 ;
        RECT 241.775 82.975 242.035 83.295 ;
        RECT 242.295 82.470 242.435 86.295 ;
        RECT 242.695 85.925 242.955 86.015 ;
        RECT 243.215 85.925 243.355 88.755 ;
        RECT 242.695 85.785 243.355 85.925 ;
        RECT 242.695 85.695 242.955 85.785 ;
        RECT 244.135 85.585 244.275 94.195 ;
        RECT 244.595 92.475 244.735 98.615 ;
        RECT 244.995 94.765 245.255 94.855 ;
        RECT 244.995 94.625 245.655 94.765 ;
        RECT 244.995 94.535 245.255 94.625 ;
        RECT 244.995 93.855 245.255 94.175 ;
        RECT 245.055 92.670 245.195 93.855 ;
        RECT 244.535 92.155 244.795 92.475 ;
        RECT 244.985 92.300 245.265 92.670 ;
        RECT 245.515 89.950 245.655 94.625 ;
        RECT 246.435 94.030 246.575 105.075 ;
        RECT 246.895 103.355 247.035 109.225 ;
        RECT 247.755 104.055 248.015 104.375 ;
        RECT 246.835 103.035 247.095 103.355 ;
        RECT 247.815 102.335 247.955 104.055 ;
        RECT 249.195 103.355 249.335 109.225 ;
        RECT 250.055 105.075 250.315 105.395 ;
        RECT 249.135 103.035 249.395 103.355 ;
        RECT 249.125 102.500 249.405 102.870 ;
        RECT 247.755 102.015 248.015 102.335 ;
        RECT 248.675 101.675 248.935 101.995 ;
        RECT 248.735 100.295 248.875 101.675 ;
        RECT 249.195 100.635 249.335 102.500 ;
        RECT 250.115 101.995 250.255 105.075 ;
        RECT 251.495 105.055 251.635 109.225 ;
        RECT 252.815 107.115 253.075 107.435 ;
        RECT 251.435 104.735 251.695 105.055 ;
        RECT 252.875 102.755 253.015 107.115 ;
        RECT 253.795 106.075 253.935 109.225 ;
        RECT 253.735 105.755 253.995 106.075 ;
        RECT 256.095 104.375 256.235 109.225 ;
        RECT 257.875 104.735 258.135 105.055 ;
        RECT 256.035 104.055 256.295 104.375 ;
        RECT 254.475 103.520 256.015 103.890 ;
        RECT 256.035 103.035 256.295 103.355 ;
        RECT 251.955 102.615 253.015 102.755 ;
        RECT 249.595 101.675 249.855 101.995 ;
        RECT 250.055 101.675 250.315 101.995 ;
        RECT 249.135 100.315 249.395 100.635 ;
        RECT 248.675 99.975 248.935 100.295 ;
        RECT 248.735 99.470 248.875 99.975 ;
        RECT 248.665 99.100 248.945 99.470 ;
        RECT 246.825 97.060 247.105 97.430 ;
        RECT 246.365 93.660 246.645 94.030 ;
        RECT 246.375 91.135 246.635 91.455 ;
        RECT 245.445 89.580 245.725 89.950 ;
        RECT 244.535 88.075 244.795 88.395 ;
        RECT 244.595 87.035 244.735 88.075 ;
        RECT 244.995 87.735 245.255 88.055 ;
        RECT 244.535 86.715 244.795 87.035 ;
        RECT 243.215 85.445 244.275 85.585 ;
        RECT 242.695 85.015 242.955 85.335 ;
        RECT 242.755 84.510 242.895 85.015 ;
        RECT 242.685 84.140 242.965 84.510 ;
        RECT 243.215 82.615 243.355 85.445 ;
        RECT 244.535 85.355 244.795 85.675 ;
        RECT 244.595 85.075 244.735 85.355 ;
        RECT 244.135 84.935 244.735 85.075 ;
        RECT 244.135 83.975 244.275 84.935 ;
        RECT 244.525 84.140 244.805 84.510 ;
        RECT 244.075 83.885 244.335 83.975 ;
        RECT 243.675 83.745 244.335 83.885 ;
        RECT 242.225 82.100 242.505 82.470 ;
        RECT 243.155 82.295 243.415 82.615 ;
        RECT 241.765 81.420 242.045 81.790 ;
        RECT 242.295 81.675 242.435 82.100 ;
        RECT 242.295 81.535 242.895 81.675 ;
        RECT 239.475 79.575 239.735 79.895 ;
        RECT 240.395 79.575 240.655 79.895 ;
        RECT 238.555 77.535 238.815 77.855 ;
        RECT 238.095 77.425 238.355 77.515 ;
        RECT 237.695 77.285 238.355 77.425 ;
        RECT 238.095 77.195 238.355 77.285 ;
        RECT 237.625 76.915 237.905 77.030 ;
        RECT 237.235 76.775 237.905 76.915 ;
        RECT 237.235 75.475 237.375 76.775 ;
        RECT 237.625 76.660 237.905 76.775 ;
        RECT 237.175 75.155 237.435 75.475 ;
        RECT 237.635 74.475 237.895 74.795 ;
        RECT 236.715 74.135 236.975 74.455 ;
        RECT 235.845 73.600 237.385 73.970 ;
        RECT 235.395 73.205 237.375 73.345 ;
        RECT 234.865 72.580 235.145 72.950 ;
        RECT 234.935 69.695 235.075 72.580 ;
        RECT 235.795 72.435 236.055 72.755 ;
        RECT 235.855 70.035 235.995 72.435 ;
        RECT 236.255 70.395 236.515 70.715 ;
        RECT 235.795 69.715 236.055 70.035 ;
        RECT 236.315 69.695 236.455 70.395 ;
        RECT 234.875 69.375 235.135 69.695 ;
        RECT 236.255 69.375 236.515 69.695 ;
        RECT 237.235 68.925 237.375 73.205 ;
        RECT 237.695 72.755 237.835 74.475 ;
        RECT 237.635 72.435 237.895 72.755 ;
        RECT 238.155 69.695 238.295 77.195 ;
        RECT 238.615 72.075 238.755 77.535 ;
        RECT 239.015 77.195 239.275 77.515 ;
        RECT 239.075 75.135 239.215 77.195 ;
        RECT 239.535 75.475 239.675 79.575 ;
        RECT 239.925 78.700 240.205 79.070 ;
        RECT 239.935 78.555 240.195 78.700 ;
        RECT 239.935 77.875 240.195 78.195 ;
        RECT 239.995 76.155 240.135 77.875 ;
        RECT 239.935 75.835 240.195 76.155 ;
        RECT 239.475 75.155 239.735 75.475 ;
        RECT 239.015 74.815 239.275 75.135 ;
        RECT 239.015 74.135 239.275 74.455 ;
        RECT 239.475 74.135 239.735 74.455 ;
        RECT 238.555 71.755 238.815 72.075 ;
        RECT 238.095 69.375 238.355 69.695 ;
        RECT 239.075 69.015 239.215 74.135 ;
        RECT 237.235 68.785 237.835 68.925 ;
        RECT 235.845 68.160 237.385 68.530 ;
        RECT 236.715 67.675 236.975 67.995 ;
        RECT 236.775 67.315 236.915 67.675 ;
        RECT 236.255 66.995 236.515 67.315 ;
        RECT 236.715 66.995 236.975 67.315 ;
        RECT 236.315 66.830 236.455 66.995 ;
        RECT 236.245 66.460 236.525 66.830 ;
        RECT 235.845 62.720 237.385 63.090 ;
        RECT 235.325 61.700 235.605 62.070 ;
        RECT 235.335 61.555 235.595 61.700 ;
        RECT 236.715 61.555 236.975 61.875 ;
        RECT 235.335 60.875 235.595 61.195 ;
        RECT 233.555 60.455 234.615 60.595 ;
        RECT 233.495 58.835 233.755 59.155 ;
        RECT 233.555 53.375 233.695 58.835 ;
        RECT 234.475 58.475 234.615 60.455 ;
        RECT 235.395 59.595 235.535 60.875 ;
        RECT 235.395 59.455 235.995 59.595 ;
        RECT 234.415 58.155 234.675 58.475 ;
        RECT 234.875 58.155 235.135 58.475 ;
        RECT 233.955 57.025 234.215 57.115 ;
        RECT 234.935 57.025 235.075 58.155 ;
        RECT 235.855 58.045 235.995 59.455 ;
        RECT 236.775 58.815 236.915 61.555 ;
        RECT 237.175 61.215 237.435 61.535 ;
        RECT 236.715 58.495 236.975 58.815 ;
        RECT 237.235 58.555 237.375 61.215 ;
        RECT 237.695 59.155 237.835 68.785 ;
        RECT 238.095 68.695 238.355 69.015 ;
        RECT 239.015 68.695 239.275 69.015 ;
        RECT 238.155 67.315 238.295 68.695 ;
        RECT 238.095 66.995 238.355 67.315 ;
        RECT 239.015 65.975 239.275 66.295 ;
        RECT 239.075 65.275 239.215 65.975 ;
        RECT 239.015 64.955 239.275 65.275 ;
        RECT 239.535 64.935 239.675 74.135 ;
        RECT 239.935 72.435 240.195 72.755 ;
        RECT 239.995 70.715 240.135 72.435 ;
        RECT 240.455 70.715 240.595 79.575 ;
        RECT 240.915 74.455 241.055 80.175 ;
        RECT 241.315 79.915 241.575 80.235 ;
        RECT 240.855 74.135 241.115 74.455 ;
        RECT 241.375 73.515 241.515 79.915 ;
        RECT 241.835 79.895 241.975 81.420 ;
        RECT 242.235 80.935 242.495 81.255 ;
        RECT 241.775 79.575 242.035 79.895 ;
        RECT 242.295 77.595 242.435 80.935 ;
        RECT 242.755 78.195 242.895 81.535 ;
        RECT 243.675 81.255 243.815 83.745 ;
        RECT 244.075 83.655 244.335 83.745 ;
        RECT 244.075 83.205 244.335 83.295 ;
        RECT 244.595 83.205 244.735 84.140 ;
        RECT 244.075 83.065 244.735 83.205 ;
        RECT 244.075 82.975 244.335 83.065 ;
        RECT 244.535 82.470 244.795 82.615 ;
        RECT 244.525 82.100 244.805 82.470 ;
        RECT 243.615 80.935 243.875 81.255 ;
        RECT 244.075 80.935 244.335 81.255 ;
        RECT 243.615 80.255 243.875 80.575 ;
        RECT 243.155 79.575 243.415 79.895 ;
        RECT 242.695 77.875 242.955 78.195 ;
        RECT 240.915 73.375 241.515 73.515 ;
        RECT 241.835 77.455 242.435 77.595 ;
        RECT 241.835 73.395 241.975 77.455 ;
        RECT 242.235 76.855 242.495 77.175 ;
        RECT 242.295 76.350 242.435 76.855 ;
        RECT 242.225 75.980 242.505 76.350 ;
        RECT 239.935 70.395 240.195 70.715 ;
        RECT 240.395 70.395 240.655 70.715 ;
        RECT 239.925 68.500 240.205 68.870 ;
        RECT 239.995 67.655 240.135 68.500 ;
        RECT 239.935 67.335 240.195 67.655 ;
        RECT 240.455 67.315 240.595 70.395 ;
        RECT 240.915 67.995 241.055 73.375 ;
        RECT 241.835 73.255 242.435 73.395 ;
        RECT 241.775 72.435 242.035 72.755 ;
        RECT 241.315 69.035 241.575 69.355 ;
        RECT 240.855 67.675 241.115 67.995 ;
        RECT 240.395 66.995 240.655 67.315 ;
        RECT 239.475 64.615 239.735 64.935 ;
        RECT 239.535 64.165 239.675 64.615 ;
        RECT 241.375 64.255 241.515 69.035 ;
        RECT 241.835 68.870 241.975 72.435 ;
        RECT 241.765 68.500 242.045 68.870 ;
        RECT 242.295 68.075 242.435 73.255 ;
        RECT 242.755 72.755 242.895 77.875 ;
        RECT 243.215 76.155 243.355 79.575 ;
        RECT 243.155 75.835 243.415 76.155 ;
        RECT 243.675 75.135 243.815 80.255 ;
        RECT 244.135 78.195 244.275 80.935 ;
        RECT 244.535 80.255 244.795 80.575 ;
        RECT 244.075 77.875 244.335 78.195 ;
        RECT 244.595 77.175 244.735 80.255 ;
        RECT 244.535 76.855 244.795 77.175 ;
        RECT 243.615 74.815 243.875 75.135 ;
        RECT 244.075 74.135 244.335 74.455 ;
        RECT 242.695 72.435 242.955 72.755 ;
        RECT 243.155 72.435 243.415 72.755 ;
        RECT 241.835 67.935 242.435 68.075 ;
        RECT 240.395 64.165 240.655 64.255 ;
        RECT 239.535 64.025 240.655 64.165 ;
        RECT 240.395 63.935 240.655 64.025 ;
        RECT 241.315 63.935 241.575 64.255 ;
        RECT 238.095 60.535 238.355 60.855 ;
        RECT 240.395 60.535 240.655 60.855 ;
        RECT 237.635 58.835 237.895 59.155 ;
        RECT 237.235 58.475 237.835 58.555 ;
        RECT 237.235 58.415 237.895 58.475 ;
        RECT 237.635 58.155 237.895 58.415 ;
        RECT 233.955 56.885 235.075 57.025 ;
        RECT 235.395 57.905 235.995 58.045 ;
        RECT 233.955 56.795 234.215 56.885 ;
        RECT 235.395 54.055 235.535 57.905 ;
        RECT 235.845 57.280 237.385 57.650 ;
        RECT 237.695 56.685 237.835 58.155 ;
        RECT 235.855 56.545 237.835 56.685 ;
        RECT 233.945 53.540 234.225 53.910 ;
        RECT 235.335 53.735 235.595 54.055 ;
        RECT 233.955 53.395 234.215 53.540 ;
        RECT 233.495 53.055 233.755 53.375 ;
        RECT 234.015 50.315 234.155 53.395 ;
        RECT 235.855 53.375 235.995 56.545 ;
        RECT 237.175 55.095 237.435 55.415 ;
        RECT 237.235 54.055 237.375 55.095 ;
        RECT 237.175 53.735 237.435 54.055 ;
        RECT 238.155 53.375 238.295 60.535 ;
        RECT 240.455 58.815 240.595 60.535 ;
        RECT 241.375 59.350 241.515 63.935 ;
        RECT 241.835 61.535 241.975 67.935 ;
        RECT 242.235 66.315 242.495 66.635 ;
        RECT 242.695 66.315 242.955 66.635 ;
        RECT 241.775 61.215 242.035 61.535 ;
        RECT 241.305 58.980 241.585 59.350 ;
        RECT 241.835 59.155 241.975 61.215 ;
        RECT 241.775 58.835 242.035 59.155 ;
        RECT 240.395 58.495 240.655 58.815 ;
        RECT 240.855 57.815 241.115 58.135 ;
        RECT 241.315 57.815 241.575 58.135 ;
        RECT 241.775 57.815 242.035 58.135 ;
        RECT 240.915 56.775 241.055 57.815 ;
        RECT 240.855 56.455 241.115 56.775 ;
        RECT 239.475 56.115 239.735 56.435 ;
        RECT 238.555 53.395 238.815 53.715 ;
        RECT 235.795 53.055 236.055 53.375 ;
        RECT 237.175 53.055 237.435 53.375 ;
        RECT 238.095 53.055 238.355 53.375 ;
        RECT 234.415 52.375 234.675 52.695 ;
        RECT 237.235 52.605 237.375 53.055 ;
        RECT 237.235 52.465 237.835 52.605 ;
        RECT 233.955 49.995 234.215 50.315 ;
        RECT 234.475 48.275 234.615 52.375 ;
        RECT 235.845 51.840 237.385 52.210 ;
        RECT 237.695 50.315 237.835 52.465 ;
        RECT 238.095 52.375 238.355 52.695 ;
        RECT 238.155 50.995 238.295 52.375 ;
        RECT 238.095 50.675 238.355 50.995 ;
        RECT 237.635 49.995 237.895 50.315 ;
        RECT 238.615 49.975 238.755 53.395 ;
        RECT 239.535 53.375 239.675 56.115 ;
        RECT 240.395 55.775 240.655 56.095 ;
        RECT 240.455 53.375 240.595 55.775 ;
        RECT 240.855 55.435 241.115 55.755 ;
        RECT 240.915 54.395 241.055 55.435 ;
        RECT 240.855 54.075 241.115 54.395 ;
        RECT 239.475 53.055 239.735 53.375 ;
        RECT 240.395 53.055 240.655 53.375 ;
        RECT 240.855 53.230 241.115 53.375 ;
        RECT 240.845 52.860 241.125 53.230 ;
        RECT 241.375 50.995 241.515 57.815 ;
        RECT 241.835 53.375 241.975 57.815 ;
        RECT 241.775 53.055 242.035 53.375 ;
        RECT 242.295 51.675 242.435 66.315 ;
        RECT 242.755 66.150 242.895 66.315 ;
        RECT 242.685 65.780 242.965 66.150 ;
        RECT 243.215 64.935 243.355 72.435 ;
        RECT 243.615 71.755 243.875 72.075 ;
        RECT 243.675 69.355 243.815 71.755 ;
        RECT 243.615 69.035 243.875 69.355 ;
        RECT 243.155 64.615 243.415 64.935 ;
        RECT 242.695 56.115 242.955 56.435 ;
        RECT 242.755 55.270 242.895 56.115 ;
        RECT 243.675 56.095 243.815 69.035 ;
        RECT 244.135 56.435 244.275 74.135 ;
        RECT 245.055 73.395 245.195 87.735 ;
        RECT 245.515 86.355 245.655 89.580 ;
        RECT 245.455 86.035 245.715 86.355 ;
        RECT 245.455 85.015 245.715 85.335 ;
        RECT 245.515 83.635 245.655 85.015 ;
        RECT 245.455 83.315 245.715 83.635 ;
        RECT 245.915 82.295 246.175 82.615 ;
        RECT 245.455 80.935 245.715 81.255 ;
        RECT 245.515 80.575 245.655 80.935 ;
        RECT 245.455 80.255 245.715 80.575 ;
        RECT 245.975 79.750 246.115 82.295 ;
        RECT 246.435 80.575 246.575 91.135 ;
        RECT 246.375 80.255 246.635 80.575 ;
        RECT 246.895 80.315 247.035 97.060 ;
        RECT 247.295 96.575 247.555 96.895 ;
        RECT 247.355 93.495 247.495 96.575 ;
        RECT 247.295 93.175 247.555 93.495 ;
        RECT 248.215 90.455 248.475 90.775 ;
        RECT 248.275 83.975 248.415 90.455 ;
        RECT 248.675 83.995 248.935 84.315 ;
        RECT 248.215 83.655 248.475 83.975 ;
        RECT 247.295 83.545 247.555 83.635 ;
        RECT 247.295 83.405 247.955 83.545 ;
        RECT 247.295 83.315 247.555 83.405 ;
        RECT 247.815 80.915 247.955 83.405 ;
        RECT 248.215 82.975 248.475 83.295 ;
        RECT 248.275 81.595 248.415 82.975 ;
        RECT 248.215 81.275 248.475 81.595 ;
        RECT 247.755 80.595 248.015 80.915 ;
        RECT 246.895 80.175 247.495 80.315 ;
        RECT 245.905 79.380 246.185 79.750 ;
        RECT 246.835 79.575 247.095 79.895 ;
        RECT 245.515 78.875 246.575 78.955 ;
        RECT 245.455 78.815 246.575 78.875 ;
        RECT 245.455 78.555 245.715 78.815 ;
        RECT 246.435 78.535 246.575 78.815 ;
        RECT 246.375 78.215 246.635 78.535 ;
        RECT 245.455 77.875 245.715 78.195 ;
        RECT 245.515 75.815 245.655 77.875 ;
        RECT 245.455 75.495 245.715 75.815 ;
        RECT 246.895 75.475 247.035 79.575 ;
        RECT 247.355 78.875 247.495 80.175 ;
        RECT 248.215 79.915 248.475 80.235 ;
        RECT 247.295 78.555 247.555 78.875 ;
        RECT 247.755 78.555 248.015 78.875 ;
        RECT 246.835 75.155 247.095 75.475 ;
        RECT 245.915 74.815 246.175 75.135 ;
        RECT 245.055 73.255 245.655 73.395 ;
        RECT 244.535 69.035 244.795 69.355 ;
        RECT 244.595 56.435 244.735 69.035 ;
        RECT 244.995 58.835 245.255 59.155 ;
        RECT 244.075 56.115 244.335 56.435 ;
        RECT 244.535 56.115 244.795 56.435 ;
        RECT 243.615 55.775 243.875 56.095 ;
        RECT 242.685 54.900 242.965 55.270 ;
        RECT 244.135 53.375 244.275 56.115 ;
        RECT 245.055 55.415 245.195 58.835 ;
        RECT 244.995 55.095 245.255 55.415 ;
        RECT 245.515 53.795 245.655 73.255 ;
        RECT 245.975 58.135 246.115 74.815 ;
        RECT 247.355 74.795 247.495 78.555 ;
        RECT 247.815 77.030 247.955 78.555 ;
        RECT 247.745 76.660 248.025 77.030 ;
        RECT 247.295 74.475 247.555 74.795 ;
        RECT 246.825 71.900 247.105 72.270 ;
        RECT 246.375 68.695 246.635 69.015 ;
        RECT 245.915 57.815 246.175 58.135 ;
        RECT 246.435 55.415 246.575 68.695 ;
        RECT 246.375 55.095 246.635 55.415 ;
        RECT 245.515 53.715 246.575 53.795 ;
        RECT 246.895 53.715 247.035 71.900 ;
        RECT 247.295 69.715 247.555 70.035 ;
        RECT 247.355 64.790 247.495 69.715 ;
        RECT 248.275 69.355 248.415 79.915 ;
        RECT 248.735 78.535 248.875 83.995 ;
        RECT 249.135 82.635 249.395 82.955 ;
        RECT 249.195 82.470 249.335 82.635 ;
        RECT 249.655 82.615 249.795 101.675 ;
        RECT 250.515 101.335 250.775 101.655 ;
        RECT 250.575 100.295 250.715 101.335 ;
        RECT 250.515 99.975 250.775 100.295 ;
        RECT 251.955 91.455 252.095 102.615 ;
        RECT 252.875 102.335 253.015 102.615 ;
        RECT 252.355 102.015 252.615 102.335 ;
        RECT 252.815 102.015 253.075 102.335 ;
        RECT 253.275 102.015 253.535 102.335 ;
        RECT 252.415 99.955 252.555 102.015 ;
        RECT 252.355 99.635 252.615 99.955 ;
        RECT 252.815 99.635 253.075 99.955 ;
        RECT 252.415 99.275 252.555 99.635 ;
        RECT 252.355 98.955 252.615 99.275 ;
        RECT 252.875 98.110 253.015 99.635 ;
        RECT 252.805 97.740 253.085 98.110 ;
        RECT 253.335 96.635 253.475 102.015 ;
        RECT 254.655 101.675 254.915 101.995 ;
        RECT 253.735 100.315 253.995 100.635 ;
        RECT 253.795 96.895 253.935 100.315 ;
        RECT 254.715 100.295 254.855 101.675 ;
        RECT 255.105 100.715 255.385 100.830 ;
        RECT 256.095 100.715 256.235 103.035 ;
        RECT 256.955 101.335 257.215 101.655 ;
        RECT 257.415 101.335 257.675 101.655 ;
        RECT 255.105 100.575 256.235 100.715 ;
        RECT 255.105 100.460 255.385 100.575 ;
        RECT 254.655 99.975 254.915 100.295 ;
        RECT 255.635 99.955 255.775 100.575 ;
        RECT 256.485 100.460 256.765 100.830 ;
        RECT 254.195 99.635 254.455 99.955 ;
        RECT 255.575 99.635 255.835 99.955 ;
        RECT 254.255 99.355 254.395 99.635 ;
        RECT 256.555 99.355 256.695 100.460 ;
        RECT 257.015 100.295 257.155 101.335 ;
        RECT 256.955 99.975 257.215 100.295 ;
        RECT 254.255 99.215 256.695 99.355 ;
        RECT 257.475 98.675 257.615 101.335 ;
        RECT 257.935 100.995 258.075 104.735 ;
        RECT 258.395 103.435 258.535 109.225 ;
        RECT 260.695 106.075 260.835 109.225 ;
        RECT 262.995 106.075 263.135 109.225 ;
        RECT 265.295 107.435 265.435 109.225 ;
        RECT 265.235 107.115 265.495 107.435 ;
        RECT 267.075 106.775 267.335 107.095 ;
        RECT 260.635 105.755 260.895 106.075 ;
        RECT 262.935 105.755 263.195 106.075 ;
        RECT 262.015 105.415 262.275 105.735 ;
        RECT 259.715 105.075 259.975 105.395 ;
        RECT 258.395 103.355 258.995 103.435 ;
        RECT 258.395 103.295 259.055 103.355 ;
        RECT 258.795 103.035 259.055 103.295 ;
        RECT 259.775 101.510 259.915 105.075 ;
        RECT 260.635 104.395 260.895 104.715 ;
        RECT 260.695 103.015 260.835 104.395 ;
        RECT 260.635 102.695 260.895 103.015 ;
        RECT 260.175 101.675 260.435 101.995 ;
        RECT 259.705 101.140 259.985 101.510 ;
        RECT 257.935 100.855 258.535 100.995 ;
        RECT 257.015 98.535 257.615 98.675 ;
        RECT 257.875 98.615 258.135 98.935 ;
        RECT 254.475 98.080 256.015 98.450 ;
        RECT 257.015 97.315 257.155 98.535 ;
        RECT 257.405 97.740 257.685 98.110 ;
        RECT 257.475 97.575 257.615 97.740 ;
        RECT 254.195 96.915 254.455 97.235 ;
        RECT 255.635 97.175 257.155 97.315 ;
        RECT 257.415 97.255 257.675 97.575 ;
        RECT 252.875 96.495 253.475 96.635 ;
        RECT 253.735 96.575 253.995 96.895 ;
        RECT 251.895 91.135 252.155 91.455 ;
        RECT 250.055 86.375 250.315 86.695 ;
        RECT 249.125 82.100 249.405 82.470 ;
        RECT 249.595 82.295 249.855 82.615 ;
        RECT 248.675 78.215 248.935 78.535 ;
        RECT 248.675 76.855 248.935 77.175 ;
        RECT 248.735 75.135 248.875 76.855 ;
        RECT 248.675 74.815 248.935 75.135 ;
        RECT 248.675 74.135 248.935 74.455 ;
        RECT 248.735 73.435 248.875 74.135 ;
        RECT 248.675 73.115 248.935 73.435 ;
        RECT 248.215 69.035 248.475 69.355 ;
        RECT 248.275 65.470 248.415 69.035 ;
        RECT 248.675 66.995 248.935 67.315 ;
        RECT 248.205 65.100 248.485 65.470 ;
        RECT 247.285 64.420 247.565 64.790 ;
        RECT 247.295 58.495 247.555 58.815 ;
        RECT 247.355 57.115 247.495 58.495 ;
        RECT 247.745 58.300 248.025 58.670 ;
        RECT 247.755 58.155 248.015 58.300 ;
        RECT 247.295 56.795 247.555 57.115 ;
        RECT 248.215 56.115 248.475 56.435 ;
        RECT 248.275 54.395 248.415 56.115 ;
        RECT 248.215 54.075 248.475 54.395 ;
        RECT 244.995 53.395 245.255 53.715 ;
        RECT 245.515 53.655 246.635 53.715 ;
        RECT 246.375 53.395 246.635 53.655 ;
        RECT 246.835 53.395 247.095 53.715 ;
        RECT 244.075 53.055 244.335 53.375 ;
        RECT 242.235 51.355 242.495 51.675 ;
        RECT 241.315 50.675 241.575 50.995 ;
        RECT 243.155 50.675 243.415 50.995 ;
        RECT 238.555 49.655 238.815 49.975 ;
        RECT 240.395 49.655 240.655 49.975 ;
        RECT 240.455 48.275 240.595 49.655 ;
        RECT 243.215 48.955 243.355 50.675 ;
        RECT 243.155 48.635 243.415 48.955 ;
        RECT 234.415 47.955 234.675 48.275 ;
        RECT 240.395 47.955 240.655 48.275 ;
        RECT 239.015 47.615 239.275 47.935 ;
        RECT 234.415 46.935 234.675 47.255 ;
        RECT 233.035 45.235 233.295 45.555 ;
        RECT 231.655 44.895 231.915 45.215 ;
        RECT 230.735 43.195 230.995 43.515 ;
        RECT 232.575 43.195 232.835 43.515 ;
        RECT 229.815 40.475 230.075 40.795 ;
        RECT 230.275 40.475 230.535 40.795 ;
        RECT 228.895 39.795 229.155 40.115 ;
        RECT 227.975 38.775 228.235 39.095 ;
        RECT 228.435 38.775 228.695 39.095 ;
        RECT 228.955 38.075 229.095 39.795 ;
        RECT 228.895 37.755 229.155 38.075 ;
        RECT 229.875 35.015 230.015 40.475 ;
        RECT 232.635 37.055 232.775 43.195 ;
        RECT 233.495 42.515 233.755 42.835 ;
        RECT 233.555 42.155 233.695 42.515 ;
        RECT 233.495 41.835 233.755 42.155 ;
        RECT 230.275 36.735 230.535 37.055 ;
        RECT 232.575 36.735 232.835 37.055 ;
        RECT 222.915 34.695 223.175 35.015 ;
        RECT 227.515 34.695 227.775 35.015 ;
        RECT 229.815 34.695 230.075 35.015 ;
        RECT 221.995 34.245 222.255 34.335 ;
        RECT 221.135 34.105 222.255 34.245 ;
        RECT 220.615 32.315 220.875 32.635 ;
        RECT 220.615 29.145 220.875 29.235 ;
        RECT 220.215 29.005 220.875 29.145 ;
        RECT 220.615 28.915 220.875 29.005 ;
        RECT 221.135 28.555 221.275 34.105 ;
        RECT 221.995 34.015 222.255 34.105 ;
        RECT 222.975 29.915 223.115 34.695 ;
        RECT 224.295 34.355 224.555 34.675 ;
        RECT 224.355 33.655 224.495 34.355 ;
        RECT 227.055 34.015 227.315 34.335 ;
        RECT 224.295 33.335 224.555 33.655 ;
        RECT 227.115 32.635 227.255 34.015 ;
        RECT 227.055 32.315 227.315 32.635 ;
        RECT 227.575 31.275 227.715 34.695 ;
        RECT 229.355 34.015 229.615 34.335 ;
        RECT 228.895 33.675 229.155 33.995 ;
        RECT 228.955 32.295 229.095 33.675 ;
        RECT 228.895 31.975 229.155 32.295 ;
        RECT 227.515 30.955 227.775 31.275 ;
        RECT 222.915 29.595 223.175 29.915 ;
        RECT 228.955 28.895 229.095 31.975 ;
        RECT 229.415 31.955 229.555 34.015 ;
        RECT 229.355 31.635 229.615 31.955 ;
        RECT 230.335 30.935 230.475 36.735 ;
        RECT 230.275 30.615 230.535 30.935 ;
        RECT 232.635 29.915 232.775 36.735 ;
        RECT 233.555 31.470 233.695 41.835 ;
        RECT 234.475 40.795 234.615 46.935 ;
        RECT 235.845 46.400 237.385 46.770 ;
        RECT 239.075 45.215 239.215 47.615 ;
        RECT 242.695 47.275 242.955 47.595 ;
        RECT 242.755 46.235 242.895 47.275 ;
        RECT 242.695 45.915 242.955 46.235 ;
        RECT 245.055 45.215 245.195 53.395 ;
        RECT 247.295 53.055 247.555 53.375 ;
        RECT 247.355 45.215 247.495 53.055 ;
        RECT 247.755 49.995 248.015 50.315 ;
        RECT 247.815 48.955 247.955 49.995 ;
        RECT 247.755 48.635 248.015 48.955 ;
        RECT 239.015 44.895 239.275 45.215 ;
        RECT 241.775 44.895 242.035 45.215 ;
        RECT 244.995 44.895 245.255 45.215 ;
        RECT 247.295 44.895 247.555 45.215 ;
        RECT 239.075 42.835 239.215 44.895 ;
        RECT 239.015 42.515 239.275 42.835 ;
        RECT 240.395 42.175 240.655 42.495 ;
        RECT 234.875 41.495 235.135 41.815 ;
        RECT 234.935 40.795 235.075 41.495 ;
        RECT 235.845 40.960 237.385 41.330 ;
        RECT 234.415 40.475 234.675 40.795 ;
        RECT 234.875 40.475 235.135 40.795 ;
        RECT 234.935 37.395 235.075 40.475 ;
        RECT 238.545 38.580 238.825 38.950 ;
        RECT 234.875 37.075 235.135 37.395 ;
        RECT 238.615 37.055 238.755 38.580 ;
        RECT 238.555 36.910 238.815 37.055 ;
        RECT 238.545 36.540 238.825 36.910 ;
        RECT 238.095 36.055 238.355 36.375 ;
        RECT 235.845 35.520 237.385 35.890 ;
        RECT 238.155 35.355 238.295 36.055 ;
        RECT 240.455 35.355 240.595 42.175 ;
        RECT 241.835 40.795 241.975 44.895 ;
        RECT 247.355 42.495 247.495 44.895 ;
        RECT 247.295 42.175 247.555 42.495 ;
        RECT 241.775 40.475 242.035 40.795 ;
        RECT 240.855 39.455 241.115 39.775 ;
        RECT 247.755 39.455 248.015 39.775 ;
        RECT 240.915 38.075 241.055 39.455 ;
        RECT 244.535 38.775 244.795 39.095 ;
        RECT 240.855 37.755 241.115 38.075 ;
        RECT 241.775 37.075 242.035 37.395 ;
        RECT 241.835 35.355 241.975 37.075 ;
        RECT 242.235 36.055 242.495 36.375 ;
        RECT 238.095 35.035 238.355 35.355 ;
        RECT 240.395 35.035 240.655 35.355 ;
        RECT 241.775 35.035 242.035 35.355 ;
        RECT 233.955 33.335 234.215 33.655 ;
        RECT 233.485 31.100 233.765 31.470 ;
        RECT 233.555 30.935 233.695 31.100 ;
        RECT 233.495 30.615 233.755 30.935 ;
        RECT 232.575 29.595 232.835 29.915 ;
        RECT 228.895 28.575 229.155 28.895 ;
        RECT 233.555 28.555 233.695 30.615 ;
        RECT 234.015 29.915 234.155 33.335 ;
        RECT 238.155 31.615 238.295 35.035 ;
        RECT 242.295 34.675 242.435 36.055 ;
        RECT 244.595 35.355 244.735 38.775 ;
        RECT 247.815 38.075 247.955 39.455 ;
        RECT 247.755 37.755 248.015 38.075 ;
        RECT 244.535 35.035 244.795 35.355 ;
        RECT 242.235 34.355 242.495 34.675 ;
        RECT 243.615 34.015 243.875 34.335 ;
        RECT 243.675 32.635 243.815 34.015 ;
        RECT 243.615 32.315 243.875 32.635 ;
        RECT 236.255 31.470 236.515 31.615 ;
        RECT 234.415 30.955 234.675 31.275 ;
        RECT 236.245 31.100 236.525 31.470 ;
        RECT 238.095 31.295 238.355 31.615 ;
        RECT 233.955 29.595 234.215 29.915 ;
        RECT 221.075 28.235 221.335 28.555 ;
        RECT 233.495 28.235 233.755 28.555 ;
        RECT 234.475 28.215 234.615 30.955 ;
        RECT 247.815 30.935 247.955 37.755 ;
        RECT 247.755 30.615 248.015 30.935 ;
        RECT 235.845 30.080 237.385 30.450 ;
        RECT 206.355 27.895 206.615 28.215 ;
        RECT 234.415 27.895 234.675 28.215 ;
        RECT 217.215 27.360 218.755 27.730 ;
        RECT 205.435 26.875 205.695 27.195 ;
        RECT 204.055 25.855 204.315 26.175 ;
        RECT 199.915 25.515 200.175 25.835 ;
        RECT 10.170 23.510 74.550 25.010 ;
        RECT 79.810 23.665 127.975 24.765 ;
        RECT 198.585 24.640 200.125 25.010 ;
        RECT 235.845 24.640 237.385 25.010 ;
        RECT 10.170 21.510 74.550 23.010 ;
        RECT 79.810 22.165 127.975 23.265 ;
        RECT 179.955 21.920 181.495 22.290 ;
        RECT 217.215 21.920 218.755 22.290 ;
        RECT 79.810 20.665 127.975 21.765 ;
        RECT 248.735 20.590 248.875 66.995 ;
        RECT 249.595 65.975 249.855 66.295 ;
        RECT 249.655 64.255 249.795 65.975 ;
        RECT 249.595 63.935 249.855 64.255 ;
        RECT 250.115 61.955 250.255 86.375 ;
        RECT 252.875 85.335 253.015 96.495 ;
        RECT 254.255 96.070 254.395 96.915 ;
        RECT 255.635 96.895 255.775 97.175 ;
        RECT 257.935 96.975 258.075 98.615 ;
        RECT 255.575 96.575 255.835 96.895 ;
        RECT 256.495 96.575 256.755 96.895 ;
        RECT 257.875 96.655 258.135 96.975 ;
        RECT 254.185 95.700 254.465 96.070 ;
        RECT 255.635 94.175 255.775 96.575 ;
        RECT 256.035 96.235 256.295 96.555 ;
        RECT 255.575 93.855 255.835 94.175 ;
        RECT 256.095 93.405 256.235 96.235 ;
        RECT 256.555 94.175 256.695 96.575 ;
        RECT 257.935 94.515 258.075 96.655 ;
        RECT 257.875 94.195 258.135 94.515 ;
        RECT 256.495 93.855 256.755 94.175 ;
        RECT 258.395 93.835 258.535 100.855 ;
        RECT 259.715 100.315 259.975 100.635 ;
        RECT 259.775 96.895 259.915 100.315 ;
        RECT 260.235 99.955 260.375 101.675 ;
        RECT 260.175 99.635 260.435 99.955 ;
        RECT 260.235 97.430 260.375 99.635 ;
        RECT 260.695 98.790 260.835 102.695 ;
        RECT 261.095 102.015 261.355 102.335 ;
        RECT 261.155 99.955 261.295 102.015 ;
        RECT 261.545 100.460 261.825 100.830 ;
        RECT 261.095 99.635 261.355 99.955 ;
        RECT 260.625 98.420 260.905 98.790 ;
        RECT 261.095 98.615 261.355 98.935 ;
        RECT 260.695 97.575 260.835 98.420 ;
        RECT 260.165 97.060 260.445 97.430 ;
        RECT 260.635 97.255 260.895 97.575 ;
        RECT 261.155 97.430 261.295 98.615 ;
        RECT 261.085 97.060 261.365 97.430 ;
        RECT 261.615 96.895 261.755 100.460 ;
        RECT 259.715 96.575 259.975 96.895 ;
        RECT 260.175 96.575 260.435 96.895 ;
        RECT 261.555 96.575 261.815 96.895 ;
        RECT 259.245 95.020 259.525 95.390 ;
        RECT 259.315 94.515 259.455 95.020 ;
        RECT 258.795 94.195 259.055 94.515 ;
        RECT 259.255 94.195 259.515 94.515 ;
        RECT 258.335 93.515 258.595 93.835 ;
        RECT 256.095 93.265 256.695 93.405 ;
        RECT 254.475 92.640 256.015 93.010 ;
        RECT 256.555 89.155 256.695 93.265 ;
        RECT 258.395 89.415 258.535 93.515 ;
        RECT 258.855 89.755 258.995 94.195 ;
        RECT 259.255 93.515 259.515 93.835 ;
        RECT 259.315 91.455 259.455 93.515 ;
        RECT 259.775 91.705 259.915 96.575 ;
        RECT 260.235 94.710 260.375 96.575 ;
        RECT 260.635 96.235 260.895 96.555 ;
        RECT 260.165 94.340 260.445 94.710 ;
        RECT 260.175 94.195 260.435 94.340 ;
        RECT 260.695 93.835 260.835 96.235 ;
        RECT 261.095 95.895 261.355 96.215 ;
        RECT 260.635 93.515 260.895 93.835 ;
        RECT 259.775 91.565 260.835 91.705 ;
        RECT 259.255 91.135 259.515 91.455 ;
        RECT 258.795 89.435 259.055 89.755 ;
        RECT 253.275 88.755 253.535 89.075 ;
        RECT 255.115 88.985 255.375 89.075 ;
        RECT 256.095 89.015 256.695 89.155 ;
        RECT 258.335 89.095 258.595 89.415 ;
        RECT 256.095 88.985 256.235 89.015 ;
        RECT 255.115 88.845 256.235 88.985 ;
        RECT 255.115 88.755 255.375 88.845 ;
        RECT 257.415 88.755 257.675 89.075 ;
        RECT 257.875 88.755 258.135 89.075 ;
        RECT 253.335 85.675 253.475 88.755 ;
        RECT 256.495 88.415 256.755 88.735 ;
        RECT 254.475 87.200 256.015 87.570 ;
        RECT 256.555 87.035 256.695 88.415 ;
        RECT 256.955 87.735 257.215 88.055 ;
        RECT 256.495 86.715 256.755 87.035 ;
        RECT 257.015 86.015 257.155 87.735 ;
        RECT 253.735 85.695 253.995 86.015 ;
        RECT 256.955 85.695 257.215 86.015 ;
        RECT 257.475 85.925 257.615 88.755 ;
        RECT 257.935 86.435 258.075 88.755 ;
        RECT 258.335 88.075 258.595 88.395 ;
        RECT 258.395 87.115 258.535 88.075 ;
        RECT 258.395 86.975 258.995 87.115 ;
        RECT 257.935 86.295 258.535 86.435 ;
        RECT 258.855 86.355 258.995 86.975 ;
        RECT 257.875 85.925 258.135 86.015 ;
        RECT 257.475 85.785 258.135 85.925 ;
        RECT 253.275 85.355 253.535 85.675 ;
        RECT 252.815 85.015 253.075 85.335 ;
        RECT 253.335 85.190 253.475 85.355 ;
        RECT 251.435 83.315 251.695 83.635 ;
        RECT 251.495 80.915 251.635 83.315 ;
        RECT 252.875 83.295 253.015 85.015 ;
        RECT 253.265 84.820 253.545 85.190 ;
        RECT 252.815 82.975 253.075 83.295 ;
        RECT 252.345 81.420 252.625 81.790 ;
        RECT 251.435 80.595 251.695 80.915 ;
        RECT 250.515 77.535 250.775 77.855 ;
        RECT 250.575 70.910 250.715 77.535 ;
        RECT 250.975 75.835 251.235 76.155 ;
        RECT 250.505 70.540 250.785 70.910 ;
        RECT 250.575 67.315 250.715 70.540 ;
        RECT 251.035 69.015 251.175 75.835 ;
        RECT 250.975 68.695 251.235 69.015 ;
        RECT 250.515 66.995 250.775 67.315 ;
        RECT 249.195 61.875 250.715 61.955 ;
        RECT 249.195 61.815 250.775 61.875 ;
        RECT 249.195 59.155 249.335 61.815 ;
        RECT 250.515 61.555 250.775 61.815 ;
        RECT 250.055 61.215 250.315 61.535 ;
        RECT 249.135 58.835 249.395 59.155 ;
        RECT 250.115 58.475 250.255 61.215 ;
        RECT 251.495 59.835 251.635 80.595 ;
        RECT 251.895 80.255 252.155 80.575 ;
        RECT 251.955 70.035 252.095 80.255 ;
        RECT 251.895 69.715 252.155 70.035 ;
        RECT 252.415 66.975 252.555 81.420 ;
        RECT 253.795 80.915 253.935 85.695 ;
        RECT 256.495 85.015 256.755 85.335 ;
        RECT 256.955 85.015 257.215 85.335 ;
        RECT 254.475 81.760 256.015 82.130 ;
        RECT 253.735 80.595 253.995 80.915 ;
        RECT 253.795 80.315 253.935 80.595 ;
        RECT 253.335 80.175 253.935 80.315 ;
        RECT 253.335 72.155 253.475 80.175 ;
        RECT 256.025 80.060 256.305 80.430 ;
        RECT 256.095 78.875 256.235 80.060 ;
        RECT 256.555 79.070 256.695 85.015 ;
        RECT 257.015 83.150 257.155 85.015 ;
        RECT 256.945 82.780 257.225 83.150 ;
        RECT 256.945 81.420 257.225 81.790 ;
        RECT 256.035 78.555 256.295 78.875 ;
        RECT 256.485 78.700 256.765 79.070 ;
        RECT 256.555 78.195 256.695 78.700 ;
        RECT 256.495 77.875 256.755 78.195 ;
        RECT 254.475 76.320 256.015 76.690 ;
        RECT 257.015 75.385 257.155 81.420 ;
        RECT 257.475 78.195 257.615 85.785 ;
        RECT 257.875 85.695 258.135 85.785 ;
        RECT 258.395 84.315 258.535 86.295 ;
        RECT 258.795 86.035 259.055 86.355 ;
        RECT 258.335 83.995 258.595 84.315 ;
        RECT 258.335 82.295 258.595 82.615 ;
        RECT 257.875 80.255 258.135 80.575 ;
        RECT 257.415 77.875 257.675 78.195 ;
        RECT 257.015 75.245 257.615 75.385 ;
        RECT 253.735 74.815 253.995 75.135 ;
        RECT 252.875 72.015 253.475 72.155 ;
        RECT 252.355 66.655 252.615 66.975 ;
        RECT 252.415 63.915 252.555 66.655 ;
        RECT 252.355 63.595 252.615 63.915 ;
        RECT 251.895 63.255 252.155 63.575 ;
        RECT 251.435 59.515 251.695 59.835 ;
        RECT 250.515 59.175 250.775 59.495 ;
        RECT 250.055 58.155 250.315 58.475 ;
        RECT 249.135 57.815 249.395 58.135 ;
        RECT 249.595 57.815 249.855 58.135 ;
        RECT 249.195 56.435 249.335 57.815 ;
        RECT 249.135 56.115 249.395 56.435 ;
        RECT 249.195 53.035 249.335 56.115 ;
        RECT 249.655 55.755 249.795 57.815 ;
        RECT 250.055 55.950 250.315 56.095 ;
        RECT 249.595 55.435 249.855 55.755 ;
        RECT 250.045 55.580 250.325 55.950 ;
        RECT 250.575 55.755 250.715 59.175 ;
        RECT 250.975 58.155 251.235 58.475 ;
        RECT 251.035 56.095 251.175 58.155 ;
        RECT 250.975 55.775 251.235 56.095 ;
        RECT 250.515 55.435 250.775 55.755 ;
        RECT 249.655 54.395 249.795 55.435 ;
        RECT 250.975 55.155 251.235 55.415 ;
        RECT 251.495 55.155 251.635 59.515 ;
        RECT 251.955 58.815 252.095 63.255 ;
        RECT 252.875 59.495 253.015 72.015 ;
        RECT 253.275 71.590 253.535 71.735 ;
        RECT 253.265 71.220 253.545 71.590 ;
        RECT 253.335 69.695 253.475 71.220 ;
        RECT 253.795 70.115 253.935 74.815 ;
        RECT 256.955 74.475 257.215 74.795 ;
        RECT 256.035 72.435 256.295 72.755 ;
        RECT 257.015 72.665 257.155 74.475 ;
        RECT 257.475 73.345 257.615 75.245 ;
        RECT 257.935 74.990 258.075 80.255 ;
        RECT 258.395 78.535 258.535 82.295 ;
        RECT 259.315 81.790 259.455 91.135 ;
        RECT 260.695 89.415 260.835 91.565 ;
        RECT 261.155 91.455 261.295 95.895 ;
        RECT 261.555 94.195 261.815 94.515 ;
        RECT 261.095 91.135 261.355 91.455 ;
        RECT 260.635 89.095 260.895 89.415 ;
        RECT 260.635 88.415 260.895 88.735 ;
        RECT 260.165 87.540 260.445 87.910 ;
        RECT 260.235 86.015 260.375 87.540 ;
        RECT 260.175 85.695 260.435 86.015 ;
        RECT 260.695 85.245 260.835 88.415 ;
        RECT 261.095 87.735 261.355 88.055 ;
        RECT 260.235 85.105 260.835 85.245 ;
        RECT 260.235 84.315 260.375 85.105 ;
        RECT 260.625 84.395 260.905 84.510 ;
        RECT 261.155 84.395 261.295 87.735 ;
        RECT 261.615 85.335 261.755 94.195 ;
        RECT 261.555 85.015 261.815 85.335 ;
        RECT 260.175 83.995 260.435 84.315 ;
        RECT 260.625 84.255 261.295 84.395 ;
        RECT 260.625 84.140 260.905 84.255 ;
        RECT 259.245 81.420 259.525 81.790 ;
        RECT 259.255 80.255 259.515 80.575 ;
        RECT 258.335 78.215 258.595 78.535 ;
        RECT 259.315 78.445 259.455 80.255 ;
        RECT 259.705 78.700 259.985 79.070 ;
        RECT 259.715 78.555 259.975 78.700 ;
        RECT 259.085 78.305 259.455 78.445 ;
        RECT 257.865 74.620 258.145 74.990 ;
        RECT 257.475 73.205 258.075 73.345 ;
        RECT 257.415 72.665 257.675 72.755 ;
        RECT 257.015 72.525 257.675 72.665 ;
        RECT 257.415 72.435 257.675 72.525 ;
        RECT 256.095 72.155 256.235 72.435 ;
        RECT 256.095 72.015 256.695 72.155 ;
        RECT 254.475 70.880 256.015 71.250 ;
        RECT 256.025 70.115 256.305 70.230 ;
        RECT 256.555 70.115 256.695 72.015 ;
        RECT 257.935 70.715 258.075 73.205 ;
        RECT 258.395 70.715 258.535 78.215 ;
        RECT 259.085 77.765 259.225 78.305 ;
        RECT 259.085 77.625 259.455 77.765 ;
        RECT 258.795 77.030 259.055 77.175 ;
        RECT 258.785 76.660 259.065 77.030 ;
        RECT 259.315 75.815 259.455 77.625 ;
        RECT 260.235 77.030 260.375 83.995 ;
        RECT 260.695 80.575 260.835 84.140 ;
        RECT 261.095 83.150 261.355 83.295 ;
        RECT 261.085 82.780 261.365 83.150 ;
        RECT 261.555 82.975 261.815 83.295 ;
        RECT 261.615 81.595 261.755 82.975 ;
        RECT 261.555 81.275 261.815 81.595 ;
        RECT 260.635 80.485 260.895 80.575 ;
        RECT 260.635 80.345 261.295 80.485 ;
        RECT 260.635 80.255 260.895 80.345 ;
        RECT 260.635 79.575 260.895 79.895 ;
        RECT 260.165 76.660 260.445 77.030 ;
        RECT 259.255 75.495 259.515 75.815 ;
        RECT 259.315 75.135 259.455 75.495 ;
        RECT 260.695 75.135 260.835 79.575 ;
        RECT 261.155 78.535 261.295 80.345 ;
        RECT 261.095 78.215 261.355 78.535 ;
        RECT 261.095 77.535 261.355 77.855 ;
        RECT 261.155 76.155 261.295 77.535 ;
        RECT 261.095 75.835 261.355 76.155 ;
        RECT 259.255 74.815 259.515 75.135 ;
        RECT 258.795 74.475 259.055 74.795 ;
        RECT 259.705 74.620 259.985 74.990 ;
        RECT 260.635 74.815 260.895 75.135 ;
        RECT 261.095 74.815 261.355 75.135 ;
        RECT 258.855 71.735 258.995 74.475 ;
        RECT 258.795 71.415 259.055 71.735 ;
        RECT 257.875 70.395 258.135 70.715 ;
        RECT 258.335 70.395 258.595 70.715 ;
        RECT 257.935 70.115 258.075 70.395 ;
        RECT 253.795 69.975 254.855 70.115 ;
        RECT 254.715 69.695 254.855 69.975 ;
        RECT 256.025 69.975 256.695 70.115 ;
        RECT 257.475 69.975 258.075 70.115 ;
        RECT 256.025 69.860 256.305 69.975 ;
        RECT 253.275 69.375 253.535 69.695 ;
        RECT 254.655 69.375 254.915 69.695 ;
        RECT 253.275 68.695 253.535 69.015 ;
        RECT 253.335 64.595 253.475 68.695 ;
        RECT 256.095 67.655 256.235 69.860 ;
        RECT 256.035 67.335 256.295 67.655 ;
        RECT 257.475 67.315 257.615 69.975 ;
        RECT 257.875 69.375 258.135 69.695 ;
        RECT 257.935 67.995 258.075 69.375 ;
        RECT 257.875 67.675 258.135 67.995 ;
        RECT 258.395 67.655 258.535 70.395 ;
        RECT 259.775 70.035 259.915 74.620 ;
        RECT 261.155 73.435 261.295 74.815 ;
        RECT 261.095 73.115 261.355 73.435 ;
        RECT 260.635 72.775 260.895 73.095 ;
        RECT 259.715 69.715 259.975 70.035 ;
        RECT 259.255 68.695 259.515 69.015 ;
        RECT 258.335 67.335 258.595 67.655 ;
        RECT 257.415 66.995 257.675 67.315 ;
        RECT 256.025 66.460 256.305 66.830 ;
        RECT 256.035 66.315 256.295 66.460 ;
        RECT 257.415 65.975 257.675 66.295 ;
        RECT 258.335 65.975 258.595 66.295 ;
        RECT 254.475 65.440 256.015 65.810 ;
        RECT 257.475 65.275 257.615 65.975 ;
        RECT 257.415 64.955 257.675 65.275 ;
        RECT 253.275 64.275 253.535 64.595 ;
        RECT 255.565 64.420 255.845 64.790 ;
        RECT 255.635 64.255 255.775 64.420 ;
        RECT 258.395 64.255 258.535 65.975 ;
        RECT 259.315 65.275 259.455 68.695 ;
        RECT 260.695 67.995 260.835 72.775 ;
        RECT 261.095 70.055 261.355 70.375 ;
        RECT 260.635 67.675 260.895 67.995 ;
        RECT 260.175 67.225 260.435 67.315 ;
        RECT 261.155 67.225 261.295 70.055 ;
        RECT 260.175 67.085 261.295 67.225 ;
        RECT 260.175 66.995 260.435 67.085 ;
        RECT 259.715 66.830 259.975 66.975 ;
        RECT 259.705 66.460 259.985 66.830 ;
        RECT 259.255 64.955 259.515 65.275 ;
        RECT 254.655 64.110 254.915 64.255 ;
        RECT 254.645 63.740 254.925 64.110 ;
        RECT 255.575 63.935 255.835 64.255 ;
        RECT 258.335 63.935 258.595 64.255 ;
        RECT 258.785 63.740 259.065 64.110 ;
        RECT 259.775 63.915 259.915 66.460 ;
        RECT 258.855 63.575 258.995 63.740 ;
        RECT 259.715 63.595 259.975 63.915 ;
        RECT 256.955 63.255 257.215 63.575 ;
        RECT 258.795 63.255 259.055 63.575 ;
        RECT 253.735 61.555 253.995 61.875 ;
        RECT 253.795 59.835 253.935 61.555 ;
        RECT 254.475 60.000 256.015 60.370 ;
        RECT 253.735 59.515 253.995 59.835 ;
        RECT 252.815 59.235 253.075 59.495 ;
        RECT 252.815 59.175 255.775 59.235 ;
        RECT 252.875 59.095 255.775 59.175 ;
        RECT 255.635 58.815 255.775 59.095 ;
        RECT 251.895 58.495 252.155 58.815 ;
        RECT 253.275 58.495 253.535 58.815 ;
        RECT 255.575 58.495 255.835 58.815 ;
        RECT 253.335 57.115 253.475 58.495 ;
        RECT 253.275 56.795 253.535 57.115 ;
        RECT 253.275 56.115 253.535 56.435 ;
        RECT 250.975 55.095 251.635 55.155 ;
        RECT 251.035 55.015 251.635 55.095 ;
        RECT 249.595 54.075 249.855 54.395 ;
        RECT 253.335 53.715 253.475 56.115 ;
        RECT 256.495 55.775 256.755 56.095 ;
        RECT 254.475 54.560 256.015 54.930 ;
        RECT 256.555 54.395 256.695 55.775 ;
        RECT 257.015 55.415 257.155 63.255 ;
        RECT 261.615 61.875 261.755 81.275 ;
        RECT 262.075 78.535 262.215 105.415 ;
        RECT 267.135 105.395 267.275 106.775 ;
        RECT 267.595 106.075 267.735 109.225 ;
        RECT 267.995 107.455 268.255 107.775 ;
        RECT 267.535 105.755 267.795 106.075 ;
        RECT 267.075 105.075 267.335 105.395 ;
        RECT 263.395 102.695 263.655 103.015 ;
        RECT 262.935 99.975 263.195 100.295 ;
        RECT 262.475 99.635 262.735 99.955 ;
        RECT 262.535 96.070 262.675 99.635 ;
        RECT 262.995 96.555 263.135 99.975 ;
        RECT 262.935 96.235 263.195 96.555 ;
        RECT 262.465 95.700 262.745 96.070 ;
        RECT 262.465 95.020 262.745 95.390 ;
        RECT 262.535 94.175 262.675 95.020 ;
        RECT 262.935 94.195 263.195 94.515 ;
        RECT 262.475 93.855 262.735 94.175 ;
        RECT 262.475 91.815 262.735 92.135 ;
        RECT 262.535 89.755 262.675 91.815 ;
        RECT 262.995 89.755 263.135 94.195 ;
        RECT 262.475 89.435 262.735 89.755 ;
        RECT 262.935 89.435 263.195 89.755 ;
        RECT 262.475 88.755 262.735 89.075 ;
        RECT 262.535 87.035 262.675 88.755 ;
        RECT 263.455 87.115 263.595 102.695 ;
        RECT 264.315 102.015 264.575 102.335 ;
        RECT 264.375 99.955 264.515 102.015 ;
        RECT 264.315 99.635 264.575 99.955 ;
        RECT 266.615 99.295 266.875 99.615 ;
        RECT 265.695 98.615 265.955 98.935 ;
        RECT 263.845 97.740 264.125 98.110 ;
        RECT 265.755 97.915 265.895 98.615 ;
        RECT 263.915 96.895 264.055 97.740 ;
        RECT 264.775 97.595 265.035 97.915 ;
        RECT 265.695 97.595 265.955 97.915 ;
        RECT 263.855 96.575 264.115 96.895 ;
        RECT 264.835 95.195 264.975 97.595 ;
        RECT 266.675 97.235 266.815 99.295 ;
        RECT 267.135 97.575 267.275 105.075 ;
        RECT 268.055 102.675 268.195 107.455 ;
        RECT 269.895 106.075 270.035 109.225 ;
        RECT 269.835 105.755 270.095 106.075 ;
        RECT 270.295 105.075 270.555 105.395 ;
        RECT 271.675 105.075 271.935 105.395 ;
        RECT 268.915 104.735 269.175 105.055 ;
        RECT 268.975 103.355 269.115 104.735 ;
        RECT 268.915 103.035 269.175 103.355 ;
        RECT 267.995 102.355 268.255 102.675 ;
        RECT 268.455 99.295 268.715 99.615 ;
        RECT 267.075 97.255 267.335 97.575 ;
        RECT 266.615 96.915 266.875 97.235 ;
        RECT 265.235 95.895 265.495 96.215 ;
        RECT 264.775 94.875 265.035 95.195 ;
        RECT 263.845 94.340 264.125 94.710 ;
        RECT 263.915 89.270 264.055 94.340 ;
        RECT 264.315 93.175 264.575 93.495 ;
        RECT 264.375 91.455 264.515 93.175 ;
        RECT 264.315 91.135 264.575 91.455 ;
        RECT 263.845 88.900 264.125 89.270 ;
        RECT 262.475 86.715 262.735 87.035 ;
        RECT 263.455 86.975 264.515 87.115 ;
        RECT 262.465 86.180 262.745 86.550 ;
        RECT 262.935 86.375 263.195 86.695 ;
        RECT 263.855 86.375 264.115 86.695 ;
        RECT 262.535 86.015 262.675 86.180 ;
        RECT 262.995 86.015 263.135 86.375 ;
        RECT 262.475 85.695 262.735 86.015 ;
        RECT 262.935 85.695 263.195 86.015 ;
        RECT 262.535 83.975 262.675 85.695 ;
        RECT 262.475 83.655 262.735 83.975 ;
        RECT 262.015 78.275 262.275 78.535 ;
        RECT 262.015 78.215 263.595 78.275 ;
        RECT 262.075 78.135 263.595 78.215 ;
        RECT 262.015 77.195 262.275 77.515 ;
        RECT 262.075 76.155 262.215 77.195 ;
        RECT 262.935 76.855 263.195 77.175 ;
        RECT 262.015 75.835 262.275 76.155 ;
        RECT 262.995 75.135 263.135 76.855 ;
        RECT 262.935 74.815 263.195 75.135 ;
        RECT 262.475 74.135 262.735 74.455 ;
        RECT 262.935 74.135 263.195 74.455 ;
        RECT 262.015 65.975 262.275 66.295 ;
        RECT 262.075 64.595 262.215 65.975 ;
        RECT 262.015 64.275 262.275 64.595 ;
        RECT 262.535 62.215 262.675 74.135 ;
        RECT 262.475 61.895 262.735 62.215 ;
        RECT 261.555 61.785 261.815 61.875 ;
        RECT 261.155 61.645 261.815 61.785 ;
        RECT 257.875 60.875 258.135 61.195 ;
        RECT 257.935 58.475 258.075 60.875 ;
        RECT 260.635 60.535 260.895 60.855 ;
        RECT 257.875 58.155 258.135 58.475 ;
        RECT 257.415 57.815 257.675 58.135 ;
        RECT 257.475 57.115 257.615 57.815 ;
        RECT 257.415 56.795 257.675 57.115 ;
        RECT 256.955 55.095 257.215 55.415 ;
        RECT 257.875 55.095 258.135 55.415 ;
        RECT 256.495 54.075 256.755 54.395 ;
        RECT 257.015 54.055 257.155 55.095 ;
        RECT 256.955 53.735 257.215 54.055 ;
        RECT 253.275 53.395 253.535 53.715 ;
        RECT 253.335 53.115 253.475 53.395 ;
        RECT 251.955 53.035 253.475 53.115 ;
        RECT 249.135 52.715 249.395 53.035 ;
        RECT 251.895 52.975 253.475 53.035 ;
        RECT 251.895 52.715 252.155 52.975 ;
        RECT 257.935 50.995 258.075 55.095 ;
        RECT 260.695 51.675 260.835 60.535 ;
        RECT 261.155 59.235 261.295 61.645 ;
        RECT 261.555 61.555 261.815 61.645 ;
        RECT 261.155 59.095 262.675 59.235 ;
        RECT 261.155 58.815 261.295 59.095 ;
        RECT 261.095 58.495 261.355 58.815 ;
        RECT 262.535 58.135 262.675 59.095 ;
        RECT 262.995 58.815 263.135 74.135 ;
        RECT 263.455 70.035 263.595 78.135 ;
        RECT 263.395 69.715 263.655 70.035 ;
        RECT 263.395 65.975 263.655 66.295 ;
        RECT 263.455 65.275 263.595 65.975 ;
        RECT 263.395 64.955 263.655 65.275 ;
        RECT 262.935 58.495 263.195 58.815 ;
        RECT 263.395 58.495 263.655 58.815 ;
        RECT 262.475 57.815 262.735 58.135 ;
        RECT 263.455 57.115 263.595 58.495 ;
        RECT 263.395 57.025 263.655 57.115 ;
        RECT 262.995 56.885 263.655 57.025 ;
        RECT 261.095 55.775 261.355 56.095 ;
        RECT 261.155 54.055 261.295 55.775 ;
        RECT 261.555 55.095 261.815 55.415 ;
        RECT 261.615 54.055 261.755 55.095 ;
        RECT 261.095 53.735 261.355 54.055 ;
        RECT 261.555 53.735 261.815 54.055 ;
        RECT 262.015 52.605 262.275 52.695 ;
        RECT 262.995 52.605 263.135 56.885 ;
        RECT 263.395 56.795 263.655 56.885 ;
        RECT 263.395 56.115 263.655 56.435 ;
        RECT 263.455 55.155 263.595 56.115 ;
        RECT 263.915 55.755 264.055 86.375 ;
        RECT 264.375 86.015 264.515 86.975 ;
        RECT 264.315 85.695 264.575 86.015 ;
        RECT 265.295 83.635 265.435 95.895 ;
        RECT 268.515 94.425 268.655 99.295 ;
        RECT 268.975 96.895 269.115 103.035 ;
        RECT 269.835 102.695 270.095 103.015 ;
        RECT 268.915 96.575 269.175 96.895 ;
        RECT 268.915 94.425 269.175 94.515 ;
        RECT 268.515 94.285 269.175 94.425 ;
        RECT 268.915 94.195 269.175 94.285 ;
        RECT 266.155 88.755 266.415 89.075 ;
        RECT 265.685 88.475 265.965 88.590 ;
        RECT 266.215 88.475 266.355 88.755 ;
        RECT 265.685 88.335 266.355 88.475 ;
        RECT 265.685 88.220 265.965 88.335 ;
        RECT 265.695 87.735 265.955 88.055 ;
        RECT 265.755 83.635 265.895 87.735 ;
        RECT 266.215 86.015 266.355 88.335 ;
        RECT 268.455 87.735 268.715 88.055 ;
        RECT 266.615 86.375 266.875 86.695 ;
        RECT 266.155 85.695 266.415 86.015 ;
        RECT 266.155 85.015 266.415 85.335 ;
        RECT 266.215 84.315 266.355 85.015 ;
        RECT 266.155 83.995 266.415 84.315 ;
        RECT 265.235 83.315 265.495 83.635 ;
        RECT 265.695 83.315 265.955 83.635 ;
        RECT 264.775 82.295 265.035 82.615 ;
        RECT 264.315 77.875 264.575 78.195 ;
        RECT 264.375 77.030 264.515 77.875 ;
        RECT 264.305 76.660 264.585 77.030 ;
        RECT 264.315 66.995 264.575 67.315 ;
        RECT 264.375 63.575 264.515 66.995 ;
        RECT 264.315 63.255 264.575 63.575 ;
        RECT 264.315 60.535 264.575 60.855 ;
        RECT 264.375 56.435 264.515 60.535 ;
        RECT 264.315 56.115 264.575 56.435 ;
        RECT 263.855 55.435 264.115 55.755 ;
        RECT 264.835 55.155 264.975 82.295 ;
        RECT 265.755 80.915 265.895 83.315 ;
        RECT 265.695 80.595 265.955 80.915 ;
        RECT 265.235 66.315 265.495 66.635 ;
        RECT 265.295 63.575 265.435 66.315 ;
        RECT 265.235 63.255 265.495 63.575 ;
        RECT 266.675 61.195 266.815 86.375 ;
        RECT 268.515 86.015 268.655 87.735 ;
        RECT 268.455 85.695 268.715 86.015 ;
        RECT 267.535 85.015 267.795 85.335 ;
        RECT 267.995 85.015 268.255 85.335 ;
        RECT 267.075 71.755 267.335 72.075 ;
        RECT 267.135 67.315 267.275 71.755 ;
        RECT 267.075 66.995 267.335 67.315 ;
        RECT 266.615 60.875 266.875 61.195 ;
        RECT 265.695 58.495 265.955 58.815 ;
        RECT 265.755 55.755 265.895 58.495 ;
        RECT 266.155 57.815 266.415 58.135 ;
        RECT 266.615 57.815 266.875 58.135 ;
        RECT 266.215 56.435 266.355 57.815 ;
        RECT 266.675 57.115 266.815 57.815 ;
        RECT 266.615 56.795 266.875 57.115 ;
        RECT 266.155 56.115 266.415 56.435 ;
        RECT 266.605 56.260 266.885 56.630 ;
        RECT 267.595 56.435 267.735 85.015 ;
        RECT 266.615 56.115 266.875 56.260 ;
        RECT 267.535 56.115 267.795 56.435 ;
        RECT 268.055 55.755 268.195 85.015 ;
        RECT 268.455 80.255 268.715 80.575 ;
        RECT 268.515 72.075 268.655 80.255 ;
        RECT 268.455 71.755 268.715 72.075 ;
        RECT 268.975 70.795 269.115 94.195 ;
        RECT 269.375 90.455 269.635 90.775 ;
        RECT 269.435 86.015 269.575 90.455 ;
        RECT 269.895 86.015 270.035 102.695 ;
        RECT 269.375 85.695 269.635 86.015 ;
        RECT 269.835 85.695 270.095 86.015 ;
        RECT 270.355 81.255 270.495 105.075 ;
        RECT 270.755 98.955 271.015 99.275 ;
        RECT 270.815 89.415 270.955 98.955 ;
        RECT 271.215 93.855 271.475 94.175 ;
        RECT 270.755 89.095 271.015 89.415 ;
        RECT 271.275 86.015 271.415 93.855 ;
        RECT 271.215 85.695 271.475 86.015 ;
        RECT 270.295 80.935 270.555 81.255 ;
        RECT 270.295 77.875 270.555 78.195 ;
        RECT 268.515 70.655 269.115 70.795 ;
        RECT 268.515 67.655 268.655 70.655 ;
        RECT 268.915 69.715 269.175 70.035 ;
        RECT 268.455 67.335 268.715 67.655 ;
        RECT 268.515 60.855 268.655 67.335 ;
        RECT 268.975 64.595 269.115 69.715 ;
        RECT 269.835 68.695 270.095 69.015 ;
        RECT 268.915 64.275 269.175 64.595 ;
        RECT 269.895 64.255 270.035 68.695 ;
        RECT 270.355 67.315 270.495 77.875 ;
        RECT 271.735 73.435 271.875 105.075 ;
        RECT 272.195 104.375 272.335 109.225 ;
        RECT 274.495 107.095 274.635 109.225 ;
        RECT 276.275 107.115 276.535 107.435 ;
        RECT 274.435 106.775 274.695 107.095 ;
        RECT 273.105 106.240 274.645 106.610 ;
        RECT 276.335 106.075 276.475 107.115 ;
        RECT 276.795 106.075 276.935 109.225 ;
        RECT 276.275 105.755 276.535 106.075 ;
        RECT 276.735 105.755 276.995 106.075 ;
        RECT 279.095 105.395 279.235 109.225 ;
        RECT 280.875 108.135 281.135 108.455 ;
        RECT 277.195 105.075 277.455 105.395 ;
        RECT 279.035 105.075 279.295 105.395 ;
        RECT 279.495 105.075 279.755 105.395 ;
        RECT 272.135 104.055 272.395 104.375 ;
        RECT 274.895 101.675 275.155 101.995 ;
        RECT 273.105 100.800 274.645 101.170 ;
        RECT 274.955 100.295 275.095 101.675 ;
        RECT 277.255 101.510 277.395 105.075 ;
        RECT 279.555 104.795 279.695 105.075 ;
        RECT 278.635 104.655 279.695 104.795 ;
        RECT 277.655 102.015 277.915 102.335 ;
        RECT 277.185 101.140 277.465 101.510 ;
        RECT 274.895 99.975 275.155 100.295 ;
        RECT 272.595 99.295 272.855 99.615 ;
        RECT 272.655 97.915 272.795 99.295 ;
        RECT 272.595 97.595 272.855 97.915 ;
        RECT 273.105 95.360 274.645 95.730 ;
        RECT 273.105 89.920 274.645 90.290 ;
        RECT 274.955 89.755 275.095 99.975 ;
        RECT 277.715 98.935 277.855 102.015 ;
        RECT 277.655 98.615 277.915 98.935 ;
        RECT 278.105 94.340 278.385 94.710 ;
        RECT 278.115 94.195 278.375 94.340 ;
        RECT 276.735 90.455 276.995 90.775 ;
        RECT 274.895 89.435 275.155 89.755 ;
        RECT 276.795 88.735 276.935 90.455 ;
        RECT 277.655 89.095 277.915 89.415 ;
        RECT 274.895 88.415 275.155 88.735 ;
        RECT 276.735 88.415 276.995 88.735 ;
        RECT 272.135 85.015 272.395 85.335 ;
        RECT 272.195 82.955 272.335 85.015 ;
        RECT 273.105 84.480 274.645 84.850 ;
        RECT 274.435 82.975 274.695 83.295 ;
        RECT 272.135 82.635 272.395 82.955 ;
        RECT 272.595 82.295 272.855 82.615 ;
        RECT 272.655 78.195 272.795 82.295 ;
        RECT 274.495 81.595 274.635 82.975 ;
        RECT 274.955 82.615 275.095 88.415 ;
        RECT 276.735 85.015 276.995 85.335 ;
        RECT 276.795 83.830 276.935 85.015 ;
        RECT 277.715 84.315 277.855 89.095 ;
        RECT 278.175 87.035 278.315 94.195 ;
        RECT 278.635 93.835 278.775 104.655 ;
        RECT 280.415 104.395 280.675 104.715 ;
        RECT 279.495 102.355 279.755 102.675 ;
        RECT 279.555 97.235 279.695 102.355 ;
        RECT 280.475 101.995 280.615 104.395 ;
        RECT 280.935 102.675 281.075 108.135 ;
        RECT 281.395 104.715 281.535 109.225 ;
        RECT 283.175 106.775 283.435 107.095 ;
        RECT 281.795 105.075 282.055 105.395 ;
        RECT 281.335 104.395 281.595 104.715 ;
        RECT 281.855 102.755 281.995 105.075 ;
        RECT 282.255 104.735 282.515 105.055 ;
        RECT 282.315 103.355 282.455 104.735 ;
        RECT 282.255 103.035 282.515 103.355 ;
        RECT 283.235 103.015 283.375 106.775 ;
        RECT 283.695 106.075 283.835 109.225 ;
        RECT 283.635 105.755 283.895 106.075 ;
        RECT 285.015 105.305 285.275 105.395 ;
        RECT 285.015 105.165 285.675 105.305 ;
        RECT 285.015 105.075 285.275 105.165 ;
        RECT 280.875 102.355 281.135 102.675 ;
        RECT 281.395 102.615 281.995 102.755 ;
        RECT 283.175 102.695 283.435 103.015 ;
        RECT 280.415 101.675 280.675 101.995 ;
        RECT 281.395 100.715 281.535 102.615 ;
        RECT 283.635 102.015 283.895 102.335 ;
        RECT 284.095 102.015 284.355 102.335 ;
        RECT 283.695 100.830 283.835 102.015 ;
        RECT 284.155 100.995 284.295 102.015 ;
        RECT 284.155 100.855 285.215 100.995 ;
        RECT 280.935 100.575 281.535 100.715 ;
        RECT 280.415 99.635 280.675 99.955 ;
        RECT 279.955 98.790 280.215 98.935 ;
        RECT 279.945 98.420 280.225 98.790 ;
        RECT 279.495 96.915 279.755 97.235 ;
        RECT 280.015 96.895 280.155 98.420 ;
        RECT 280.475 97.915 280.615 99.635 ;
        RECT 280.415 97.595 280.675 97.915 ;
        RECT 280.935 97.315 281.075 100.575 ;
        RECT 283.625 100.460 283.905 100.830 ;
        RECT 283.175 99.975 283.435 100.295 ;
        RECT 280.475 97.175 281.075 97.315 ;
        RECT 279.955 96.575 280.215 96.895 ;
        RECT 279.495 95.895 279.755 96.215 ;
        RECT 279.035 94.195 279.295 94.515 ;
        RECT 278.575 93.515 278.835 93.835 ;
        RECT 278.115 86.715 278.375 87.035 ;
        RECT 278.115 85.695 278.375 86.015 ;
        RECT 277.655 83.995 277.915 84.315 ;
        RECT 276.725 83.460 277.005 83.830 ;
        RECT 277.195 83.655 277.455 83.975 ;
        RECT 274.895 82.295 275.155 82.615 ;
        RECT 274.435 81.275 274.695 81.595 ;
        RECT 275.355 80.255 275.615 80.575 ;
        RECT 274.895 79.575 275.155 79.895 ;
        RECT 273.105 79.040 274.645 79.410 ;
        RECT 274.955 78.875 275.095 79.575 ;
        RECT 274.895 78.555 275.155 78.875 ;
        RECT 272.595 77.875 272.855 78.195 ;
        RECT 275.415 76.155 275.555 80.255 ;
        RECT 277.255 80.235 277.395 83.655 ;
        RECT 277.195 79.915 277.455 80.235 ;
        RECT 277.255 78.535 277.395 79.915 ;
        RECT 277.195 78.215 277.455 78.535 ;
        RECT 275.805 77.340 276.085 77.710 ;
        RECT 275.355 75.835 275.615 76.155 ;
        RECT 275.355 75.155 275.615 75.475 ;
        RECT 273.105 73.600 274.645 73.970 ;
        RECT 271.675 73.115 271.935 73.435 ;
        RECT 271.735 69.550 271.875 73.115 ;
        RECT 275.415 70.035 275.555 75.155 ;
        RECT 275.875 75.135 276.015 77.340 ;
        RECT 276.275 76.855 276.535 77.175 ;
        RECT 276.335 75.135 276.475 76.855 ;
        RECT 275.815 74.815 276.075 75.135 ;
        RECT 276.275 74.990 276.535 75.135 ;
        RECT 276.265 74.620 276.545 74.990 ;
        RECT 277.195 72.775 277.455 73.095 ;
        RECT 276.735 70.395 276.995 70.715 ;
        RECT 275.355 69.715 275.615 70.035 ;
        RECT 271.665 69.180 271.945 69.550 ;
        RECT 273.105 68.160 274.645 68.530 ;
        RECT 271.215 67.335 271.475 67.655 ;
        RECT 273.055 67.565 273.315 67.655 ;
        RECT 272.655 67.425 273.315 67.565 ;
        RECT 270.295 66.995 270.555 67.315 ;
        RECT 269.835 63.935 270.095 64.255 ;
        RECT 271.275 62.555 271.415 67.335 ;
        RECT 272.655 63.915 272.795 67.425 ;
        RECT 273.055 67.335 273.315 67.425 ;
        RECT 274.895 66.655 275.155 66.975 ;
        RECT 272.595 63.595 272.855 63.915 ;
        RECT 271.215 62.235 271.475 62.555 ;
        RECT 270.755 61.215 271.015 61.535 ;
        RECT 268.455 60.535 268.715 60.855 ;
        RECT 265.695 55.435 265.955 55.755 ;
        RECT 267.995 55.435 268.255 55.755 ;
        RECT 263.455 55.015 264.975 55.155 ;
        RECT 268.455 55.095 268.715 55.415 ;
        RECT 265.695 52.715 265.955 53.035 ;
        RECT 262.015 52.465 263.135 52.605 ;
        RECT 262.015 52.375 262.275 52.465 ;
        RECT 260.635 51.355 260.895 51.675 ;
        RECT 262.995 51.335 263.135 52.465 ;
        RECT 265.235 52.375 265.495 52.695 ;
        RECT 262.935 51.015 263.195 51.335 ;
        RECT 257.875 50.675 258.135 50.995 ;
        RECT 265.295 50.655 265.435 52.375 ;
        RECT 253.735 50.335 253.995 50.655 ;
        RECT 256.955 50.335 257.215 50.655 ;
        RECT 262.935 50.335 263.195 50.655 ;
        RECT 265.235 50.335 265.495 50.655 ;
        RECT 249.135 45.915 249.395 46.235 ;
        RECT 249.195 39.095 249.335 45.915 ;
        RECT 253.795 45.555 253.935 50.335 ;
        RECT 254.475 49.120 256.015 49.490 ;
        RECT 257.015 48.275 257.155 50.335 ;
        RECT 259.715 49.655 259.975 49.975 ;
        RECT 259.775 48.955 259.915 49.655 ;
        RECT 262.995 48.955 263.135 50.335 ;
        RECT 259.715 48.635 259.975 48.955 ;
        RECT 262.935 48.635 263.195 48.955 ;
        RECT 256.955 47.955 257.215 48.275 ;
        RECT 259.255 47.955 259.515 48.275 ;
        RECT 257.875 45.915 258.135 46.235 ;
        RECT 253.735 45.235 253.995 45.555 ;
        RECT 256.955 44.215 257.215 44.535 ;
        RECT 254.475 43.680 256.015 44.050 ;
        RECT 250.975 42.515 251.235 42.835 ;
        RECT 249.135 38.775 249.395 39.095 ;
        RECT 249.195 36.715 249.335 38.775 ;
        RECT 249.135 36.395 249.395 36.715 ;
        RECT 249.195 34.675 249.335 36.395 ;
        RECT 251.035 35.355 251.175 42.515 ;
        RECT 256.495 42.235 256.755 42.495 ;
        RECT 257.015 42.235 257.155 44.215 ;
        RECT 257.935 42.495 258.075 45.915 ;
        RECT 258.335 44.895 258.595 45.215 ;
        RECT 258.395 43.175 258.535 44.895 ;
        RECT 258.335 42.855 258.595 43.175 ;
        RECT 256.495 42.175 257.155 42.235 ;
        RECT 257.875 42.175 258.135 42.495 ;
        RECT 256.555 42.095 257.155 42.175 ;
        RECT 259.315 42.155 259.455 47.955 ;
        RECT 260.635 46.935 260.895 47.255 ;
        RECT 260.695 42.835 260.835 46.935 ;
        RECT 261.095 44.895 261.355 45.215 ;
        RECT 260.635 42.515 260.895 42.835 ;
        RECT 258.335 41.835 258.595 42.155 ;
        RECT 259.255 41.835 259.515 42.155 ;
        RECT 251.435 41.495 251.695 41.815 ;
        RECT 257.415 41.495 257.675 41.815 ;
        RECT 251.495 40.455 251.635 41.495 ;
        RECT 257.475 40.455 257.615 41.495 ;
        RECT 258.395 40.455 258.535 41.835 ;
        RECT 259.315 40.795 259.455 41.835 ;
        RECT 259.255 40.475 259.515 40.795 ;
        RECT 251.435 40.135 251.695 40.455 ;
        RECT 252.355 40.135 252.615 40.455 ;
        RECT 257.415 40.135 257.675 40.455 ;
        RECT 258.335 40.135 258.595 40.455 ;
        RECT 252.415 39.095 252.555 40.135 ;
        RECT 252.355 38.775 252.615 39.095 ;
        RECT 252.415 37.055 252.555 38.775 ;
        RECT 254.475 38.240 256.015 38.610 ;
        RECT 253.735 37.755 253.995 38.075 ;
        RECT 252.355 36.735 252.615 37.055 ;
        RECT 250.975 35.035 251.235 35.355 ;
        RECT 249.135 34.355 249.395 34.675 ;
        RECT 251.435 33.335 251.695 33.655 ;
        RECT 251.495 31.955 251.635 33.335 ;
        RECT 251.435 31.635 251.695 31.955 ;
        RECT 253.795 31.615 253.935 37.755 ;
        RECT 255.115 36.735 255.375 37.055 ;
        RECT 255.175 35.355 255.315 36.735 ;
        RECT 258.395 36.375 258.535 40.135 ;
        RECT 261.155 37.395 261.295 44.895 ;
        RECT 265.295 44.875 265.435 50.335 ;
        RECT 265.755 47.595 265.895 52.715 ;
        RECT 268.515 51.335 268.655 55.095 ;
        RECT 270.815 54.055 270.955 61.215 ;
        RECT 272.135 57.815 272.395 58.135 ;
        RECT 272.195 55.415 272.335 57.815 ;
        RECT 272.655 56.435 272.795 63.595 ;
        RECT 273.105 62.720 274.645 63.090 ;
        RECT 274.955 62.555 275.095 66.655 ;
        RECT 275.415 62.555 275.555 69.715 ;
        RECT 276.795 67.315 276.935 70.395 ;
        RECT 277.255 70.230 277.395 72.775 ;
        RECT 278.175 72.755 278.315 85.695 ;
        RECT 279.095 85.335 279.235 94.195 ;
        RECT 279.555 92.475 279.695 95.895 ;
        RECT 280.475 95.275 280.615 97.175 ;
        RECT 282.255 96.915 282.515 97.235 ;
        RECT 280.875 96.750 281.135 96.895 ;
        RECT 280.865 96.380 281.145 96.750 ;
        RECT 280.475 95.135 281.075 95.275 ;
        RECT 280.415 94.425 280.675 94.515 ;
        RECT 280.015 94.285 280.675 94.425 ;
        RECT 279.495 92.155 279.755 92.475 ;
        RECT 279.555 91.115 279.695 92.155 ;
        RECT 279.495 90.795 279.755 91.115 ;
        RECT 279.035 85.015 279.295 85.335 ;
        RECT 278.575 80.255 278.835 80.575 ;
        RECT 278.635 76.155 278.775 80.255 ;
        RECT 278.575 75.835 278.835 76.155 ;
        RECT 278.115 72.435 278.375 72.755 ;
        RECT 279.495 72.435 279.755 72.755 ;
        RECT 277.185 69.860 277.465 70.230 ;
        RECT 278.175 67.655 278.315 72.435 ;
        RECT 278.575 72.095 278.835 72.415 ;
        RECT 278.635 69.695 278.775 72.095 ;
        RECT 279.555 69.695 279.695 72.435 ;
        RECT 280.015 70.715 280.155 94.285 ;
        RECT 280.415 94.195 280.675 94.285 ;
        RECT 280.935 76.155 281.075 95.135 ;
        RECT 282.315 94.175 282.455 96.915 ;
        RECT 282.715 95.895 282.975 96.215 ;
        RECT 282.775 95.195 282.915 95.895 ;
        RECT 283.235 95.195 283.375 99.975 ;
        RECT 283.625 97.060 283.905 97.430 ;
        RECT 283.635 96.915 283.895 97.060 ;
        RECT 284.095 96.915 284.355 97.235 ;
        RECT 283.635 96.235 283.895 96.555 ;
        RECT 283.695 95.195 283.835 96.235 ;
        RECT 284.155 96.215 284.295 96.915 ;
        RECT 284.095 95.895 284.355 96.215 ;
        RECT 282.715 94.875 282.975 95.195 ;
        RECT 283.175 94.875 283.435 95.195 ;
        RECT 283.635 94.875 283.895 95.195 ;
        RECT 282.255 93.855 282.515 94.175 ;
        RECT 281.795 93.515 282.055 93.835 ;
        RECT 281.855 91.795 281.995 93.515 ;
        RECT 281.795 91.475 282.055 91.795 ;
        RECT 282.715 91.135 282.975 91.455 ;
        RECT 282.775 89.755 282.915 91.135 ;
        RECT 285.075 91.115 285.215 100.855 ;
        RECT 285.015 90.795 285.275 91.115 ;
        RECT 283.175 90.455 283.435 90.775 ;
        RECT 284.555 90.455 284.815 90.775 ;
        RECT 282.715 89.435 282.975 89.755 ;
        RECT 283.235 89.415 283.375 90.455 ;
        RECT 283.175 89.095 283.435 89.415 ;
        RECT 282.715 88.075 282.975 88.395 ;
        RECT 282.775 87.035 282.915 88.075 ;
        RECT 282.715 86.715 282.975 87.035 ;
        RECT 284.615 86.355 284.755 90.455 ;
        RECT 285.075 88.055 285.215 90.795 ;
        RECT 285.015 87.735 285.275 88.055 ;
        RECT 285.015 86.715 285.275 87.035 ;
        RECT 284.555 86.035 284.815 86.355 ;
        RECT 282.255 83.655 282.515 83.975 ;
        RECT 281.785 82.780 282.065 83.150 ;
        RECT 281.795 82.635 282.055 82.780 ;
        RECT 280.875 75.835 281.135 76.155 ;
        RECT 281.855 75.475 281.995 82.635 ;
        RECT 282.315 78.535 282.455 83.655 ;
        RECT 285.075 80.915 285.215 86.715 ;
        RECT 285.015 80.595 285.275 80.915 ;
        RECT 284.555 79.915 284.815 80.235 ;
        RECT 284.615 78.875 284.755 79.915 ;
        RECT 284.555 78.555 284.815 78.875 ;
        RECT 285.075 78.535 285.215 80.595 ;
        RECT 282.255 78.215 282.515 78.535 ;
        RECT 285.015 78.215 285.275 78.535 ;
        RECT 285.535 77.595 285.675 105.165 ;
        RECT 285.995 104.375 286.135 109.225 ;
        RECT 288.295 107.775 288.435 109.225 ;
        RECT 288.235 107.455 288.495 107.775 ;
        RECT 290.075 107.115 290.335 107.435 ;
        RECT 288.235 105.075 288.495 105.395 ;
        RECT 289.155 105.075 289.415 105.395 ;
        RECT 285.935 104.055 286.195 104.375 ;
        RECT 288.295 102.675 288.435 105.075 ;
        RECT 288.235 102.355 288.495 102.675 ;
        RECT 286.395 101.675 286.655 101.995 ;
        RECT 287.775 101.675 288.035 101.995 ;
        RECT 286.455 98.935 286.595 101.675 ;
        RECT 286.855 101.335 287.115 101.655 ;
        RECT 286.395 98.615 286.655 98.935 ;
        RECT 285.925 97.060 286.205 97.430 ;
        RECT 285.935 96.915 286.195 97.060 ;
        RECT 286.915 89.755 287.055 101.335 ;
        RECT 287.835 100.830 287.975 101.675 ;
        RECT 288.295 101.655 288.435 102.355 ;
        RECT 288.235 101.335 288.495 101.655 ;
        RECT 289.215 100.995 289.355 105.075 ;
        RECT 289.615 104.055 289.875 104.375 ;
        RECT 289.675 103.355 289.815 104.055 ;
        RECT 290.135 103.355 290.275 107.115 ;
        RECT 290.595 106.075 290.735 109.225 ;
        RECT 292.895 107.095 293.035 109.225 ;
        RECT 292.835 106.775 293.095 107.095 ;
        RECT 290.535 105.755 290.795 106.075 ;
        RECT 294.215 105.075 294.475 105.395 ;
        RECT 291.735 103.520 293.275 103.890 ;
        RECT 289.615 103.035 289.875 103.355 ;
        RECT 290.075 103.035 290.335 103.355 ;
        RECT 289.215 100.855 289.815 100.995 ;
        RECT 287.765 100.460 288.045 100.830 ;
        RECT 287.775 100.315 288.035 100.460 ;
        RECT 289.145 99.780 289.425 100.150 ;
        RECT 288.235 98.615 288.495 98.935 ;
        RECT 288.295 96.895 288.435 98.615 ;
        RECT 288.235 96.575 288.495 96.895 ;
        RECT 289.215 96.555 289.355 99.780 ;
        RECT 289.675 97.915 289.815 100.855 ;
        RECT 289.615 97.595 289.875 97.915 ;
        RECT 289.155 96.235 289.415 96.555 ;
        RECT 289.675 95.195 289.815 97.595 ;
        RECT 290.135 96.895 290.275 103.035 ;
        RECT 290.535 99.975 290.795 100.295 ;
        RECT 290.075 96.575 290.335 96.895 ;
        RECT 290.595 95.195 290.735 99.975 ;
        RECT 293.755 98.615 294.015 98.935 ;
        RECT 291.735 98.080 293.275 98.450 ;
        RECT 292.375 97.595 292.635 97.915 ;
        RECT 290.995 96.235 291.255 96.555 ;
        RECT 289.615 94.875 289.875 95.195 ;
        RECT 290.535 94.875 290.795 95.195 ;
        RECT 289.155 91.475 289.415 91.795 ;
        RECT 286.855 89.435 287.115 89.755 ;
        RECT 285.925 88.900 286.205 89.270 ;
        RECT 285.935 88.755 286.195 88.900 ;
        RECT 286.395 88.415 286.655 88.735 ;
        RECT 286.455 86.355 286.595 88.415 ;
        RECT 286.915 87.035 287.055 89.435 ;
        RECT 288.235 88.755 288.495 89.075 ;
        RECT 288.295 87.035 288.435 88.755 ;
        RECT 289.215 88.735 289.355 91.475 ;
        RECT 291.055 91.455 291.195 96.235 ;
        RECT 292.435 96.215 292.575 97.595 ;
        RECT 292.835 96.915 293.095 97.235 ;
        RECT 291.915 95.895 292.175 96.215 ;
        RECT 292.375 95.895 292.635 96.215 ;
        RECT 291.975 95.195 292.115 95.895 ;
        RECT 291.915 94.875 292.175 95.195 ;
        RECT 292.435 93.495 292.575 95.895 ;
        RECT 292.895 94.175 293.035 96.915 ;
        RECT 293.815 96.895 293.955 98.615 ;
        RECT 293.755 96.575 294.015 96.895 ;
        RECT 292.835 93.855 293.095 94.175 ;
        RECT 293.815 93.495 293.955 96.575 ;
        RECT 292.375 93.175 292.635 93.495 ;
        RECT 293.755 93.175 294.015 93.495 ;
        RECT 291.735 92.640 293.275 93.010 ;
        RECT 290.995 91.135 291.255 91.455 ;
        RECT 291.905 90.940 292.185 91.310 ;
        RECT 291.915 90.795 292.175 90.940 ;
        RECT 290.075 90.455 290.335 90.775 ;
        RECT 290.135 89.415 290.275 90.455 ;
        RECT 290.075 89.095 290.335 89.415 ;
        RECT 289.155 88.415 289.415 88.735 ;
        RECT 293.755 87.735 294.015 88.055 ;
        RECT 291.735 87.200 293.275 87.570 ;
        RECT 293.815 87.035 293.955 87.735 ;
        RECT 286.855 86.715 287.115 87.035 ;
        RECT 288.235 86.715 288.495 87.035 ;
        RECT 293.755 86.715 294.015 87.035 ;
        RECT 286.395 86.035 286.655 86.355 ;
        RECT 293.295 85.695 293.555 86.015 ;
        RECT 294.275 85.755 294.415 105.075 ;
        RECT 295.195 103.355 295.335 109.225 ;
        RECT 297.495 106.075 297.635 109.225 ;
        RECT 297.895 108.135 298.155 108.455 ;
        RECT 297.435 105.755 297.695 106.075 ;
        RECT 296.515 104.735 296.775 105.055 ;
        RECT 295.135 103.035 295.395 103.355 ;
        RECT 295.135 101.675 295.395 101.995 ;
        RECT 295.195 100.295 295.335 101.675 ;
        RECT 295.135 99.975 295.395 100.295 ;
        RECT 295.195 94.855 295.335 99.975 ;
        RECT 295.135 94.535 295.395 94.855 ;
        RECT 295.195 89.415 295.335 94.535 ;
        RECT 295.595 91.475 295.855 91.795 ;
        RECT 295.135 89.095 295.395 89.415 ;
        RECT 294.675 86.375 294.935 86.695 ;
        RECT 292.375 85.355 292.635 85.675 ;
        RECT 292.435 83.975 292.575 85.355 ;
        RECT 293.355 84.315 293.495 85.695 ;
        RECT 293.815 85.615 294.415 85.755 ;
        RECT 293.295 83.995 293.555 84.315 ;
        RECT 292.375 83.655 292.635 83.975 ;
        RECT 288.235 83.315 288.495 83.635 ;
        RECT 286.855 82.295 287.115 82.615 ;
        RECT 286.915 80.915 287.055 82.295 ;
        RECT 288.295 81.595 288.435 83.315 ;
        RECT 291.735 81.760 293.275 82.130 ;
        RECT 288.235 81.275 288.495 81.595 ;
        RECT 293.815 81.110 293.955 85.615 ;
        RECT 294.735 83.715 294.875 86.375 ;
        RECT 295.195 85.675 295.335 89.095 ;
        RECT 295.655 86.355 295.795 91.475 ;
        RECT 295.595 86.035 295.855 86.355 ;
        RECT 295.135 85.355 295.395 85.675 ;
        RECT 296.055 85.355 296.315 85.675 ;
        RECT 296.115 83.975 296.255 85.355 ;
        RECT 294.735 83.575 295.335 83.715 ;
        RECT 296.055 83.655 296.315 83.975 ;
        RECT 294.675 82.975 294.935 83.295 ;
        RECT 286.855 80.595 287.115 80.915 ;
        RECT 289.145 80.740 289.425 81.110 ;
        RECT 285.935 77.875 286.195 78.195 ;
        RECT 283.695 77.455 285.675 77.595 ;
        RECT 281.795 75.155 282.055 75.475 ;
        RECT 280.415 72.095 280.675 72.415 ;
        RECT 279.955 70.395 280.215 70.715 ;
        RECT 278.575 69.375 278.835 69.695 ;
        RECT 279.495 69.375 279.755 69.695 ;
        RECT 278.115 67.335 278.375 67.655 ;
        RECT 276.735 66.995 276.995 67.315 ;
        RECT 277.655 66.655 277.915 66.975 ;
        RECT 277.715 64.595 277.855 66.655 ;
        RECT 277.655 64.275 277.915 64.595 ;
        RECT 274.895 62.235 275.155 62.555 ;
        RECT 275.355 62.235 275.615 62.555 ;
        RECT 275.415 61.535 275.555 62.235 ;
        RECT 278.635 61.875 278.775 69.375 ;
        RECT 279.555 66.295 279.695 69.375 ;
        RECT 280.475 66.975 280.615 72.095 ;
        RECT 281.335 68.695 281.595 69.015 ;
        RECT 281.395 67.655 281.535 68.695 ;
        RECT 281.335 67.335 281.595 67.655 ;
        RECT 280.415 66.655 280.675 66.975 ;
        RECT 279.495 65.975 279.755 66.295 ;
        RECT 279.555 61.875 279.695 65.975 ;
        RECT 283.695 64.255 283.835 77.455 ;
        RECT 285.015 74.815 285.275 75.135 ;
        RECT 284.095 74.475 284.355 74.795 ;
        RECT 284.155 64.935 284.295 74.475 ;
        RECT 284.555 74.135 284.815 74.455 ;
        RECT 284.615 73.435 284.755 74.135 ;
        RECT 284.555 73.115 284.815 73.435 ;
        RECT 285.075 70.715 285.215 74.815 ;
        RECT 285.475 72.775 285.735 73.095 ;
        RECT 285.015 70.395 285.275 70.715 ;
        RECT 284.545 69.860 284.825 70.230 ;
        RECT 284.615 69.695 284.755 69.860 ;
        RECT 284.555 69.375 284.815 69.695 ;
        RECT 284.615 68.075 284.755 69.375 ;
        RECT 284.615 67.995 285.215 68.075 ;
        RECT 284.615 67.935 285.275 67.995 ;
        RECT 285.015 67.675 285.275 67.935 ;
        RECT 284.095 64.615 284.355 64.935 ;
        RECT 285.535 64.255 285.675 72.775 ;
        RECT 285.995 72.755 286.135 77.875 ;
        RECT 288.695 74.135 288.955 74.455 ;
        RECT 286.395 73.115 286.655 73.435 ;
        RECT 285.935 72.435 286.195 72.755 ;
        RECT 283.635 63.935 283.895 64.255 ;
        RECT 285.015 63.935 285.275 64.255 ;
        RECT 285.475 63.935 285.735 64.255 ;
        RECT 284.555 63.595 284.815 63.915 ;
        RECT 283.175 63.255 283.435 63.575 ;
        RECT 284.095 63.255 284.355 63.575 ;
        RECT 283.235 61.875 283.375 63.255 ;
        RECT 283.635 61.955 283.895 62.215 ;
        RECT 284.155 61.955 284.295 63.255 ;
        RECT 283.635 61.895 284.295 61.955 ;
        RECT 278.575 61.555 278.835 61.875 ;
        RECT 279.495 61.555 279.755 61.875 ;
        RECT 283.175 61.555 283.435 61.875 ;
        RECT 283.695 61.815 284.295 61.895 ;
        RECT 275.355 61.215 275.615 61.535 ;
        RECT 282.255 60.535 282.515 60.855 ;
        RECT 282.315 59.835 282.455 60.535 ;
        RECT 282.255 59.515 282.515 59.835 ;
        RECT 280.415 58.495 280.675 58.815 ;
        RECT 273.105 57.280 274.645 57.650 ;
        RECT 280.475 57.115 280.615 58.495 ;
        RECT 280.415 56.795 280.675 57.115 ;
        RECT 272.595 56.115 272.855 56.435 ;
        RECT 283.235 56.095 283.375 61.555 ;
        RECT 284.615 61.535 284.755 63.595 ;
        RECT 285.075 62.555 285.215 63.935 ;
        RECT 285.015 62.235 285.275 62.555 ;
        RECT 284.095 61.215 284.355 61.535 ;
        RECT 284.555 61.390 284.815 61.535 ;
        RECT 284.155 60.765 284.295 61.215 ;
        RECT 284.545 61.020 284.825 61.390 ;
        RECT 285.075 60.765 285.215 62.235 ;
        RECT 284.155 60.625 285.215 60.765 ;
        RECT 283.175 55.775 283.435 56.095 ;
        RECT 272.135 55.095 272.395 55.415 ;
        RECT 270.755 53.735 271.015 54.055 ;
        RECT 268.915 51.355 269.175 51.675 ;
        RECT 268.455 51.015 268.715 51.335 ;
        RECT 266.155 48.295 266.415 48.615 ;
        RECT 265.695 47.275 265.955 47.595 ;
        RECT 265.235 44.555 265.495 44.875 ;
        RECT 265.695 44.215 265.955 44.535 ;
        RECT 265.755 42.835 265.895 44.215 ;
        RECT 265.695 42.515 265.955 42.835 ;
        RECT 266.215 42.235 266.355 48.295 ;
        RECT 266.615 47.275 266.875 47.595 ;
        RECT 265.755 42.155 266.355 42.235 ;
        RECT 265.695 42.095 266.355 42.155 ;
        RECT 266.675 43.085 266.815 47.275 ;
        RECT 268.455 46.935 268.715 47.255 ;
        RECT 268.515 45.555 268.655 46.935 ;
        RECT 268.975 45.895 269.115 51.355 ;
        RECT 269.375 51.015 269.635 51.335 ;
        RECT 269.435 48.615 269.575 51.015 ;
        RECT 270.815 50.655 270.955 53.735 ;
        RECT 272.195 53.715 272.335 55.095 ;
        RECT 272.135 53.395 272.395 53.715 ;
        RECT 281.325 53.540 281.605 53.910 ;
        RECT 281.395 53.375 281.535 53.540 ;
        RECT 285.995 53.375 286.135 72.435 ;
        RECT 286.455 63.915 286.595 73.115 ;
        RECT 288.235 70.395 288.495 70.715 ;
        RECT 288.295 69.015 288.435 70.395 ;
        RECT 288.755 69.695 288.895 74.135 ;
        RECT 288.695 69.375 288.955 69.695 ;
        RECT 288.235 68.695 288.495 69.015 ;
        RECT 286.395 63.595 286.655 63.915 ;
        RECT 288.295 63.575 288.435 68.695 ;
        RECT 288.235 63.255 288.495 63.575 ;
        RECT 288.295 61.875 288.435 63.255 ;
        RECT 289.215 62.215 289.355 80.740 ;
        RECT 290.075 80.595 290.335 80.915 ;
        RECT 293.745 80.740 294.025 81.110 ;
        RECT 290.135 70.035 290.275 80.595 ;
        RECT 293.755 80.255 294.015 80.575 ;
        RECT 292.835 79.915 293.095 80.235 ;
        RECT 290.995 77.875 291.255 78.195 ;
        RECT 291.055 77.595 291.195 77.875 ;
        RECT 292.895 77.595 293.035 79.915 ;
        RECT 291.055 77.455 293.035 77.595 ;
        RECT 291.055 74.795 291.195 77.455 ;
        RECT 291.735 76.320 293.275 76.690 ;
        RECT 290.995 74.475 291.255 74.795 ;
        RECT 290.075 69.715 290.335 70.035 ;
        RECT 290.135 66.495 290.275 69.715 ;
        RECT 291.055 67.655 291.195 74.475 ;
        RECT 293.815 73.435 293.955 80.255 ;
        RECT 294.735 78.195 294.875 82.975 ;
        RECT 295.195 78.875 295.335 83.575 ;
        RECT 296.055 80.935 296.315 81.255 ;
        RECT 295.135 78.555 295.395 78.875 ;
        RECT 294.675 77.875 294.935 78.195 ;
        RECT 294.215 74.135 294.475 74.455 ;
        RECT 294.675 74.135 294.935 74.455 ;
        RECT 293.755 73.115 294.015 73.435 ;
        RECT 294.275 72.415 294.415 74.135 ;
        RECT 294.215 72.095 294.475 72.415 ;
        RECT 291.735 70.880 293.275 71.250 ;
        RECT 294.275 70.035 294.415 72.095 ;
        RECT 294.735 72.075 294.875 74.135 ;
        RECT 296.115 73.095 296.255 80.935 ;
        RECT 296.055 72.775 296.315 73.095 ;
        RECT 294.675 71.755 294.935 72.075 ;
        RECT 294.215 69.715 294.475 70.035 ;
        RECT 290.995 67.335 291.255 67.655 ;
        RECT 294.275 67.315 294.415 69.715 ;
        RECT 293.755 66.995 294.015 67.315 ;
        RECT 294.215 66.995 294.475 67.315 ;
        RECT 290.135 66.355 291.195 66.495 ;
        RECT 291.055 64.595 291.195 66.355 ;
        RECT 291.735 65.440 293.275 65.810 ;
        RECT 293.815 65.275 293.955 66.995 ;
        RECT 296.575 66.495 296.715 104.735 ;
        RECT 296.975 99.295 297.235 99.615 ;
        RECT 297.035 97.235 297.175 99.295 ;
        RECT 297.955 97.235 298.095 108.135 ;
        RECT 299.795 106.075 299.935 109.225 ;
        RECT 300.195 107.455 300.455 107.775 ;
        RECT 300.255 106.075 300.395 107.455 ;
        RECT 302.095 106.075 302.235 109.225 ;
        RECT 302.495 106.775 302.755 107.095 ;
        RECT 299.735 105.755 299.995 106.075 ;
        RECT 300.195 105.755 300.455 106.075 ;
        RECT 302.035 105.755 302.295 106.075 ;
        RECT 301.115 105.075 301.375 105.395 ;
        RECT 300.195 104.735 300.455 105.055 ;
        RECT 299.275 98.955 299.535 99.275 ;
        RECT 296.975 96.915 297.235 97.235 ;
        RECT 297.895 96.915 298.155 97.235 ;
        RECT 296.975 93.175 297.235 93.495 ;
        RECT 297.035 86.015 297.175 93.175 ;
        RECT 297.955 91.795 298.095 96.915 ;
        RECT 299.335 96.750 299.475 98.955 ;
        RECT 299.265 96.380 299.545 96.750 ;
        RECT 297.895 91.475 298.155 91.795 ;
        RECT 299.335 87.035 299.475 96.380 ;
        RECT 300.255 88.055 300.395 104.735 ;
        RECT 300.655 94.195 300.915 94.515 ;
        RECT 300.715 89.075 300.855 94.195 ;
        RECT 300.655 88.755 300.915 89.075 ;
        RECT 300.195 87.735 300.455 88.055 ;
        RECT 299.275 86.715 299.535 87.035 ;
        RECT 296.975 85.695 297.235 86.015 ;
        RECT 297.435 85.015 297.695 85.335 ;
        RECT 297.495 83.975 297.635 85.015 ;
        RECT 300.715 84.315 300.855 88.755 ;
        RECT 300.655 83.995 300.915 84.315 ;
        RECT 297.435 83.655 297.695 83.975 ;
        RECT 301.175 83.715 301.315 105.075 ;
        RECT 302.555 104.375 302.695 106.775 ;
        RECT 302.955 104.395 303.215 104.715 ;
        RECT 302.495 104.055 302.755 104.375 ;
        RECT 302.035 101.675 302.295 101.995 ;
        RECT 302.495 101.675 302.755 101.995 ;
        RECT 302.095 100.995 302.235 101.675 ;
        RECT 301.635 100.855 302.235 100.995 ;
        RECT 301.635 97.915 301.775 100.855 ;
        RECT 302.035 98.615 302.295 98.935 ;
        RECT 301.575 97.595 301.835 97.915 ;
        RECT 302.095 96.895 302.235 98.615 ;
        RECT 302.035 96.575 302.295 96.895 ;
        RECT 302.035 95.895 302.295 96.215 ;
        RECT 302.095 95.195 302.235 95.895 ;
        RECT 302.035 94.875 302.295 95.195 ;
        RECT 302.035 93.855 302.295 94.175 ;
        RECT 301.575 91.815 301.835 92.135 ;
        RECT 301.635 89.415 301.775 91.815 ;
        RECT 301.575 89.095 301.835 89.415 ;
        RECT 302.095 87.035 302.235 93.855 ;
        RECT 302.555 91.455 302.695 101.675 ;
        RECT 303.015 93.495 303.155 104.395 ;
        RECT 303.415 102.015 303.675 102.335 ;
        RECT 303.475 94.855 303.615 102.015 ;
        RECT 303.875 101.335 304.135 101.655 ;
        RECT 303.935 100.635 304.075 101.335 ;
        RECT 303.875 100.315 304.135 100.635 ;
        RECT 303.865 99.100 304.145 99.470 ;
        RECT 303.935 95.195 304.075 99.100 ;
        RECT 304.395 98.935 304.535 109.225 ;
        RECT 304.795 105.075 305.055 105.395 ;
        RECT 304.335 98.615 304.595 98.935 ;
        RECT 303.875 94.875 304.135 95.195 ;
        RECT 303.415 94.535 303.675 94.855 ;
        RECT 302.955 93.175 303.215 93.495 ;
        RECT 302.495 91.135 302.755 91.455 ;
        RECT 302.555 88.735 302.695 91.135 ;
        RECT 303.935 89.755 304.075 94.875 ;
        RECT 303.875 89.435 304.135 89.755 ;
        RECT 302.495 88.415 302.755 88.735 ;
        RECT 302.035 86.715 302.295 87.035 ;
        RECT 303.935 85.675 304.075 89.435 ;
        RECT 303.875 85.355 304.135 85.675 ;
        RECT 300.715 83.575 301.315 83.715 ;
        RECT 303.415 83.655 303.675 83.975 ;
        RECT 296.975 82.975 297.235 83.295 ;
        RECT 298.355 82.975 298.615 83.295 ;
        RECT 297.035 80.575 297.175 82.975 ;
        RECT 298.415 80.915 298.555 82.975 ;
        RECT 298.355 80.595 298.615 80.915 ;
        RECT 296.975 80.255 297.235 80.575 ;
        RECT 297.895 77.535 298.155 77.855 ;
        RECT 297.955 74.795 298.095 77.535 ;
        RECT 298.415 75.475 298.555 80.595 ;
        RECT 299.735 75.495 299.995 75.815 ;
        RECT 298.355 75.155 298.615 75.475 ;
        RECT 299.795 75.135 299.935 75.495 ;
        RECT 299.735 74.815 299.995 75.135 ;
        RECT 297.895 74.475 298.155 74.795 ;
        RECT 297.435 74.135 297.695 74.455 ;
        RECT 298.355 74.135 298.615 74.455 ;
        RECT 297.495 69.015 297.635 74.135 ;
        RECT 298.415 70.035 298.555 74.135 ;
        RECT 298.355 69.715 298.615 70.035 ;
        RECT 297.435 68.695 297.695 69.015 ;
        RECT 296.115 66.355 296.715 66.495 ;
        RECT 293.755 64.955 294.015 65.275 ;
        RECT 296.115 64.790 296.255 66.355 ;
        RECT 290.995 64.275 291.255 64.595 ;
        RECT 296.045 64.420 296.325 64.790 ;
        RECT 296.115 62.555 296.255 64.420 ;
        RECT 296.515 64.275 296.775 64.595 ;
        RECT 296.055 62.235 296.315 62.555 ;
        RECT 289.155 61.895 289.415 62.215 ;
        RECT 288.235 61.555 288.495 61.875 ;
        RECT 289.215 59.835 289.355 61.895 ;
        RECT 293.755 61.555 294.015 61.875 ;
        RECT 290.075 60.535 290.335 60.855 ;
        RECT 289.155 59.515 289.415 59.835 ;
        RECT 290.135 58.815 290.275 60.535 ;
        RECT 291.735 60.000 293.275 60.370 ;
        RECT 293.815 59.835 293.955 61.555 ;
        RECT 294.215 61.215 294.475 61.535 ;
        RECT 293.755 59.515 294.015 59.835 ;
        RECT 290.075 58.495 290.335 58.815 ;
        RECT 288.695 58.155 288.955 58.475 ;
        RECT 288.235 56.795 288.495 57.115 ;
        RECT 288.295 53.375 288.435 56.795 ;
        RECT 288.755 56.775 288.895 58.155 ;
        RECT 289.615 57.815 289.875 58.135 ;
        RECT 289.675 56.775 289.815 57.815 ;
        RECT 288.695 56.455 288.955 56.775 ;
        RECT 289.615 56.455 289.875 56.775 ;
        RECT 288.755 56.095 288.895 56.455 ;
        RECT 294.275 56.095 294.415 61.215 ;
        RECT 296.115 58.815 296.255 62.235 ;
        RECT 296.575 60.855 296.715 64.275 ;
        RECT 296.515 60.535 296.775 60.855 ;
        RECT 296.575 59.155 296.715 60.535 ;
        RECT 296.515 58.835 296.775 59.155 ;
        RECT 296.055 58.495 296.315 58.815 ;
        RECT 297.495 58.475 297.635 68.695 ;
        RECT 297.885 67.140 298.165 67.510 ;
        RECT 297.955 66.495 298.095 67.140 ;
        RECT 300.715 66.495 300.855 83.575 ;
        RECT 301.115 82.975 301.375 83.295 ;
        RECT 301.175 81.595 301.315 82.975 ;
        RECT 301.575 82.295 301.835 82.615 ;
        RECT 301.115 81.275 301.375 81.595 ;
        RECT 301.115 79.575 301.375 79.895 ;
        RECT 301.175 70.715 301.315 79.575 ;
        RECT 301.635 78.390 301.775 82.295 ;
        RECT 303.475 80.235 303.615 83.655 ;
        RECT 303.415 79.915 303.675 80.235 ;
        RECT 303.475 78.535 303.615 79.915 ;
        RECT 301.565 78.020 301.845 78.390 ;
        RECT 303.415 78.215 303.675 78.535 ;
        RECT 301.635 75.135 301.775 78.020 ;
        RECT 301.575 74.815 301.835 75.135 ;
        RECT 303.475 73.095 303.615 78.215 ;
        RECT 303.415 72.775 303.675 73.095 ;
        RECT 301.115 70.395 301.375 70.715 ;
        RECT 303.475 69.695 303.615 72.775 ;
        RECT 303.935 70.375 304.075 85.355 ;
        RECT 304.855 81.595 304.995 105.075 ;
        RECT 305.255 99.635 305.515 99.955 ;
        RECT 304.795 81.275 305.055 81.595 ;
        RECT 305.315 80.995 305.455 99.635 ;
        RECT 305.715 99.295 305.975 99.615 ;
        RECT 305.775 85.335 305.915 99.295 ;
        RECT 306.695 97.915 306.835 109.225 ;
        RECT 308.475 105.075 308.735 105.395 ;
        RECT 307.555 101.675 307.815 101.995 ;
        RECT 307.615 100.995 307.755 101.675 ;
        RECT 307.155 100.855 307.755 100.995 ;
        RECT 306.635 97.595 306.895 97.915 ;
        RECT 305.715 85.015 305.975 85.335 ;
        RECT 306.175 85.015 306.435 85.335 ;
        RECT 304.855 80.855 305.455 80.995 ;
        RECT 304.335 80.255 304.595 80.575 ;
        RECT 304.395 73.435 304.535 80.255 ;
        RECT 304.855 74.795 304.995 80.855 ;
        RECT 305.255 80.255 305.515 80.575 ;
        RECT 305.315 76.155 305.455 80.255 ;
        RECT 305.775 77.855 305.915 85.015 ;
        RECT 305.715 77.535 305.975 77.855 ;
        RECT 305.255 75.835 305.515 76.155 ;
        RECT 304.795 74.475 305.055 74.795 ;
        RECT 304.335 73.115 304.595 73.435 ;
        RECT 304.855 70.715 304.995 74.475 ;
        RECT 304.795 70.395 305.055 70.715 ;
        RECT 303.875 70.055 304.135 70.375 ;
        RECT 303.415 69.375 303.675 69.695 ;
        RECT 303.475 67.655 303.615 69.375 ;
        RECT 303.935 67.995 304.075 70.055 ;
        RECT 304.335 69.375 304.595 69.695 ;
        RECT 303.875 67.675 304.135 67.995 ;
        RECT 303.415 67.335 303.675 67.655 ;
        RECT 297.955 66.355 300.855 66.495 ;
        RECT 298.415 63.575 298.555 66.355 ;
        RECT 303.875 65.975 304.135 66.295 ;
        RECT 303.935 64.255 304.075 65.975 ;
        RECT 303.875 63.935 304.135 64.255 ;
        RECT 298.355 63.255 298.615 63.575 ;
        RECT 299.275 63.255 299.535 63.575 ;
        RECT 297.435 58.155 297.695 58.475 ;
        RECT 298.415 57.115 298.555 63.255 ;
        RECT 299.335 58.815 299.475 63.255 ;
        RECT 299.275 58.495 299.535 58.815 ;
        RECT 298.815 57.815 299.075 58.135 ;
        RECT 298.355 56.795 298.615 57.115 ;
        RECT 298.875 56.775 299.015 57.815 ;
        RECT 298.815 56.455 299.075 56.775 ;
        RECT 295.595 56.115 295.855 56.435 ;
        RECT 288.695 55.775 288.955 56.095 ;
        RECT 294.215 55.775 294.475 56.095 ;
        RECT 294.215 55.095 294.475 55.415 ;
        RECT 291.735 54.560 293.275 54.930 ;
        RECT 294.275 53.375 294.415 55.095 ;
        RECT 274.895 53.055 275.155 53.375 ;
        RECT 278.115 53.055 278.375 53.375 ;
        RECT 281.335 53.055 281.595 53.375 ;
        RECT 285.935 53.055 286.195 53.375 ;
        RECT 288.235 53.055 288.495 53.375 ;
        RECT 293.755 53.055 294.015 53.375 ;
        RECT 294.215 53.055 294.475 53.375 ;
        RECT 273.105 51.840 274.645 52.210 ;
        RECT 270.755 50.335 271.015 50.655 ;
        RECT 273.515 49.995 273.775 50.315 ;
        RECT 269.835 49.655 270.095 49.975 ;
        RECT 270.295 49.655 270.555 49.975 ;
        RECT 269.895 49.150 270.035 49.655 ;
        RECT 269.825 48.780 270.105 49.150 ;
        RECT 269.375 48.295 269.635 48.615 ;
        RECT 269.835 47.790 270.095 47.935 ;
        RECT 269.825 47.420 270.105 47.790 ;
        RECT 269.835 46.935 270.095 47.255 ;
        RECT 269.895 46.235 270.035 46.935 ;
        RECT 269.835 45.915 270.095 46.235 ;
        RECT 268.915 45.575 269.175 45.895 ;
        RECT 268.455 45.235 268.715 45.555 ;
        RECT 269.365 45.380 269.645 45.750 ;
        RECT 270.355 45.555 270.495 49.655 ;
        RECT 271.735 49.575 273.255 49.715 ;
        RECT 271.735 48.955 271.875 49.575 ;
        RECT 271.675 48.635 271.935 48.955 ;
        RECT 272.135 48.635 272.395 48.955 ;
        RECT 271.215 47.615 271.475 47.935 ;
        RECT 271.675 47.615 271.935 47.935 ;
        RECT 269.435 45.215 269.575 45.380 ;
        RECT 270.295 45.235 270.555 45.555 ;
        RECT 269.375 44.895 269.635 45.215 ;
        RECT 271.275 43.515 271.415 47.615 ;
        RECT 271.735 45.895 271.875 47.615 ;
        RECT 272.195 45.895 272.335 48.635 ;
        RECT 273.115 48.615 273.255 49.575 ;
        RECT 273.055 48.295 273.315 48.615 ;
        RECT 273.575 47.935 273.715 49.995 ;
        RECT 274.955 49.975 275.095 53.055 ;
        RECT 278.175 50.655 278.315 53.055 ;
        RECT 280.415 52.375 280.675 52.695 ;
        RECT 280.475 50.995 280.615 52.375 ;
        RECT 285.995 51.335 286.135 53.055 ;
        RECT 288.295 51.335 288.435 53.055 ;
        RECT 288.695 52.715 288.955 53.035 ;
        RECT 285.935 51.015 286.195 51.335 ;
        RECT 288.235 51.015 288.495 51.335 ;
        RECT 279.495 50.675 279.755 50.995 ;
        RECT 280.415 50.675 280.675 50.995 ;
        RECT 277.655 50.335 277.915 50.655 ;
        RECT 278.115 50.335 278.375 50.655 ;
        RECT 274.895 49.655 275.155 49.975 ;
        RECT 276.735 49.655 276.995 49.975 ;
        RECT 272.595 47.615 272.855 47.935 ;
        RECT 273.515 47.615 273.775 47.935 ;
        RECT 271.675 45.575 271.935 45.895 ;
        RECT 272.135 45.575 272.395 45.895 ;
        RECT 272.135 44.215 272.395 44.535 ;
        RECT 271.215 43.195 271.475 43.515 ;
        RECT 267.535 43.085 267.795 43.175 ;
        RECT 266.675 42.945 267.795 43.085 ;
        RECT 265.695 41.835 265.955 42.095 ;
        RECT 262.015 41.495 262.275 41.815 ;
        RECT 262.075 40.115 262.215 41.495 ;
        RECT 262.015 39.795 262.275 40.115 ;
        RECT 264.775 39.455 265.035 39.775 ;
        RECT 261.555 38.775 261.815 39.095 ;
        RECT 261.095 37.075 261.355 37.395 ;
        RECT 261.615 36.715 261.755 38.775 ;
        RECT 264.835 37.395 264.975 39.455 ;
        RECT 264.775 37.075 265.035 37.395 ;
        RECT 261.555 36.395 261.815 36.715 ;
        RECT 258.335 36.055 258.595 36.375 ;
        RECT 255.115 35.035 255.375 35.355 ;
        RECT 260.635 35.035 260.895 35.355 ;
        RECT 254.475 32.800 256.015 33.170 ;
        RECT 260.695 32.295 260.835 35.035 ;
        RECT 260.635 31.975 260.895 32.295 ;
        RECT 253.735 31.295 253.995 31.615 ;
        RECT 264.835 29.235 264.975 37.075 ;
        RECT 265.755 35.015 265.895 41.835 ;
        RECT 265.695 34.695 265.955 35.015 ;
        RECT 265.235 34.355 265.495 34.675 ;
        RECT 265.295 32.635 265.435 34.355 ;
        RECT 265.235 32.315 265.495 32.635 ;
        RECT 265.755 31.615 265.895 34.695 ;
        RECT 265.695 31.295 265.955 31.615 ;
        RECT 264.775 28.915 265.035 29.235 ;
        RECT 254.475 27.360 256.015 27.730 ;
        RECT 265.755 27.195 265.895 31.295 ;
        RECT 265.695 26.875 265.955 27.195 ;
        RECT 266.675 26.175 266.815 42.945 ;
        RECT 267.535 42.855 267.795 42.945 ;
        RECT 268.915 42.175 269.175 42.495 ;
        RECT 268.975 40.795 269.115 42.175 ;
        RECT 268.915 40.475 269.175 40.795 ;
        RECT 272.195 40.455 272.335 44.215 ;
        RECT 272.655 42.155 272.795 47.615 ;
        RECT 274.895 46.935 275.155 47.255 ;
        RECT 273.105 46.400 274.645 46.770 ;
        RECT 274.955 46.235 275.095 46.935 ;
        RECT 274.895 45.915 275.155 46.235 ;
        RECT 276.795 42.495 276.935 49.655 ;
        RECT 277.185 47.420 277.465 47.790 ;
        RECT 277.255 43.175 277.395 47.420 ;
        RECT 277.715 46.235 277.855 50.335 ;
        RECT 278.175 47.935 278.315 50.335 ;
        RECT 278.115 47.615 278.375 47.935 ;
        RECT 277.655 45.915 277.915 46.235 ;
        RECT 277.195 42.855 277.455 43.175 ;
        RECT 276.735 42.175 276.995 42.495 ;
        RECT 272.595 41.835 272.855 42.155 ;
        RECT 273.105 40.960 274.645 41.330 ;
        RECT 277.715 40.455 277.855 45.915 ;
        RECT 278.175 45.750 278.315 47.615 ;
        RECT 279.555 47.595 279.695 50.675 ;
        RECT 283.175 49.995 283.435 50.315 ;
        RECT 282.255 49.655 282.515 49.975 ;
        RECT 281.785 48.780 282.065 49.150 ;
        RECT 281.855 47.935 281.995 48.780 ;
        RECT 280.875 47.615 281.135 47.935 ;
        RECT 281.795 47.615 282.055 47.935 ;
        RECT 279.495 47.275 279.755 47.595 ;
        RECT 278.575 46.935 278.835 47.255 ;
        RECT 278.105 45.380 278.385 45.750 ;
        RECT 272.135 40.135 272.395 40.455 ;
        RECT 277.655 40.135 277.915 40.455 ;
        RECT 271.215 39.455 271.475 39.775 ;
        RECT 270.755 38.775 271.015 39.095 ;
        RECT 270.815 37.055 270.955 38.775 ;
        RECT 271.275 38.075 271.415 39.455 ;
        RECT 271.215 37.755 271.475 38.075 ;
        RECT 270.755 36.735 271.015 37.055 ;
        RECT 267.075 36.285 267.335 36.375 ;
        RECT 267.075 36.145 267.735 36.285 ;
        RECT 267.075 36.055 267.335 36.145 ;
        RECT 267.595 29.575 267.735 36.145 ;
        RECT 269.835 36.055 270.095 36.375 ;
        RECT 269.895 35.015 270.035 36.055 ;
        RECT 269.835 34.695 270.095 35.015 ;
        RECT 270.815 34.870 270.955 36.735 ;
        RECT 270.745 34.500 271.025 34.870 ;
        RECT 272.195 34.675 272.335 40.135 ;
        RECT 278.175 37.395 278.315 45.380 ;
        RECT 278.635 40.115 278.775 46.935 ;
        RECT 279.555 42.495 279.695 47.275 ;
        RECT 280.935 43.175 281.075 47.615 ;
        RECT 282.315 43.515 282.455 49.655 ;
        RECT 282.255 43.195 282.515 43.515 ;
        RECT 280.875 42.855 281.135 43.175 ;
        RECT 279.495 42.405 279.755 42.495 ;
        RECT 279.495 42.265 280.155 42.405 ;
        RECT 279.495 42.175 279.755 42.265 ;
        RECT 280.015 40.115 280.155 42.265 ;
        RECT 280.935 40.795 281.075 42.855 ;
        RECT 281.335 41.835 281.595 42.155 ;
        RECT 280.875 40.475 281.135 40.795 ;
        RECT 281.395 40.115 281.535 41.835 ;
        RECT 281.795 41.495 282.055 41.815 ;
        RECT 278.575 39.795 278.835 40.115 ;
        RECT 279.955 39.795 280.215 40.115 ;
        RECT 281.335 39.795 281.595 40.115 ;
        RECT 280.015 39.435 280.155 39.795 ;
        RECT 279.955 39.115 280.215 39.435 ;
        RECT 281.855 37.395 281.995 41.495 ;
        RECT 282.315 40.115 282.455 43.195 ;
        RECT 283.235 42.155 283.375 49.995 ;
        RECT 285.475 49.655 285.735 49.975 ;
        RECT 285.535 47.255 285.675 49.655 ;
        RECT 285.475 46.935 285.735 47.255 ;
        RECT 288.755 45.895 288.895 52.715 ;
        RECT 290.995 52.375 291.255 52.695 ;
        RECT 290.535 47.275 290.795 47.595 ;
        RECT 290.595 46.235 290.735 47.275 ;
        RECT 290.535 45.915 290.795 46.235 ;
        RECT 287.775 45.575 288.035 45.895 ;
        RECT 288.695 45.575 288.955 45.895 ;
        RECT 284.095 44.555 284.355 44.875 ;
        RECT 284.155 42.835 284.295 44.555 ;
        RECT 284.095 42.515 284.355 42.835 ;
        RECT 285.935 42.175 286.195 42.495 ;
        RECT 283.175 41.835 283.435 42.155 ;
        RECT 285.995 40.795 286.135 42.175 ;
        RECT 285.935 40.475 286.195 40.795 ;
        RECT 282.255 39.795 282.515 40.115 ;
        RECT 283.635 37.755 283.895 38.075 ;
        RECT 282.255 37.415 282.515 37.735 ;
        RECT 278.115 37.075 278.375 37.395 ;
        RECT 281.795 37.075 282.055 37.395 ;
        RECT 276.275 36.735 276.535 37.055 ;
        RECT 272.595 36.395 272.855 36.715 ;
        RECT 272.135 34.355 272.395 34.675 ;
        RECT 269.375 33.335 269.635 33.655 ;
        RECT 269.435 30.935 269.575 33.335 ;
        RECT 269.375 30.615 269.635 30.935 ;
        RECT 267.535 29.255 267.795 29.575 ;
        RECT 269.435 28.895 269.575 30.615 ;
        RECT 272.195 29.575 272.335 34.355 ;
        RECT 272.655 31.275 272.795 36.395 ;
        RECT 273.105 35.520 274.645 35.890 ;
        RECT 275.815 33.565 276.075 33.655 ;
        RECT 276.335 33.565 276.475 36.735 ;
        RECT 279.495 36.395 279.755 36.715 ;
        RECT 279.955 36.395 280.215 36.715 ;
        RECT 277.195 36.055 277.455 36.375 ;
        RECT 275.815 33.425 276.475 33.565 ;
        RECT 275.815 33.335 276.075 33.425 ;
        RECT 276.335 31.615 276.475 33.425 ;
        RECT 276.735 32.315 276.995 32.635 ;
        RECT 276.275 31.295 276.535 31.615 ;
        RECT 272.595 30.955 272.855 31.275 ;
        RECT 273.105 30.080 274.645 30.450 ;
        RECT 272.135 29.255 272.395 29.575 ;
        RECT 276.795 28.895 276.935 32.315 ;
        RECT 277.255 29.915 277.395 36.055 ;
        RECT 279.035 34.355 279.295 34.675 ;
        RECT 279.095 31.955 279.235 34.355 ;
        RECT 279.555 31.955 279.695 36.395 ;
        RECT 280.015 34.335 280.155 36.395 ;
        RECT 281.335 36.055 281.595 36.375 ;
        RECT 280.875 34.695 281.135 35.015 ;
        RECT 279.955 34.015 280.215 34.335 ;
        RECT 280.015 32.295 280.155 34.015 ;
        RECT 279.955 31.975 280.215 32.295 ;
        RECT 279.035 31.635 279.295 31.955 ;
        RECT 279.495 31.635 279.755 31.955 ;
        RECT 279.035 30.955 279.295 31.275 ;
        RECT 277.655 30.615 277.915 30.935 ;
        RECT 277.715 29.915 277.855 30.615 ;
        RECT 277.195 29.595 277.455 29.915 ;
        RECT 277.655 29.595 277.915 29.915 ;
        RECT 279.095 29.315 279.235 30.955 ;
        RECT 278.635 29.235 279.235 29.315 ;
        RECT 278.575 29.175 279.235 29.235 ;
        RECT 278.575 28.915 278.835 29.175 ;
        RECT 269.375 28.575 269.635 28.895 ;
        RECT 276.735 28.575 276.995 28.895 ;
        RECT 279.555 28.555 279.695 31.635 ;
        RECT 280.935 29.915 281.075 34.695 ;
        RECT 281.395 29.915 281.535 36.055 ;
        RECT 282.315 31.955 282.455 37.415 ;
        RECT 283.695 37.055 283.835 37.755 ;
        RECT 283.635 36.735 283.895 37.055 ;
        RECT 286.395 36.735 286.655 37.055 ;
        RECT 285.935 36.395 286.195 36.715 ;
        RECT 283.635 36.055 283.895 36.375 ;
        RECT 283.695 32.295 283.835 36.055 ;
        RECT 285.995 35.355 286.135 36.395 ;
        RECT 285.935 35.035 286.195 35.355 ;
        RECT 285.475 34.015 285.735 34.335 ;
        RECT 284.095 33.335 284.355 33.655 ;
        RECT 283.635 31.975 283.895 32.295 ;
        RECT 282.255 31.635 282.515 31.955 ;
        RECT 282.315 31.355 282.455 31.635 ;
        RECT 282.315 31.215 283.375 31.355 ;
        RECT 282.255 30.615 282.515 30.935 ;
        RECT 282.715 30.615 282.975 30.935 ;
        RECT 282.315 29.915 282.455 30.615 ;
        RECT 282.775 29.915 282.915 30.615 ;
        RECT 280.875 29.595 281.135 29.915 ;
        RECT 281.335 29.595 281.595 29.915 ;
        RECT 282.255 29.595 282.515 29.915 ;
        RECT 282.715 29.595 282.975 29.915 ;
        RECT 283.235 29.575 283.375 31.215 ;
        RECT 283.175 29.255 283.435 29.575 ;
        RECT 284.155 29.235 284.295 33.335 ;
        RECT 285.535 32.635 285.675 34.015 ;
        RECT 286.455 33.995 286.595 36.735 ;
        RECT 286.395 33.675 286.655 33.995 ;
        RECT 285.475 32.315 285.735 32.635 ;
        RECT 287.835 31.995 287.975 45.575 ;
        RECT 288.755 33.995 288.895 45.575 ;
        RECT 291.055 45.555 291.195 52.375 ;
        RECT 291.735 49.120 293.275 49.490 ;
        RECT 293.815 48.955 293.955 53.055 ;
        RECT 295.655 51.675 295.795 56.115 ;
        RECT 302.955 54.075 303.215 54.395 ;
        RECT 298.355 52.715 298.615 53.035 ;
        RECT 295.595 51.355 295.855 51.675 ;
        RECT 294.215 51.015 294.475 51.335 ;
        RECT 293.755 48.635 294.015 48.955 ;
        RECT 291.915 46.935 292.175 47.255 ;
        RECT 291.975 45.555 292.115 46.935 ;
        RECT 293.815 46.315 293.955 48.635 ;
        RECT 294.275 48.275 294.415 51.015 ;
        RECT 297.895 50.335 298.155 50.655 ;
        RECT 295.135 49.995 295.395 50.315 ;
        RECT 294.675 49.655 294.935 49.975 ;
        RECT 294.215 47.955 294.475 48.275 ;
        RECT 294.735 47.595 294.875 49.655 ;
        RECT 294.675 47.275 294.935 47.595 ;
        RECT 293.815 46.175 294.415 46.315 ;
        RECT 295.195 46.235 295.335 49.995 ;
        RECT 295.595 47.275 295.855 47.595 ;
        RECT 296.055 47.275 296.315 47.595 ;
        RECT 290.995 45.235 291.255 45.555 ;
        RECT 291.915 45.235 292.175 45.555 ;
        RECT 293.755 45.235 294.015 45.555 ;
        RECT 289.155 44.895 289.415 45.215 ;
        RECT 289.215 43.515 289.355 44.895 ;
        RECT 291.735 43.680 293.275 44.050 ;
        RECT 289.155 43.195 289.415 43.515 ;
        RECT 291.915 43.195 292.175 43.515 ;
        RECT 289.615 41.835 289.875 42.155 ;
        RECT 289.155 41.495 289.415 41.815 ;
        RECT 288.695 33.675 288.955 33.995 ;
        RECT 289.215 33.655 289.355 41.495 ;
        RECT 289.675 40.795 289.815 41.835 ;
        RECT 289.615 40.475 289.875 40.795 ;
        RECT 291.975 40.115 292.115 43.195 ;
        RECT 293.815 40.795 293.955 45.235 ;
        RECT 294.275 43.515 294.415 46.175 ;
        RECT 295.135 45.915 295.395 46.235 ;
        RECT 294.215 43.195 294.475 43.515 ;
        RECT 295.195 40.795 295.335 45.915 ;
        RECT 295.655 41.725 295.795 47.275 ;
        RECT 296.115 46.235 296.255 47.275 ;
        RECT 297.955 47.255 298.095 50.335 ;
        RECT 297.895 46.935 298.155 47.255 ;
        RECT 296.055 45.915 296.315 46.235 ;
        RECT 297.955 45.895 298.095 46.935 ;
        RECT 297.895 45.575 298.155 45.895 ;
        RECT 297.895 42.515 298.155 42.835 ;
        RECT 296.055 41.725 296.315 41.815 ;
        RECT 295.655 41.585 296.315 41.725 ;
        RECT 296.055 41.495 296.315 41.585 ;
        RECT 296.975 41.495 297.235 41.815 ;
        RECT 293.755 40.475 294.015 40.795 ;
        RECT 295.135 40.475 295.395 40.795 ;
        RECT 290.535 39.795 290.795 40.115 ;
        RECT 291.915 39.795 292.175 40.115 ;
        RECT 295.135 39.795 295.395 40.115 ;
        RECT 289.615 37.755 289.875 38.075 ;
        RECT 289.675 35.355 289.815 37.755 ;
        RECT 290.595 37.395 290.735 39.795 ;
        RECT 291.735 38.240 293.275 38.610 ;
        RECT 295.195 38.075 295.335 39.795 ;
        RECT 295.135 37.755 295.395 38.075 ;
        RECT 296.115 37.735 296.255 41.495 ;
        RECT 296.515 39.455 296.775 39.775 ;
        RECT 296.055 37.415 296.315 37.735 ;
        RECT 296.575 37.395 296.715 39.455 ;
        RECT 290.535 37.075 290.795 37.395 ;
        RECT 296.515 37.075 296.775 37.395 ;
        RECT 297.035 36.910 297.175 41.495 ;
        RECT 295.135 36.395 295.395 36.715 ;
        RECT 296.965 36.540 297.245 36.910 ;
        RECT 289.615 35.035 289.875 35.355 ;
        RECT 294.665 34.500 294.945 34.870 ;
        RECT 290.995 33.675 291.255 33.995 ;
        RECT 289.155 33.335 289.415 33.655 ;
        RECT 287.375 31.855 287.975 31.995 ;
        RECT 291.055 31.955 291.195 33.675 ;
        RECT 293.755 33.335 294.015 33.655 ;
        RECT 291.735 32.800 293.275 33.170 ;
        RECT 293.815 32.635 293.955 33.335 ;
        RECT 294.735 32.635 294.875 34.500 ;
        RECT 293.755 32.315 294.015 32.635 ;
        RECT 294.675 32.315 294.935 32.635 ;
        RECT 287.375 31.615 287.515 31.855 ;
        RECT 290.995 31.635 291.255 31.955 ;
        RECT 287.315 31.295 287.575 31.615 ;
        RECT 295.195 29.915 295.335 36.395 ;
        RECT 297.035 35.015 297.175 36.540 ;
        RECT 296.975 34.695 297.235 35.015 ;
        RECT 295.135 29.595 295.395 29.915 ;
        RECT 297.955 29.235 298.095 42.515 ;
        RECT 298.415 42.495 298.555 52.715 ;
        RECT 303.015 51.675 303.155 54.075 ;
        RECT 302.955 51.355 303.215 51.675 ;
        RECT 300.655 44.215 300.915 44.535 ;
        RECT 300.715 42.495 300.855 44.215 ;
        RECT 304.395 43.515 304.535 69.375 ;
        RECT 305.715 68.695 305.975 69.015 ;
        RECT 305.255 61.555 305.515 61.875 ;
        RECT 305.315 58.475 305.455 61.555 ;
        RECT 305.255 58.155 305.515 58.475 ;
        RECT 305.315 56.435 305.455 58.155 ;
        RECT 305.255 56.115 305.515 56.435 ;
        RECT 305.315 51.335 305.455 56.115 ;
        RECT 305.255 51.015 305.515 51.335 ;
        RECT 305.315 47.595 305.455 51.015 ;
        RECT 305.775 50.655 305.915 68.695 ;
        RECT 305.715 50.335 305.975 50.655 ;
        RECT 305.255 47.275 305.515 47.595 ;
        RECT 305.315 45.895 305.455 47.275 ;
        RECT 305.255 45.575 305.515 45.895 ;
        RECT 305.315 43.515 305.455 45.575 ;
        RECT 304.335 43.195 304.595 43.515 ;
        RECT 305.255 43.195 305.515 43.515 ;
        RECT 298.355 42.175 298.615 42.495 ;
        RECT 300.655 42.175 300.915 42.495 ;
        RECT 302.035 39.795 302.295 40.115 ;
        RECT 299.735 38.775 299.995 39.095 ;
        RECT 299.795 37.395 299.935 38.775 ;
        RECT 302.095 37.735 302.235 39.795 ;
        RECT 302.035 37.415 302.295 37.735 ;
        RECT 299.735 37.075 299.995 37.395 ;
        RECT 298.355 36.395 298.615 36.715 ;
        RECT 298.815 36.395 299.075 36.715 ;
        RECT 298.415 35.355 298.555 36.395 ;
        RECT 298.355 35.035 298.615 35.355 ;
        RECT 298.875 34.335 299.015 36.395 ;
        RECT 300.195 35.035 300.455 35.355 ;
        RECT 300.255 34.870 300.395 35.035 ;
        RECT 302.095 35.015 302.235 37.415 ;
        RECT 304.395 37.055 304.535 43.195 ;
        RECT 305.255 42.515 305.515 42.835 ;
        RECT 305.315 38.075 305.455 42.515 ;
        RECT 305.255 37.755 305.515 38.075 ;
        RECT 304.335 36.735 304.595 37.055 ;
        RECT 303.415 36.055 303.675 36.375 ;
        RECT 303.475 35.355 303.615 36.055 ;
        RECT 303.415 35.035 303.675 35.355 ;
        RECT 300.185 34.500 300.465 34.870 ;
        RECT 302.035 34.695 302.295 35.015 ;
        RECT 298.815 34.015 299.075 34.335 ;
        RECT 303.875 31.295 304.135 31.615 ;
        RECT 303.935 29.915 304.075 31.295 ;
        RECT 305.315 31.275 305.455 37.755 ;
        RECT 306.235 31.995 306.375 85.015 ;
        RECT 306.635 74.135 306.895 74.455 ;
        RECT 306.695 64.595 306.835 74.135 ;
        RECT 306.635 64.275 306.895 64.595 ;
        RECT 307.155 54.395 307.295 100.855 ;
        RECT 308.015 96.575 308.275 96.895 ;
        RECT 308.075 82.615 308.215 96.575 ;
        RECT 308.535 90.775 308.675 105.075 ;
        RECT 308.995 100.635 309.135 109.225 ;
        RECT 310.365 106.240 311.905 106.610 ;
        RECT 309.395 101.675 309.655 101.995 ;
        RECT 308.935 100.315 309.195 100.635 ;
        RECT 309.455 100.150 309.595 101.675 ;
        RECT 310.365 100.800 311.905 101.170 ;
        RECT 309.385 99.780 309.665 100.150 ;
        RECT 310.365 95.360 311.905 95.730 ;
        RECT 308.475 90.455 308.735 90.775 ;
        RECT 308.535 89.755 308.675 90.455 ;
        RECT 310.365 89.920 311.905 90.290 ;
        RECT 308.475 89.435 308.735 89.755 ;
        RECT 310.765 86.180 311.045 86.550 ;
        RECT 310.775 86.035 311.035 86.180 ;
        RECT 310.365 84.480 311.905 84.850 ;
        RECT 308.015 82.295 308.275 82.615 ;
        RECT 310.365 79.040 311.905 79.410 ;
        RECT 310.365 73.600 311.905 73.970 ;
        RECT 310.765 69.860 311.045 70.230 ;
        RECT 310.775 69.715 311.035 69.860 ;
        RECT 310.365 68.160 311.905 68.530 ;
        RECT 310.365 62.720 311.905 63.090 ;
        RECT 310.365 57.280 311.905 57.650 ;
        RECT 310.775 56.115 311.035 56.435 ;
        RECT 308.475 55.095 308.735 55.415 ;
        RECT 307.095 54.075 307.355 54.395 ;
        RECT 307.095 52.375 307.355 52.695 ;
        RECT 307.155 45.555 307.295 52.375 ;
        RECT 307.095 45.235 307.355 45.555 ;
        RECT 308.535 40.795 308.675 55.095 ;
        RECT 310.835 54.590 310.975 56.115 ;
        RECT 310.765 54.220 311.045 54.590 ;
        RECT 308.935 53.055 309.195 53.375 ;
        RECT 308.995 51.675 309.135 53.055 ;
        RECT 310.365 51.840 311.905 52.210 ;
        RECT 308.935 51.355 309.195 51.675 ;
        RECT 310.365 46.400 311.905 46.770 ;
        RECT 308.935 44.895 309.195 45.215 ;
        RECT 308.475 40.475 308.735 40.795 ;
        RECT 308.995 40.115 309.135 44.895 ;
        RECT 310.365 40.960 311.905 41.330 ;
        RECT 308.935 39.795 309.195 40.115 ;
        RECT 308.995 34.675 309.135 39.795 ;
        RECT 310.365 35.520 311.905 35.890 ;
        RECT 316.555 35.745 318.485 36.545 ;
        RECT 308.935 34.355 309.195 34.675 ;
        RECT 308.995 31.995 309.135 34.355 ;
        RECT 305.775 31.855 306.375 31.995 ;
        RECT 308.535 31.955 309.135 31.995 ;
        RECT 308.475 31.855 309.135 31.955 ;
        RECT 305.255 30.955 305.515 31.275 ;
        RECT 305.315 29.915 305.455 30.955 ;
        RECT 303.875 29.595 304.135 29.915 ;
        RECT 305.255 29.595 305.515 29.915 ;
        RECT 305.775 29.575 305.915 31.855 ;
        RECT 308.475 31.635 308.735 31.855 ;
        RECT 305.715 29.255 305.975 29.575 ;
        RECT 308.535 29.235 308.675 31.635 ;
        RECT 310.365 30.080 311.905 30.450 ;
        RECT 284.095 28.915 284.355 29.235 ;
        RECT 297.895 28.915 298.155 29.235 ;
        RECT 308.475 28.915 308.735 29.235 ;
        RECT 279.495 28.235 279.755 28.555 ;
        RECT 291.735 27.360 293.275 27.730 ;
        RECT 266.615 25.855 266.875 26.175 ;
        RECT 273.105 24.640 274.645 25.010 ;
        RECT 310.365 24.640 311.905 25.010 ;
        RECT 254.475 21.920 256.015 22.290 ;
        RECT 291.735 21.920 293.275 22.290 ;
        RECT 10.170 18.105 74.550 20.485 ;
        RECT 79.810 19.165 127.975 20.265 ;
        RECT 248.665 20.220 248.945 20.590 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 198.585 19.200 200.125 19.570 ;
        RECT 235.845 19.200 237.385 19.570 ;
        RECT 273.105 19.200 274.645 19.570 ;
        RECT 310.365 19.200 311.905 19.570 ;
        RECT 10.170 15.580 74.550 17.080 ;
        RECT 179.955 16.480 181.495 16.850 ;
        RECT 217.215 16.480 218.755 16.850 ;
        RECT 254.475 16.480 256.015 16.850 ;
        RECT 291.735 16.480 293.275 16.850 ;
        RECT 10.170 13.580 74.550 15.080 ;
        RECT 198.585 13.760 200.125 14.130 ;
        RECT 235.845 13.760 237.385 14.130 ;
        RECT 273.105 13.760 274.645 14.130 ;
        RECT 310.365 13.760 311.905 14.130 ;
        RECT 10.170 11.580 74.550 13.080 ;
        RECT 10.170 9.555 74.550 10.555 ;
        RECT 80.745 9.665 82.345 10.465 ;
        RECT 7.065 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.965 5.690 130.565 8.890 ;
      LAYER met3 ;
        RECT 125.730 225.710 126.530 225.760 ;
        RECT 23.260 225.160 23.660 225.560 ;
        RECT 1.000 224.760 23.660 225.160 ;
        RECT 45.340 224.760 45.740 225.560 ;
        RECT 64.710 225.310 65.510 225.710 ;
        RECT 125.730 225.410 252.160 225.710 ;
        RECT 125.730 225.360 126.530 225.410 ;
        RECT 59.190 224.760 59.990 225.160 ;
        RECT 1.000 221.560 1.400 224.760 ;
        RECT 67.470 224.710 68.270 225.110 ;
        RECT 129.395 225.050 130.195 225.100 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.110 71.030 224.510 ;
        RECT 72.990 223.510 73.790 223.910 ;
        RECT 75.700 223.310 76.100 224.860 ;
        RECT 75.700 222.910 76.500 223.310 ;
        RECT 78.545 222.710 78.945 224.860 ;
        RECT 78.545 222.310 79.345 222.710 ;
        RECT 83.980 222.110 84.380 224.860 ;
        RECT 83.980 221.710 84.780 222.110 ;
        RECT 1.000 220.760 1.800 221.560 ;
        RECT 86.740 221.510 87.140 224.860 ;
        RECT 86.740 221.110 87.540 221.510 ;
        RECT 92.260 220.910 92.660 224.860 ;
        RECT 129.375 224.750 251.225 225.050 ;
        RECT 129.395 224.700 130.195 224.750 ;
        RECT 108.865 224.515 109.665 224.615 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.915 106.460 224.450 ;
        RECT 108.865 224.215 129.040 224.515 ;
        RECT 95.070 221.515 95.370 223.650 ;
        RECT 97.830 222.115 98.130 223.650 ;
        RECT 100.590 222.715 100.890 223.650 ;
        RECT 103.350 223.315 103.650 223.650 ;
        RECT 106.060 223.615 125.010 223.915 ;
        RECT 103.350 223.015 120.980 223.315 ;
        RECT 100.590 222.415 116.950 222.715 ;
        RECT 97.830 221.815 112.920 222.115 ;
        RECT 95.070 221.215 108.890 221.515 ;
        RECT 92.260 220.510 93.060 220.910 ;
        RECT 1.000 218.590 12.150 220.190 ;
        RECT 106.340 217.515 107.940 219.915 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.920 188.640 10.720 211.890 ;
        RECT 15.720 198.970 38.920 209.370 ;
        RECT 9.520 187.840 11.120 188.640 ;
        RECT 15.720 186.970 38.920 197.370 ;
        RECT 44.120 188.440 44.920 211.890 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.520 182.990 11.120 183.790 ;
        RECT 3.600 176.050 7.510 179.250 ;
        RECT 9.920 163.040 10.720 182.990 ;
        RECT 15.720 174.970 38.920 185.370 ;
        RECT 45.870 181.190 46.670 210.555 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 47.470 182.790 48.270 204.590 ;
        RECT 108.590 202.625 108.890 221.215 ;
        RECT 109.240 207.925 109.640 219.305 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 111.820 207.925 112.220 219.305 ;
        RECT 109.240 207.525 110.490 207.925 ;
        RECT 108.540 201.825 108.940 202.625 ;
        RECT 63.550 200.610 98.400 200.615 ;
        RECT 63.550 199.815 106.330 200.610 ;
        RECT 98.400 199.810 106.330 199.815 ;
        RECT 68.970 196.830 100.300 197.630 ;
        RECT 74.545 193.735 98.000 194.535 ;
        RECT 66.295 190.655 95.650 191.455 ;
        RECT 52.860 188.465 53.660 190.065 ;
        RECT 55.320 184.940 56.920 186.540 ;
        RECT 47.470 181.990 54.670 182.790 ;
        RECT 45.870 180.390 53.020 181.190 ;
        RECT 9.520 162.240 11.120 163.040 ;
        RECT 15.720 162.970 38.920 173.370 ;
        RECT 52.220 170.440 53.020 180.390 ;
        RECT 53.870 175.290 54.670 181.990 ;
        RECT 53.870 164.840 54.670 174.240 ;
        RECT 55.720 166.640 56.520 184.940 ;
        RECT 57.020 177.390 57.820 178.990 ;
        RECT 61.980 174.370 90.220 175.170 ;
        RECT 57.020 168.290 57.820 169.890 ;
        RECT 55.320 165.840 56.920 166.640 ;
        RECT 53.470 164.040 55.070 164.840 ;
        RECT 9.920 153.790 10.720 162.240 ;
        RECT 9.520 152.990 11.120 153.790 ;
        RECT 9.920 152.915 10.720 152.990 ;
        RECT 15.720 150.970 38.920 161.370 ;
        RECT 51.570 160.190 53.170 160.990 ;
        RECT 51.970 155.790 52.770 160.190 ;
        RECT 51.570 154.990 53.170 155.790 ;
        RECT 41.830 149.410 46.630 150.210 ;
        RECT 51.970 148.290 52.770 154.990 ;
        RECT 53.870 151.990 54.670 164.040 ;
        RECT 53.470 151.190 55.070 151.990 ;
        RECT 55.720 150.240 56.520 165.840 ;
        RECT 54.920 149.440 56.520 150.240 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 61.980 143.690 62.780 174.370 ;
        RECT 3.600 132.225 7.510 135.425 ;
        RECT 9.095 134.635 18.955 143.035 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 28.140 142.890 62.780 143.690 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 20.650 131.410 21.050 138.770 ;
        RECT 61.980 135.095 62.780 142.890 ;
        RECT 70.165 172.130 84.650 172.930 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 12.915 45.565 14.515 119.215 ;
        RECT 16.165 56.765 17.765 121.615 ;
        RECT 21.615 95.165 22.415 132.545 ;
        RECT 27.065 95.165 27.865 130.795 ;
        RECT 70.165 128.125 70.965 172.130 ;
        RECT 74.940 154.795 86.100 155.595 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 145.235 75.740 154.795 ;
        RECT 94.850 150.520 95.650 190.655 ;
        RECT 80.010 149.520 95.650 150.520 ;
        RECT 74.940 144.435 86.100 145.235 ;
        RECT 63.315 103.770 64.915 123.715 ;
        RECT 65.865 110.280 67.465 127.485 ;
        RECT 75.510 123.715 77.110 135.155 ;
        RECT 80.125 133.320 80.925 144.435 ;
        RECT 94.850 131.745 95.650 149.520 ;
        RECT 97.200 137.420 98.000 193.735 ;
        RECT 99.500 129.995 100.300 196.830 ;
        RECT 102.950 168.255 103.750 186.540 ;
        RECT 105.530 170.890 106.330 199.810 ;
        RECT 109.240 198.885 109.640 205.545 ;
        RECT 110.090 197.895 110.490 207.525 ;
        RECT 109.240 197.495 110.490 197.895 ;
        RECT 110.970 207.525 112.220 207.925 ;
        RECT 110.970 197.895 111.370 207.525 ;
        RECT 111.820 198.885 112.220 206.755 ;
        RECT 112.620 202.625 112.920 221.815 ;
        RECT 113.270 207.925 113.670 219.305 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 115.850 207.925 116.250 219.305 ;
        RECT 113.270 207.525 114.520 207.925 ;
        RECT 112.570 201.825 112.970 202.625 ;
        RECT 113.270 198.885 113.670 205.545 ;
        RECT 114.120 197.895 114.520 207.525 ;
        RECT 110.970 197.495 112.220 197.895 ;
        RECT 109.240 183.970 109.640 197.495 ;
        RECT 111.820 191.285 112.220 197.495 ;
        RECT 113.270 197.495 114.520 197.895 ;
        RECT 115.000 207.525 116.250 207.925 ;
        RECT 115.000 197.895 115.400 207.525 ;
        RECT 115.850 198.885 116.250 206.755 ;
        RECT 116.650 202.625 116.950 222.415 ;
        RECT 117.300 207.925 117.700 219.305 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 119.880 207.925 120.280 219.305 ;
        RECT 117.300 207.525 118.550 207.925 ;
        RECT 116.600 201.825 117.000 202.625 ;
        RECT 117.300 198.885 117.700 205.545 ;
        RECT 118.150 197.895 118.550 207.525 ;
        RECT 115.000 197.495 116.250 197.895 ;
        RECT 110.530 187.540 110.930 189.140 ;
        RECT 113.270 183.990 113.670 197.495 ;
        RECT 115.850 191.285 116.250 197.495 ;
        RECT 117.300 197.495 118.550 197.895 ;
        RECT 119.030 207.525 120.280 207.925 ;
        RECT 119.030 197.895 119.430 207.525 ;
        RECT 119.880 198.885 120.280 206.755 ;
        RECT 120.680 202.625 120.980 223.015 ;
        RECT 121.330 207.925 121.730 219.305 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 123.910 207.925 124.310 219.305 ;
        RECT 121.330 207.525 122.580 207.925 ;
        RECT 120.630 201.825 121.030 202.625 ;
        RECT 121.330 198.885 121.730 205.545 ;
        RECT 122.180 197.895 122.580 207.525 ;
        RECT 119.030 197.495 120.280 197.895 ;
        RECT 114.560 187.540 114.960 189.140 ;
        RECT 111.685 183.590 113.670 183.990 ;
        RECT 105.530 168.255 106.730 170.890 ;
        RECT 107.380 168.490 107.780 170.890 ;
        RECT 103.350 152.765 103.750 160.495 ;
        RECT 103.350 143.435 103.750 145.835 ;
        RECT 104.640 140.165 105.040 167.190 ;
        RECT 105.385 157.365 105.785 158.165 ;
        RECT 106.330 145.835 106.730 168.255 ;
        RECT 107.380 152.765 107.780 160.495 ;
        RECT 108.670 147.135 109.070 178.990 ;
        RECT 109.960 168.490 110.760 170.890 ;
        RECT 109.415 156.165 109.815 156.965 ;
        RECT 110.360 145.835 110.760 168.490 ;
        RECT 111.685 157.765 112.085 183.590 ;
        RECT 117.300 182.580 117.700 197.495 ;
        RECT 119.880 191.285 120.280 197.495 ;
        RECT 121.330 197.495 122.580 197.895 ;
        RECT 123.060 207.525 124.310 207.925 ;
        RECT 123.060 197.895 123.460 207.525 ;
        RECT 123.910 198.885 124.310 206.755 ;
        RECT 124.710 202.625 125.010 223.615 ;
        RECT 125.360 207.925 125.760 219.305 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 127.940 207.925 128.340 219.305 ;
        RECT 125.360 207.525 126.610 207.925 ;
        RECT 124.660 201.825 125.060 202.625 ;
        RECT 125.360 198.885 125.760 205.545 ;
        RECT 126.210 197.895 126.610 207.525 ;
        RECT 123.060 197.495 124.310 197.895 ;
        RECT 118.590 187.540 118.990 189.140 ;
        RECT 113.085 182.180 117.700 182.580 ;
        RECT 113.085 156.165 113.485 182.180 ;
        RECT 121.330 181.545 121.730 197.495 ;
        RECT 123.910 191.285 124.310 197.495 ;
        RECT 125.360 197.495 126.610 197.895 ;
        RECT 127.090 207.525 128.340 207.925 ;
        RECT 127.090 197.895 127.490 207.525 ;
        RECT 127.940 198.885 128.340 206.755 ;
        RECT 128.740 202.625 129.040 224.215 ;
        RECT 132.720 220.715 133.120 221.515 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 129.390 207.925 129.790 219.305 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 131.970 207.925 132.370 219.305 ;
        RECT 129.390 207.525 130.640 207.925 ;
        RECT 128.690 201.825 129.090 202.625 ;
        RECT 129.390 198.885 129.790 205.545 ;
        RECT 130.240 197.895 130.640 207.525 ;
        RECT 127.090 197.495 128.340 197.895 ;
        RECT 122.620 187.540 123.020 189.140 ;
        RECT 116.415 181.145 121.730 181.545 ;
        RECT 116.415 176.215 116.815 181.145 ;
        RECT 125.360 180.565 125.760 197.495 ;
        RECT 127.940 191.285 128.340 197.495 ;
        RECT 129.390 197.495 130.640 197.895 ;
        RECT 131.120 207.525 132.370 207.925 ;
        RECT 131.120 197.895 131.520 207.525 ;
        RECT 131.970 198.885 132.370 206.755 ;
        RECT 132.770 202.625 133.070 220.715 ;
        RECT 133.420 207.925 133.820 219.305 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 136.000 207.925 136.400 219.305 ;
        RECT 133.420 207.525 134.670 207.925 ;
        RECT 132.720 201.825 133.120 202.625 ;
        RECT 133.420 198.885 133.820 205.545 ;
        RECT 134.270 197.895 134.670 207.525 ;
        RECT 131.120 197.495 132.370 197.895 ;
        RECT 126.650 187.540 127.050 189.140 ;
        RECT 121.035 180.165 125.760 180.565 ;
        RECT 121.035 176.215 121.435 180.165 ;
        RECT 129.390 179.490 129.790 197.495 ;
        RECT 131.970 191.285 132.370 197.495 ;
        RECT 133.420 197.495 134.670 197.895 ;
        RECT 135.150 207.525 136.400 207.925 ;
        RECT 135.150 197.895 135.550 207.525 ;
        RECT 136.000 198.885 136.400 206.755 ;
        RECT 136.800 202.625 137.100 220.715 ;
        RECT 137.450 207.925 137.850 219.305 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 140.030 207.925 140.430 219.305 ;
        RECT 137.450 207.525 138.700 207.925 ;
        RECT 136.750 201.825 137.150 202.625 ;
        RECT 137.450 198.885 137.850 205.545 ;
        RECT 138.300 197.895 138.700 207.525 ;
        RECT 135.150 197.495 136.400 197.895 ;
        RECT 130.680 187.540 131.080 189.140 ;
        RECT 125.660 179.090 129.790 179.490 ;
        RECT 125.660 176.215 126.060 179.090 ;
        RECT 133.420 178.920 133.820 197.495 ;
        RECT 136.000 191.285 136.400 197.495 ;
        RECT 137.450 197.495 138.700 197.895 ;
        RECT 139.180 207.525 140.430 207.925 ;
        RECT 139.180 197.895 139.580 207.525 ;
        RECT 140.030 198.885 140.430 206.755 ;
        RECT 140.830 202.625 141.130 220.715 ;
        RECT 141.480 207.925 141.880 219.305 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 144.060 207.925 144.460 219.305 ;
        RECT 141.480 207.525 142.730 207.925 ;
        RECT 140.780 201.825 141.180 202.625 ;
        RECT 141.480 198.885 141.880 205.545 ;
        RECT 142.330 197.895 142.730 207.525 ;
        RECT 139.180 197.495 140.430 197.895 ;
        RECT 134.710 187.540 135.110 189.140 ;
        RECT 137.450 178.920 137.850 197.495 ;
        RECT 140.030 191.285 140.430 197.495 ;
        RECT 141.480 197.495 142.730 197.895 ;
        RECT 143.210 207.525 144.460 207.925 ;
        RECT 143.210 197.895 143.610 207.525 ;
        RECT 144.060 198.885 144.460 206.755 ;
        RECT 144.860 202.625 145.160 220.715 ;
        RECT 145.510 207.925 145.910 219.305 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 148.090 207.925 148.490 219.305 ;
        RECT 145.510 207.525 146.760 207.925 ;
        RECT 144.810 201.825 145.210 202.625 ;
        RECT 145.510 198.885 145.910 205.545 ;
        RECT 146.360 197.895 146.760 207.525 ;
        RECT 143.210 197.495 144.460 197.895 ;
        RECT 138.740 187.540 139.140 189.140 ;
        RECT 141.480 178.920 141.880 197.495 ;
        RECT 144.060 191.285 144.460 197.495 ;
        RECT 145.510 197.495 146.760 197.895 ;
        RECT 147.240 207.525 148.490 207.925 ;
        RECT 147.240 197.895 147.640 207.525 ;
        RECT 148.090 198.885 148.490 206.755 ;
        RECT 148.890 202.625 149.190 220.715 ;
        RECT 162.100 220.260 162.500 220.910 ;
        RECT 163.100 220.860 163.500 221.510 ;
        RECT 164.100 221.460 164.500 222.110 ;
        RECT 164.100 221.160 250.220 221.460 ;
        RECT 163.100 220.560 249.370 220.860 ;
        RECT 162.100 219.960 248.285 220.260 ;
        RECT 149.540 207.925 149.940 219.305 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 152.120 207.925 152.520 219.305 ;
        RECT 246.615 217.650 247.015 218.450 ;
        RECT 149.540 207.525 150.790 207.925 ;
        RECT 148.840 201.825 149.240 202.625 ;
        RECT 149.540 198.885 149.940 205.545 ;
        RECT 150.390 197.895 150.790 207.525 ;
        RECT 147.240 197.495 148.490 197.895 ;
        RECT 142.770 187.540 143.170 189.140 ;
        RECT 145.510 178.920 145.910 197.495 ;
        RECT 148.090 191.285 148.490 197.495 ;
        RECT 149.540 197.495 150.790 197.895 ;
        RECT 151.270 207.525 152.520 207.925 ;
        RECT 151.270 197.895 151.670 207.525 ;
        RECT 152.120 198.885 152.520 206.755 ;
        RECT 173.615 201.325 175.195 201.655 ;
        RECT 192.125 201.325 193.705 201.655 ;
        RECT 210.635 201.325 212.215 201.655 ;
        RECT 229.145 201.325 230.725 201.655 ;
        RECT 182.870 198.605 184.450 198.935 ;
        RECT 201.380 198.605 202.960 198.935 ;
        RECT 219.890 198.605 221.470 198.935 ;
        RECT 238.400 198.605 239.980 198.935 ;
        RECT 162.390 197.900 164.390 198.050 ;
        RECT 166.595 197.900 166.925 197.915 ;
        RECT 151.270 197.495 152.520 197.895 ;
        RECT 146.800 187.540 147.200 189.140 ;
        RECT 149.540 178.920 149.940 197.495 ;
        RECT 152.120 191.285 152.520 197.495 ;
        RECT 159.185 197.600 166.925 197.900 ;
        RECT 150.830 187.540 151.230 189.140 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 158.335 187.580 158.735 188.380 ;
        RECT 130.275 178.520 133.820 178.920 ;
        RECT 134.895 178.520 137.850 178.920 ;
        RECT 139.510 178.520 141.880 178.920 ;
        RECT 144.135 178.520 145.910 178.920 ;
        RECT 148.755 178.520 149.940 178.920 ;
        RECT 130.275 176.215 130.675 178.520 ;
        RECT 134.895 176.215 135.295 178.520 ;
        RECT 139.510 176.215 139.910 178.520 ;
        RECT 144.135 176.215 144.535 178.520 ;
        RECT 148.755 176.215 149.155 178.520 ;
        RECT 116.215 175.815 117.015 176.215 ;
        RECT 120.835 175.815 121.635 176.215 ;
        RECT 125.455 175.815 126.255 176.215 ;
        RECT 130.075 175.815 130.875 176.215 ;
        RECT 134.695 175.815 135.495 176.215 ;
        RECT 139.315 175.815 140.115 176.215 ;
        RECT 143.935 175.815 144.735 176.215 ;
        RECT 148.555 175.815 149.355 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 115.815 173.070 117.415 173.870 ;
        RECT 120.435 173.070 122.035 173.870 ;
        RECT 125.055 173.070 126.655 173.870 ;
        RECT 129.675 173.070 131.275 173.870 ;
        RECT 134.295 173.070 135.895 173.870 ;
        RECT 138.915 173.070 140.515 173.870 ;
        RECT 143.535 173.070 145.135 173.870 ;
        RECT 148.155 173.070 149.755 173.870 ;
        RECT 105.930 143.435 106.730 145.835 ;
        RECT 104.640 139.365 105.440 140.165 ;
        RECT 107.380 136.325 107.780 145.835 ;
        RECT 109.960 143.435 110.760 145.835 ;
        RECT 116.310 144.730 116.910 173.070 ;
        RECT 120.930 147.530 121.530 173.070 ;
        RECT 125.550 148.690 126.150 173.070 ;
        RECT 130.175 149.890 130.775 173.070 ;
        RECT 134.795 160.260 135.395 173.070 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 133.275 152.100 134.875 152.200 ;
        RECT 136.875 152.100 137.475 161.650 ;
        RECT 133.275 151.500 137.475 152.100 ;
        RECT 133.275 151.400 134.875 151.500 ;
        RECT 133.275 150.930 134.875 151.030 ;
        RECT 139.410 150.930 140.010 173.070 ;
        RECT 144.035 162.450 144.635 173.070 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 148.655 161.210 149.255 173.070 ;
        RECT 133.275 150.330 140.010 150.930 ;
        RECT 141.715 160.610 149.255 161.210 ;
        RECT 133.275 150.230 134.875 150.330 ;
        RECT 130.175 149.290 136.695 149.890 ;
        RECT 125.550 148.090 133.635 148.690 ;
        RECT 130.615 147.530 132.215 147.630 ;
        RECT 120.930 146.930 132.215 147.530 ;
        RECT 130.615 146.830 132.215 146.930 ;
        RECT 122.645 144.730 124.245 144.830 ;
        RECT 116.310 144.130 124.245 144.730 ;
        RECT 122.645 144.030 124.245 144.130 ;
        RECT 133.035 144.520 133.635 148.090 ;
        RECT 136.095 148.010 136.695 149.290 ;
        RECT 138.525 148.010 140.125 148.110 ;
        RECT 136.095 147.410 140.125 148.010 ;
        RECT 138.525 147.310 140.125 147.410 ;
        RECT 138.525 144.520 140.125 144.620 ;
        RECT 133.035 143.920 140.125 144.520 ;
        RECT 141.715 144.040 142.315 160.610 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 138.525 143.820 140.125 143.920 ;
        RECT 109.960 138.220 110.360 143.435 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 142.690 142.815 142.790 ;
        RECT 145.625 142.690 146.225 159.460 ;
        RECT 141.215 142.090 146.225 142.690 ;
        RECT 141.215 141.990 142.815 142.090 ;
        RECT 109.560 137.420 110.760 138.220 ;
        RECT 107.380 135.525 108.180 136.325 ;
        RECT 72.765 103.865 74.365 122.215 ;
        RECT 75.510 114.215 77.115 123.715 ;
        RECT 75.515 100.215 77.115 114.215 ;
        RECT 21.215 51.675 22.815 95.165 ;
        RECT 26.665 61.465 28.265 95.165 ;
        RECT 97.165 93.265 98.765 119.215 ;
        RECT 100.515 117.715 101.315 128.925 ;
        RECT 100.115 96.415 101.715 117.715 ;
        RECT 103.315 111.365 104.915 123.165 ;
        RECT 116.915 121.965 118.515 122.765 ;
        RECT 105.965 103.965 107.565 120.665 ;
        RECT 109.865 108.365 111.465 119.215 ;
        RECT 117.115 108.365 118.715 118.265 ;
        RECT 121.565 113.015 123.165 127.485 ;
        RECT 116.965 104.015 118.565 104.815 ;
        RECT 42.740 71.190 53.140 83.050 ;
        RECT 55.740 71.190 66.140 83.050 ;
        RECT 68.740 71.190 79.140 83.050 ;
        RECT 81.740 71.190 92.140 83.050 ;
        RECT 94.740 71.190 105.140 83.050 ;
        RECT 42.740 57.830 53.140 69.690 ;
        RECT 55.740 57.830 66.140 69.690 ;
        RECT 68.740 57.830 79.140 69.690 ;
        RECT 81.740 57.830 92.140 69.690 ;
        RECT 94.740 57.830 105.140 69.690 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 3.600 36.430 8.665 39.630 ;
        RECT 3.600 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 34.940 ;
        RECT 65.765 15.915 67.365 44.215 ;
        RECT 68.865 11.965 70.465 41.615 ;
        RECT 72.095 9.665 73.695 38.865 ;
        RECT 80.745 9.665 82.345 37.635 ;
        RECT 84.015 22.315 85.615 41.615 ;
        RECT 87.165 26.815 88.765 44.215 ;
        RECT 90.715 19.315 92.315 47.165 ;
        RECT 116.115 42.615 117.715 90.815 ;
        RECT 119.215 40.015 120.815 84.315 ;
        RECT 123.215 23.815 124.815 94.865 ;
        RECT 126.165 25.365 127.765 98.015 ;
        RECT 128.965 5.690 130.565 8.890 ;
        RECT 2.705 1.285 98.380 2.085 ;
        RECT 131.665 1.800 132.465 136.325 ;
        RECT 133.265 111.795 134.065 130.795 ;
        RECT 134.865 110.315 135.665 132.545 ;
        RECT 136.465 114.770 137.265 134.120 ;
        RECT 137.945 133.410 138.745 133.810 ;
        RECT 137.945 131.410 138.345 133.410 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.970 125.690 142.100 127.290 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 133.525 109.515 138.400 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 136.495 29.375 138.195 94.305 ;
        RECT 139.355 30.545 141.055 114.150 ;
        RECT 141.900 110.315 142.700 117.170 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 141.495 20.015 143.195 110.315 ;
        RECT 143.640 32.885 145.340 114.150 ;
        RECT 146.950 110.315 147.750 138.220 ;
        RECT 149.945 116.370 150.745 170.845 ;
        RECT 146.490 104.255 148.190 110.315 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 151.560 1.800 152.360 140.165 ;
        RECT 153.945 129.145 154.345 184.370 ;
        RECT 157.560 178.060 157.960 178.860 ;
        RECT 157.560 28.035 157.860 178.060 ;
        RECT 158.335 60.675 158.635 187.580 ;
        RECT 159.185 93.465 159.485 197.600 ;
        RECT 162.390 197.450 164.390 197.600 ;
        RECT 166.595 197.585 166.925 197.600 ;
        RECT 173.615 195.885 175.195 196.215 ;
        RECT 192.125 195.885 193.705 196.215 ;
        RECT 210.635 195.885 212.215 196.215 ;
        RECT 229.145 195.885 230.725 196.215 ;
        RECT 190.975 195.190 191.305 195.195 ;
        RECT 190.975 195.180 191.560 195.190 ;
        RECT 190.975 194.880 191.760 195.180 ;
        RECT 190.975 194.870 191.560 194.880 ;
        RECT 190.975 194.865 191.305 194.870 ;
        RECT 182.870 193.165 184.450 193.495 ;
        RECT 201.380 193.165 202.960 193.495 ;
        RECT 219.890 193.165 221.470 193.495 ;
        RECT 238.400 193.165 239.980 193.495 ;
        RECT 173.615 190.445 175.195 190.775 ;
        RECT 192.125 190.445 193.705 190.775 ;
        RECT 210.635 190.445 212.215 190.775 ;
        RECT 229.145 190.445 230.725 190.775 ;
        RECT 213.300 190.120 224.640 190.420 ;
        RECT 175.335 189.750 175.665 189.755 ;
        RECT 175.335 189.740 175.920 189.750 ;
        RECT 187.500 189.740 187.880 189.750 ;
        RECT 175.335 189.440 176.120 189.740 ;
        RECT 179.260 189.440 187.880 189.740 ;
        RECT 175.335 189.430 175.920 189.440 ;
        RECT 175.335 189.425 175.665 189.430 ;
        RECT 170.735 189.060 171.065 189.075 ;
        RECT 179.260 189.060 179.560 189.440 ;
        RECT 187.500 189.430 187.880 189.440 ;
        RECT 196.495 189.740 196.825 189.755 ;
        RECT 213.300 189.740 213.600 190.120 ;
        RECT 196.495 189.440 213.600 189.740 ;
        RECT 216.940 189.740 217.320 189.750 ;
        RECT 224.340 189.740 224.640 190.120 ;
        RECT 227.315 189.740 227.645 189.755 ;
        RECT 216.940 189.440 220.040 189.740 ;
        RECT 224.340 189.440 227.645 189.740 ;
        RECT 196.495 189.425 196.825 189.440 ;
        RECT 216.940 189.430 217.320 189.440 ;
        RECT 170.735 188.760 179.560 189.060 ;
        RECT 180.395 189.060 180.725 189.075 ;
        RECT 181.980 189.060 182.360 189.070 ;
        RECT 180.395 188.760 182.360 189.060 ;
        RECT 170.735 188.745 171.065 188.760 ;
        RECT 180.395 188.745 180.725 188.760 ;
        RECT 181.980 188.750 182.360 188.760 ;
        RECT 210.295 189.060 210.625 189.075 ;
        RECT 218.780 189.060 219.160 189.070 ;
        RECT 210.295 188.760 219.160 189.060 ;
        RECT 219.740 189.060 220.040 189.440 ;
        RECT 227.315 189.425 227.645 189.440 ;
        RECT 230.075 189.060 230.405 189.075 ;
        RECT 219.740 188.760 230.405 189.060 ;
        RECT 210.295 188.745 210.625 188.760 ;
        RECT 218.780 188.750 219.160 188.760 ;
        RECT 230.075 188.745 230.405 188.760 ;
        RECT 162.390 188.430 164.390 188.530 ;
        RECT 161.590 188.380 164.390 188.430 ;
        RECT 166.595 188.380 166.925 188.395 ;
        RECT 161.590 188.080 166.925 188.380 ;
        RECT 161.590 188.030 164.390 188.080 ;
        RECT 166.595 188.065 166.925 188.080 ;
        RECT 169.815 188.380 170.145 188.395 ;
        RECT 177.175 188.380 177.505 188.395 ;
        RECT 169.815 188.080 177.505 188.380 ;
        RECT 169.815 188.065 170.145 188.080 ;
        RECT 177.175 188.065 177.505 188.080 ;
        RECT 190.260 188.380 190.640 188.390 ;
        RECT 191.895 188.380 192.225 188.395 ;
        RECT 190.260 188.080 192.225 188.380 ;
        RECT 190.260 188.070 190.640 188.080 ;
        RECT 191.895 188.065 192.225 188.080 ;
        RECT 162.390 187.930 164.390 188.030 ;
        RECT 182.870 187.725 184.450 188.055 ;
        RECT 201.380 187.725 202.960 188.055 ;
        RECT 219.890 187.725 221.470 188.055 ;
        RECT 238.400 187.725 239.980 188.055 ;
        RECT 190.515 187.700 190.845 187.715 ;
        RECT 200.175 187.700 200.505 187.715 ;
        RECT 190.515 187.400 200.505 187.700 ;
        RECT 190.515 187.385 190.845 187.400 ;
        RECT 200.175 187.385 200.505 187.400 ;
        RECT 227.315 187.700 227.645 187.715 ;
        RECT 234.215 187.700 234.545 187.715 ;
        RECT 227.315 187.400 234.545 187.700 ;
        RECT 227.315 187.385 227.645 187.400 ;
        RECT 234.215 187.385 234.545 187.400 ;
        RECT 175.335 187.020 175.665 187.035 ;
        RECT 207.995 187.020 208.325 187.035 ;
        RECT 175.335 186.720 208.325 187.020 ;
        RECT 175.335 186.705 175.665 186.720 ;
        RECT 207.995 186.705 208.325 186.720 ;
        RECT 212.135 187.020 212.465 187.035 ;
        RECT 213.260 187.020 213.640 187.030 ;
        RECT 212.135 186.720 213.640 187.020 ;
        RECT 212.135 186.705 212.465 186.720 ;
        RECT 213.260 186.710 213.640 186.720 ;
        RECT 227.775 187.020 228.105 187.035 ;
        RECT 233.755 187.020 234.085 187.035 ;
        RECT 227.775 186.720 234.085 187.020 ;
        RECT 227.775 186.705 228.105 186.720 ;
        RECT 233.755 186.705 234.085 186.720 ;
        RECT 179.015 186.340 179.345 186.355 ;
        RECT 184.535 186.340 184.865 186.355 ;
        RECT 179.015 186.040 184.865 186.340 ;
        RECT 179.015 186.025 179.345 186.040 ;
        RECT 184.535 186.025 184.865 186.040 ;
        RECT 199.255 186.340 199.585 186.355 ;
        RECT 231.915 186.340 232.245 186.355 ;
        RECT 199.255 186.040 232.245 186.340 ;
        RECT 199.255 186.025 199.585 186.040 ;
        RECT 231.915 186.025 232.245 186.040 ;
        RECT 180.395 185.660 180.725 185.675 ;
        RECT 185.660 185.660 186.040 185.670 ;
        RECT 190.515 185.660 190.845 185.675 ;
        RECT 180.395 185.360 186.040 185.660 ;
        RECT 180.395 185.345 180.725 185.360 ;
        RECT 185.660 185.350 186.040 185.360 ;
        RECT 186.620 185.360 190.845 185.660 ;
        RECT 173.615 185.005 175.195 185.335 ;
        RECT 182.235 184.980 182.565 184.995 ;
        RECT 184.740 184.980 185.120 184.990 ;
        RECT 182.235 184.680 185.120 184.980 ;
        RECT 182.235 184.665 182.565 184.680 ;
        RECT 184.740 184.670 185.120 184.680 ;
        RECT 173.955 184.300 174.285 184.315 ;
        RECT 186.620 184.300 186.920 185.360 ;
        RECT 190.515 185.345 190.845 185.360 ;
        RECT 215.815 185.660 216.145 185.675 ;
        RECT 225.015 185.660 225.345 185.675 ;
        RECT 215.815 185.360 225.345 185.660 ;
        RECT 215.815 185.345 216.145 185.360 ;
        RECT 225.015 185.345 225.345 185.360 ;
        RECT 192.125 185.005 193.705 185.335 ;
        RECT 210.635 185.005 212.215 185.335 ;
        RECT 229.145 185.005 230.725 185.335 ;
        RECT 187.500 184.670 187.880 184.990 ;
        RECT 188.215 184.980 188.545 184.995 ;
        RECT 191.435 184.980 191.765 184.995 ;
        RECT 188.215 184.680 191.765 184.980 ;
        RECT 173.955 184.000 186.920 184.300 ;
        RECT 187.540 184.315 187.840 184.670 ;
        RECT 188.215 184.665 188.545 184.680 ;
        RECT 191.435 184.665 191.765 184.680 ;
        RECT 195.115 184.980 195.445 184.995 ;
        RECT 202.015 184.980 202.345 184.995 ;
        RECT 195.115 184.680 202.345 184.980 ;
        RECT 195.115 184.665 195.445 184.680 ;
        RECT 202.015 184.665 202.345 184.680 ;
        RECT 213.515 184.980 213.845 184.995 ;
        RECT 223.635 184.980 223.965 184.995 ;
        RECT 213.515 184.680 223.965 184.980 ;
        RECT 213.515 184.665 213.845 184.680 ;
        RECT 223.635 184.665 223.965 184.680 ;
        RECT 187.540 184.000 188.085 184.315 ;
        RECT 199.715 184.300 200.045 184.315 ;
        RECT 173.955 183.985 174.285 184.000 ;
        RECT 187.755 183.985 188.085 184.000 ;
        RECT 197.660 184.000 200.045 184.300 ;
        RECT 168.435 183.620 168.765 183.635 ;
        RECT 196.495 183.620 196.825 183.635 ;
        RECT 168.435 183.320 196.825 183.620 ;
        RECT 168.435 183.305 168.765 183.320 ;
        RECT 196.495 183.305 196.825 183.320 ;
        RECT 172.575 182.940 172.905 182.955 ;
        RECT 178.555 182.940 178.885 182.955 ;
        RECT 180.855 182.940 181.185 182.955 ;
        RECT 172.575 182.640 174.960 182.940 ;
        RECT 172.575 182.625 172.905 182.640 ;
        RECT 174.660 182.260 174.960 182.640 ;
        RECT 178.555 182.640 181.185 182.940 ;
        RECT 178.555 182.625 178.885 182.640 ;
        RECT 180.855 182.625 181.185 182.640 ;
        RECT 182.870 182.285 184.450 182.615 ;
        RECT 178.555 182.260 178.885 182.275 ;
        RECT 174.660 181.960 178.885 182.260 ;
        RECT 178.555 181.945 178.885 181.960 ;
        RECT 190.055 182.260 190.385 182.275 ;
        RECT 197.660 182.260 197.960 184.000 ;
        RECT 199.715 183.985 200.045 184.000 ;
        RECT 214.895 184.300 215.225 184.315 ;
        RECT 234.215 184.300 234.545 184.315 ;
        RECT 214.895 184.000 234.545 184.300 ;
        RECT 214.895 183.985 215.225 184.000 ;
        RECT 234.215 183.985 234.545 184.000 ;
        RECT 211.675 183.620 212.005 183.635 ;
        RECT 222.460 183.620 222.840 183.630 ;
        RECT 211.675 183.320 222.840 183.620 ;
        RECT 211.675 183.305 212.005 183.320 ;
        RECT 222.460 183.310 222.840 183.320 ;
        RECT 225.015 183.620 225.345 183.635 ;
        RECT 226.395 183.620 226.725 183.635 ;
        RECT 232.375 183.620 232.705 183.635 ;
        RECT 225.015 183.320 226.725 183.620 ;
        RECT 225.015 183.305 225.345 183.320 ;
        RECT 226.395 183.305 226.725 183.320 ;
        RECT 227.100 183.320 232.705 183.620 ;
        RECT 215.100 182.940 215.480 182.950 ;
        RECT 218.115 182.940 218.445 182.955 ;
        RECT 215.100 182.640 218.445 182.940 ;
        RECT 215.100 182.630 215.480 182.640 ;
        RECT 218.115 182.625 218.445 182.640 ;
        RECT 223.175 182.940 223.505 182.955 ;
        RECT 227.100 182.940 227.400 183.320 ;
        RECT 232.375 183.305 232.705 183.320 ;
        RECT 223.175 182.640 227.400 182.940 ;
        RECT 227.775 182.940 228.105 182.955 ;
        RECT 232.835 182.940 233.165 182.955 ;
        RECT 227.775 182.640 233.165 182.940 ;
        RECT 223.175 182.625 223.505 182.640 ;
        RECT 227.775 182.625 228.105 182.640 ;
        RECT 232.835 182.625 233.165 182.640 ;
        RECT 201.380 182.285 202.960 182.615 ;
        RECT 219.890 182.285 221.470 182.615 ;
        RECT 238.400 182.285 239.980 182.615 ;
        RECT 190.055 181.960 197.960 182.260 ;
        RECT 213.515 182.260 213.845 182.275 ;
        RECT 213.515 181.960 219.350 182.260 ;
        RECT 190.055 181.945 190.385 181.960 ;
        RECT 213.515 181.945 213.845 181.960 ;
        RECT 197.415 181.580 197.745 181.595 ;
        RECT 215.815 181.580 216.145 181.595 ;
        RECT 182.020 181.280 197.745 181.580 ;
        RECT 179.935 180.900 180.265 180.915 ;
        RECT 182.020 180.900 182.320 181.280 ;
        RECT 197.415 181.265 197.745 181.280 ;
        RECT 203.180 181.280 216.145 181.580 ;
        RECT 219.050 181.580 219.350 181.960 ;
        RECT 221.335 181.580 221.665 181.595 ;
        RECT 219.050 181.280 221.665 181.580 ;
        RECT 203.180 180.915 203.480 181.280 ;
        RECT 215.815 181.265 216.145 181.280 ;
        RECT 221.335 181.265 221.665 181.280 ;
        RECT 224.095 181.580 224.425 181.595 ;
        RECT 232.835 181.580 233.165 181.595 ;
        RECT 224.095 181.280 233.165 181.580 ;
        RECT 224.095 181.265 224.425 181.280 ;
        RECT 232.835 181.265 233.165 181.280 ;
        RECT 179.935 180.600 182.320 180.900 ;
        RECT 182.695 180.900 183.025 180.915 ;
        RECT 198.335 180.900 198.665 180.915 ;
        RECT 182.695 180.600 198.665 180.900 ;
        RECT 179.935 180.585 180.265 180.600 ;
        RECT 182.695 180.585 183.025 180.600 ;
        RECT 198.335 180.585 198.665 180.600 ;
        RECT 202.935 180.600 203.480 180.915 ;
        RECT 211.675 180.900 212.005 180.915 ;
        RECT 215.815 180.900 216.145 180.915 ;
        RECT 219.035 180.900 219.365 180.915 ;
        RECT 211.675 180.600 213.370 180.900 ;
        RECT 202.935 180.585 203.265 180.600 ;
        RECT 211.675 180.585 212.005 180.600 ;
        RECT 183.615 180.220 183.945 180.235 ;
        RECT 185.915 180.230 186.245 180.235 ;
        RECT 184.740 180.220 185.120 180.230 ;
        RECT 183.615 179.920 185.120 180.220 ;
        RECT 183.615 179.905 183.945 179.920 ;
        RECT 184.740 179.910 185.120 179.920 ;
        RECT 185.660 180.220 186.245 180.230 ;
        RECT 185.660 179.920 186.470 180.220 ;
        RECT 185.660 179.910 186.245 179.920 ;
        RECT 191.180 179.910 191.560 180.230 ;
        RECT 213.070 180.220 213.370 180.600 ;
        RECT 215.815 180.600 219.365 180.900 ;
        RECT 215.815 180.585 216.145 180.600 ;
        RECT 219.035 180.585 219.365 180.600 ;
        RECT 225.935 180.900 226.265 180.915 ;
        RECT 228.695 180.900 229.025 180.915 ;
        RECT 225.935 180.600 229.025 180.900 ;
        RECT 225.935 180.585 226.265 180.600 ;
        RECT 228.695 180.585 229.025 180.600 ;
        RECT 231.915 180.900 232.245 180.915 ;
        RECT 237.435 180.900 237.765 180.915 ;
        RECT 231.915 180.600 237.765 180.900 ;
        RECT 231.915 180.585 232.245 180.600 ;
        RECT 237.435 180.585 237.765 180.600 ;
        RECT 215.815 180.220 216.145 180.235 ;
        RECT 213.070 179.920 216.145 180.220 ;
        RECT 185.915 179.905 186.245 179.910 ;
        RECT 173.615 179.565 175.195 179.895 ;
        RECT 162.390 178.910 164.390 179.010 ;
        RECT 161.590 178.860 164.390 178.910 ;
        RECT 167.055 178.860 167.385 178.875 ;
        RECT 161.590 178.560 167.385 178.860 ;
        RECT 191.220 178.860 191.520 179.910 ;
        RECT 215.815 179.905 216.145 179.920 ;
        RECT 192.125 179.565 193.705 179.895 ;
        RECT 210.635 179.565 212.215 179.895 ;
        RECT 229.145 179.565 230.725 179.895 ;
        RECT 208.455 179.540 208.785 179.555 ;
        RECT 209.835 179.540 210.165 179.555 ;
        RECT 208.455 179.240 210.165 179.540 ;
        RECT 208.455 179.225 208.785 179.240 ;
        RECT 209.835 179.225 210.165 179.240 ;
        RECT 212.595 179.540 212.925 179.555 ;
        RECT 213.260 179.540 213.640 179.550 ;
        RECT 212.595 179.240 213.640 179.540 ;
        RECT 212.595 179.225 212.925 179.240 ;
        RECT 213.260 179.230 213.640 179.240 ;
        RECT 223.175 179.540 223.505 179.555 ;
        RECT 224.555 179.540 224.885 179.555 ;
        RECT 223.175 179.240 224.885 179.540 ;
        RECT 223.175 179.225 223.505 179.240 ;
        RECT 224.555 179.225 224.885 179.240 ;
        RECT 211.675 178.860 212.005 178.875 ;
        RECT 216.940 178.860 217.320 178.870 ;
        RECT 222.255 178.860 222.585 178.875 ;
        RECT 191.220 178.560 210.840 178.860 ;
        RECT 161.590 178.510 164.390 178.560 ;
        RECT 167.055 178.545 167.385 178.560 ;
        RECT 162.390 178.410 164.390 178.510 ;
        RECT 188.675 178.180 189.005 178.195 ;
        RECT 188.460 177.865 189.005 178.180 ;
        RECT 190.975 178.180 191.305 178.195 ;
        RECT 199.255 178.180 199.585 178.195 ;
        RECT 207.075 178.180 207.405 178.195 ;
        RECT 190.975 177.880 199.585 178.180 ;
        RECT 190.975 177.865 191.305 177.880 ;
        RECT 199.255 177.865 199.585 177.880 ;
        RECT 200.420 177.880 207.405 178.180 ;
        RECT 210.540 178.180 210.840 178.560 ;
        RECT 211.675 178.560 217.320 178.860 ;
        RECT 211.675 178.545 212.005 178.560 ;
        RECT 216.940 178.550 217.320 178.560 ;
        RECT 219.740 178.560 222.585 178.860 ;
        RECT 217.655 178.180 217.985 178.195 ;
        RECT 210.540 177.880 217.985 178.180 ;
        RECT 182.870 176.845 184.450 177.175 ;
        RECT 188.460 176.835 188.760 177.865 ;
        RECT 189.595 177.500 189.925 177.515 ;
        RECT 197.875 177.500 198.205 177.515 ;
        RECT 189.595 177.200 198.205 177.500 ;
        RECT 189.595 177.185 189.925 177.200 ;
        RECT 197.875 177.185 198.205 177.200 ;
        RECT 181.980 176.510 182.360 176.830 ;
        RECT 188.460 176.520 189.005 176.835 ;
        RECT 200.420 176.820 200.720 177.880 ;
        RECT 207.075 177.865 207.405 177.880 ;
        RECT 217.655 177.865 217.985 177.880 ;
        RECT 219.035 178.180 219.365 178.195 ;
        RECT 219.740 178.180 220.040 178.560 ;
        RECT 222.255 178.545 222.585 178.560 ;
        RECT 219.035 177.880 220.040 178.180 ;
        RECT 220.875 178.180 221.205 178.195 ;
        RECT 233.755 178.180 234.085 178.195 ;
        RECT 220.875 177.880 234.085 178.180 ;
        RECT 219.035 177.865 219.365 177.880 ;
        RECT 220.875 177.865 221.205 177.880 ;
        RECT 233.755 177.865 234.085 177.880 ;
        RECT 207.995 177.500 208.325 177.515 ;
        RECT 215.355 177.500 215.685 177.515 ;
        RECT 217.195 177.500 217.525 177.515 ;
        RECT 207.995 177.200 215.685 177.500 ;
        RECT 207.995 177.185 208.325 177.200 ;
        RECT 215.355 177.185 215.685 177.200 ;
        RECT 216.060 177.200 217.525 177.500 ;
        RECT 201.380 176.845 202.960 177.175 ;
        RECT 174.415 176.140 174.745 176.155 ;
        RECT 175.540 176.140 175.920 176.150 ;
        RECT 174.415 175.840 175.920 176.140 ;
        RECT 182.020 176.140 182.320 176.510 ;
        RECT 188.675 176.505 189.005 176.520 ;
        RECT 192.140 176.520 200.720 176.820 ;
        RECT 207.075 176.820 207.405 176.835 ;
        RECT 216.060 176.820 216.360 177.200 ;
        RECT 217.195 177.185 217.525 177.200 ;
        RECT 222.460 177.500 222.840 177.510 ;
        RECT 228.695 177.500 229.025 177.515 ;
        RECT 222.460 177.200 229.025 177.500 ;
        RECT 222.460 177.190 222.840 177.200 ;
        RECT 228.695 177.185 229.025 177.200 ;
        RECT 229.615 177.500 229.945 177.515 ;
        RECT 235.595 177.500 235.925 177.515 ;
        RECT 229.615 177.200 235.925 177.500 ;
        RECT 229.615 177.185 229.945 177.200 ;
        RECT 235.595 177.185 235.925 177.200 ;
        RECT 219.890 176.845 221.470 177.175 ;
        RECT 238.400 176.845 239.980 177.175 ;
        RECT 207.075 176.520 216.360 176.820 ;
        RECT 224.095 176.820 224.425 176.835 ;
        RECT 234.675 176.820 235.005 176.835 ;
        RECT 224.095 176.520 235.005 176.820 ;
        RECT 192.140 176.140 192.440 176.520 ;
        RECT 207.075 176.505 207.405 176.520 ;
        RECT 224.095 176.505 224.425 176.520 ;
        RECT 234.675 176.505 235.005 176.520 ;
        RECT 182.020 175.840 192.440 176.140 ;
        RECT 212.135 176.140 212.465 176.155 ;
        RECT 215.100 176.140 215.480 176.150 ;
        RECT 212.135 175.840 215.480 176.140 ;
        RECT 174.415 175.825 174.745 175.840 ;
        RECT 175.540 175.830 175.920 175.840 ;
        RECT 212.135 175.825 212.465 175.840 ;
        RECT 215.100 175.830 215.480 175.840 ;
        RECT 218.575 176.140 218.905 176.155 ;
        RECT 232.375 176.140 232.705 176.155 ;
        RECT 218.575 175.840 232.705 176.140 ;
        RECT 218.575 175.825 218.905 175.840 ;
        RECT 232.375 175.825 232.705 175.840 ;
        RECT 190.260 175.460 190.640 175.470 ;
        RECT 192.815 175.460 193.145 175.475 ;
        RECT 190.260 175.160 193.145 175.460 ;
        RECT 190.260 175.150 190.640 175.160 ;
        RECT 192.815 175.145 193.145 175.160 ;
        RECT 218.780 174.780 219.160 174.790 ;
        RECT 236.055 174.780 236.385 174.795 ;
        RECT 218.780 174.480 236.385 174.780 ;
        RECT 218.780 174.470 219.160 174.480 ;
        RECT 236.055 174.465 236.385 174.480 ;
        RECT 246.665 152.705 246.965 217.650 ;
        RECT 247.985 153.875 248.285 219.960 ;
        RECT 249.070 154.925 249.370 220.560 ;
        RECT 249.920 155.950 250.220 221.160 ;
        RECT 250.925 157.080 251.225 224.750 ;
        RECT 251.860 158.175 252.160 225.410 ;
        RECT 251.860 157.875 318.785 158.175 ;
        RECT 250.925 156.780 317.675 157.080 ;
        RECT 249.920 155.650 316.845 155.950 ;
        RECT 249.070 154.625 316.145 154.925 ;
        RECT 247.985 153.575 315.370 153.875 ;
        RECT 246.665 152.405 314.635 152.705 ;
        RECT 198.565 106.260 200.145 106.590 ;
        RECT 235.825 106.260 237.405 106.590 ;
        RECT 273.085 106.260 274.665 106.590 ;
        RECT 310.345 106.260 311.925 106.590 ;
        RECT 181.480 104.875 181.810 104.890 ;
        RECT 186.285 104.875 186.665 104.885 ;
        RECT 181.480 104.575 186.665 104.875 ;
        RECT 181.480 104.560 181.810 104.575 ;
        RECT 186.285 104.565 186.665 104.575 ;
        RECT 179.935 103.540 181.515 103.870 ;
        RECT 217.195 103.540 218.775 103.870 ;
        RECT 254.455 103.540 256.035 103.870 ;
        RECT 291.715 103.540 293.295 103.870 ;
        RECT 190.220 102.835 190.550 102.850 ;
        RECT 249.100 102.835 249.430 102.850 ;
        RECT 190.220 102.535 249.430 102.835 ;
        RECT 190.220 102.520 190.550 102.535 ;
        RECT 249.100 102.520 249.430 102.535 ;
        RECT 237.600 102.155 237.930 102.170 ;
        RECT 238.725 102.155 239.105 102.165 ;
        RECT 237.600 101.855 239.105 102.155 ;
        RECT 237.600 101.840 237.930 101.855 ;
        RECT 238.725 101.845 239.105 101.855 ;
        RECT 314.335 101.625 314.635 152.405 ;
        RECT 174.120 101.485 174.450 101.490 ;
        RECT 229.320 101.485 229.650 101.490 ;
        RECT 259.680 101.485 260.010 101.490 ;
        RECT 277.160 101.485 277.490 101.490 ;
        RECT 174.120 101.475 174.705 101.485 ;
        RECT 229.320 101.475 229.905 101.485 ;
        RECT 259.680 101.475 260.265 101.485 ;
        RECT 174.120 101.175 174.905 101.475 ;
        RECT 229.320 101.175 230.105 101.475 ;
        RECT 259.455 101.175 260.265 101.475 ;
        RECT 174.120 101.165 174.705 101.175 ;
        RECT 229.320 101.165 229.905 101.175 ;
        RECT 259.680 101.165 260.265 101.175 ;
        RECT 277.160 101.475 277.745 101.485 ;
        RECT 277.160 101.175 277.945 101.475 ;
        RECT 277.160 101.165 277.745 101.175 ;
        RECT 174.120 101.160 174.450 101.165 ;
        RECT 229.320 101.160 229.650 101.165 ;
        RECT 259.680 101.160 260.010 101.165 ;
        RECT 277.160 101.160 277.490 101.165 ;
        RECT 198.565 100.820 200.145 101.150 ;
        RECT 235.825 100.820 237.405 101.150 ;
        RECT 273.085 100.820 274.665 101.150 ;
        RECT 310.345 100.820 311.925 101.150 ;
        RECT 312.335 101.025 314.635 101.625 ;
        RECT 239.440 100.795 239.770 100.810 ;
        RECT 255.080 100.795 255.410 100.810 ;
        RECT 239.440 100.495 255.410 100.795 ;
        RECT 239.440 100.480 239.770 100.495 ;
        RECT 255.080 100.480 255.410 100.495 ;
        RECT 256.460 100.795 256.790 100.810 ;
        RECT 261.520 100.795 261.850 100.810 ;
        RECT 256.460 100.495 261.850 100.795 ;
        RECT 256.460 100.480 256.790 100.495 ;
        RECT 261.520 100.480 261.850 100.495 ;
        RECT 283.600 100.795 283.930 100.810 ;
        RECT 287.740 100.795 288.070 100.810 ;
        RECT 283.600 100.495 288.070 100.795 ;
        RECT 283.600 100.480 283.930 100.495 ;
        RECT 287.740 100.480 288.070 100.495 ;
        RECT 198.960 100.115 199.290 100.130 ;
        RECT 208.365 100.115 208.745 100.125 ;
        RECT 223.340 100.115 223.670 100.130 ;
        RECT 289.120 100.115 289.450 100.130 ;
        RECT 198.960 99.815 221.585 100.115 ;
        RECT 198.960 99.800 199.290 99.815 ;
        RECT 208.365 99.805 208.745 99.815 ;
        RECT 205.400 99.435 205.730 99.450 ;
        RECT 220.580 99.435 220.910 99.450 ;
        RECT 205.400 99.135 220.910 99.435 ;
        RECT 205.400 99.120 205.730 99.135 ;
        RECT 220.580 99.120 220.910 99.135 ;
        RECT 221.285 98.755 221.585 99.815 ;
        RECT 223.340 99.815 289.450 100.115 ;
        RECT 223.340 99.800 223.670 99.815 ;
        RECT 289.120 99.800 289.450 99.815 ;
        RECT 309.360 100.115 309.690 100.130 ;
        RECT 312.365 100.115 312.665 101.025 ;
        RECT 309.360 99.815 312.665 100.115 ;
        RECT 309.360 99.800 309.690 99.815 ;
        RECT 248.640 99.435 248.970 99.450 ;
        RECT 303.840 99.435 304.170 99.450 ;
        RECT 248.640 99.135 304.170 99.435 ;
        RECT 248.640 99.120 248.970 99.135 ;
        RECT 303.840 99.120 304.170 99.135 ;
        RECT 241.280 98.755 241.610 98.770 ;
        RECT 221.285 98.455 241.610 98.755 ;
        RECT 241.280 98.440 241.610 98.455 ;
        RECT 260.600 98.755 260.930 98.770 ;
        RECT 279.920 98.755 280.250 98.770 ;
        RECT 260.600 98.455 280.250 98.755 ;
        RECT 260.600 98.440 260.930 98.455 ;
        RECT 279.920 98.440 280.250 98.455 ;
        RECT 179.935 98.100 181.515 98.430 ;
        RECT 217.195 98.100 218.775 98.430 ;
        RECT 254.455 98.100 256.035 98.430 ;
        RECT 291.715 98.100 293.295 98.430 ;
        RECT 220.580 98.075 220.910 98.090 ;
        RECT 252.780 98.075 253.110 98.090 ;
        RECT 220.580 97.775 253.110 98.075 ;
        RECT 220.580 97.760 220.910 97.775 ;
        RECT 252.780 97.760 253.110 97.775 ;
        RECT 257.380 98.075 257.710 98.090 ;
        RECT 263.820 98.075 264.150 98.090 ;
        RECT 257.380 97.775 264.150 98.075 ;
        RECT 257.380 97.760 257.710 97.775 ;
        RECT 263.820 97.760 264.150 97.775 ;
        RECT 186.080 97.395 186.410 97.410 ;
        RECT 198.040 97.395 198.370 97.410 ;
        RECT 186.080 97.095 198.370 97.395 ;
        RECT 186.080 97.080 186.410 97.095 ;
        RECT 198.040 97.080 198.370 97.095 ;
        RECT 219.660 97.395 219.990 97.410 ;
        RECT 228.400 97.395 228.730 97.410 ;
        RECT 219.660 97.095 228.730 97.395 ;
        RECT 219.660 97.080 219.990 97.095 ;
        RECT 228.400 97.080 228.730 97.095 ;
        RECT 234.380 97.395 234.710 97.410 ;
        RECT 237.140 97.395 237.470 97.410 ;
        RECT 246.800 97.395 247.130 97.410 ;
        RECT 260.140 97.395 260.470 97.410 ;
        RECT 261.060 97.405 261.390 97.410 ;
        RECT 234.380 97.095 260.470 97.395 ;
        RECT 234.380 97.080 234.710 97.095 ;
        RECT 237.140 97.080 237.470 97.095 ;
        RECT 246.800 97.080 247.130 97.095 ;
        RECT 260.140 97.080 260.470 97.095 ;
        RECT 260.805 97.395 261.390 97.405 ;
        RECT 283.600 97.395 283.930 97.410 ;
        RECT 285.900 97.395 286.230 97.410 ;
        RECT 260.805 97.095 261.615 97.395 ;
        RECT 283.600 97.095 286.230 97.395 ;
        RECT 260.805 97.085 261.390 97.095 ;
        RECT 261.060 97.080 261.390 97.085 ;
        RECT 283.600 97.080 283.930 97.095 ;
        RECT 285.900 97.080 286.230 97.095 ;
        RECT 177.340 96.715 177.670 96.730 ;
        RECT 238.060 96.715 238.390 96.730 ;
        RECT 177.340 96.415 238.390 96.715 ;
        RECT 177.340 96.400 177.670 96.415 ;
        RECT 238.060 96.400 238.390 96.415 ;
        RECT 241.280 96.715 241.610 96.730 ;
        RECT 280.840 96.715 281.170 96.730 ;
        RECT 299.240 96.715 299.570 96.730 ;
        RECT 241.280 96.415 299.570 96.715 ;
        RECT 241.280 96.400 241.610 96.415 ;
        RECT 280.840 96.400 281.170 96.415 ;
        RECT 299.240 96.400 299.570 96.415 ;
        RECT 203.560 96.035 203.890 96.050 ;
        RECT 254.160 96.035 254.490 96.050 ;
        RECT 262.440 96.035 262.770 96.050 ;
        RECT 203.560 95.735 235.385 96.035 ;
        RECT 203.560 95.720 203.890 95.735 ;
        RECT 198.565 95.380 200.145 95.710 ;
        RECT 208.160 95.355 208.490 95.370 ;
        RECT 210.460 95.355 210.790 95.370 ;
        RECT 231.620 95.355 231.950 95.370 ;
        RECT 208.160 95.055 231.950 95.355 ;
        RECT 208.160 95.040 208.490 95.055 ;
        RECT 210.460 95.040 210.790 95.055 ;
        RECT 231.620 95.040 231.950 95.055 ;
        RECT 235.085 94.690 235.385 95.735 ;
        RECT 254.160 95.735 262.770 96.035 ;
        RECT 254.160 95.720 254.490 95.735 ;
        RECT 262.440 95.720 262.770 95.735 ;
        RECT 235.825 95.380 237.405 95.710 ;
        RECT 273.085 95.380 274.665 95.710 ;
        RECT 310.345 95.380 311.925 95.710 ;
        RECT 244.040 95.355 244.370 95.370 ;
        RECT 259.220 95.355 259.550 95.370 ;
        RECT 262.440 95.355 262.770 95.370 ;
        RECT 244.040 95.055 262.770 95.355 ;
        RECT 244.040 95.040 244.370 95.055 ;
        RECT 259.220 95.040 259.550 95.055 ;
        RECT 262.440 95.040 262.770 95.055 ;
        RECT 218.280 94.675 218.610 94.690 ;
        RECT 221.245 94.675 221.625 94.685 ;
        RECT 218.280 94.375 221.625 94.675 ;
        RECT 218.280 94.360 218.610 94.375 ;
        RECT 221.245 94.365 221.625 94.375 ;
        RECT 222.420 94.675 222.750 94.690 ;
        RECT 227.685 94.675 228.065 94.685 ;
        RECT 222.420 94.375 228.065 94.675 ;
        RECT 235.085 94.375 235.630 94.690 ;
        RECT 222.420 94.360 222.750 94.375 ;
        RECT 227.685 94.365 228.065 94.375 ;
        RECT 235.300 94.360 235.630 94.375 ;
        RECT 238.060 94.675 238.390 94.690 ;
        RECT 260.140 94.675 260.470 94.690 ;
        RECT 238.060 94.375 260.470 94.675 ;
        RECT 238.060 94.360 238.390 94.375 ;
        RECT 260.140 94.360 260.470 94.375 ;
        RECT 263.820 94.675 264.150 94.690 ;
        RECT 278.080 94.675 278.410 94.690 ;
        RECT 263.820 94.375 278.410 94.675 ;
        RECT 263.820 94.360 264.150 94.375 ;
        RECT 278.080 94.360 278.410 94.375 ;
        RECT 204.940 93.995 205.270 94.010 ;
        RECT 210.920 93.995 211.250 94.010 ;
        RECT 246.340 93.995 246.670 94.010 ;
        RECT 204.940 93.695 246.670 93.995 ;
        RECT 204.940 93.680 205.270 93.695 ;
        RECT 210.920 93.680 211.250 93.695 ;
        RECT 246.340 93.680 246.670 93.695 ;
        RECT 159.185 93.315 161.335 93.465 ;
        RECT 163.540 93.315 163.870 93.330 ;
        RECT 159.185 93.015 163.870 93.315 ;
        RECT 159.185 92.865 161.335 93.015 ;
        RECT 163.540 93.000 163.870 93.015 ;
        RECT 224.720 93.315 225.050 93.330 ;
        RECT 242.200 93.315 242.530 93.330 ;
        RECT 224.720 93.015 242.530 93.315 ;
        RECT 224.720 93.000 225.050 93.015 ;
        RECT 242.200 93.000 242.530 93.015 ;
        RECT 179.935 92.660 181.515 92.990 ;
        RECT 217.195 92.660 218.775 92.990 ;
        RECT 254.455 92.660 256.035 92.990 ;
        RECT 291.715 92.660 293.295 92.990 ;
        RECT 221.245 92.635 221.625 92.645 ;
        RECT 244.960 92.635 245.290 92.650 ;
        RECT 221.245 92.335 245.290 92.635 ;
        RECT 221.245 92.325 221.625 92.335 ;
        RECT 244.960 92.320 245.290 92.335 ;
        RECT 177.340 91.955 177.670 91.970 ;
        RECT 242.200 91.955 242.530 91.970 ;
        RECT 177.340 91.655 242.530 91.955 ;
        RECT 177.340 91.640 177.670 91.655 ;
        RECT 242.200 91.640 242.530 91.655 ;
        RECT 220.580 91.275 220.910 91.290 ;
        RECT 224.260 91.275 224.590 91.290 ;
        RECT 291.880 91.275 292.210 91.290 ;
        RECT 220.580 90.975 292.210 91.275 ;
        RECT 220.580 90.960 220.910 90.975 ;
        RECT 224.260 90.960 224.590 90.975 ;
        RECT 291.880 90.960 292.210 90.975 ;
        RECT 198.565 89.940 200.145 90.270 ;
        RECT 235.825 89.940 237.405 90.270 ;
        RECT 273.085 89.940 274.665 90.270 ;
        RECT 310.345 89.940 311.925 90.270 ;
        RECT 245.420 89.915 245.750 89.930 ;
        RECT 245.420 89.615 269.885 89.915 ;
        RECT 245.420 89.600 245.750 89.615 ;
        RECT 208.620 89.235 208.950 89.250 ;
        RECT 263.820 89.235 264.150 89.250 ;
        RECT 208.620 88.935 264.150 89.235 ;
        RECT 269.585 89.235 269.885 89.615 ;
        RECT 285.900 89.235 286.230 89.250 ;
        RECT 269.585 88.935 286.230 89.235 ;
        RECT 208.620 88.920 208.950 88.935 ;
        RECT 263.820 88.920 264.150 88.935 ;
        RECT 285.900 88.920 286.230 88.935 ;
        RECT 175.040 88.555 175.370 88.570 ;
        RECT 265.660 88.555 265.990 88.570 ;
        RECT 175.040 88.255 265.990 88.555 ;
        RECT 175.040 88.240 175.370 88.255 ;
        RECT 265.660 88.240 265.990 88.255 ;
        RECT 237.600 87.875 237.930 87.890 ;
        RECT 239.440 87.875 239.770 87.890 ;
        RECT 237.600 87.575 239.770 87.875 ;
        RECT 237.600 87.560 237.930 87.575 ;
        RECT 239.440 87.560 239.770 87.575 ;
        RECT 260.140 87.875 260.470 87.890 ;
        RECT 260.805 87.875 261.185 87.885 ;
        RECT 260.140 87.575 261.185 87.875 ;
        RECT 260.140 87.560 260.470 87.575 ;
        RECT 260.805 87.565 261.185 87.575 ;
        RECT 179.935 87.220 181.515 87.550 ;
        RECT 217.195 87.220 218.775 87.550 ;
        RECT 254.455 87.220 256.035 87.550 ;
        RECT 291.715 87.220 293.295 87.550 ;
        RECT 208.620 87.205 208.950 87.210 ;
        RECT 208.365 87.195 208.950 87.205 ;
        RECT 222.420 87.195 222.750 87.210 ;
        RECT 238.520 87.195 238.850 87.210 ;
        RECT 208.365 86.895 209.175 87.195 ;
        RECT 222.420 86.895 238.850 87.195 ;
        RECT 208.365 86.885 208.950 86.895 ;
        RECT 208.620 86.880 208.950 86.885 ;
        RECT 222.420 86.880 222.750 86.895 ;
        RECT 238.520 86.880 238.850 86.895 ;
        RECT 186.540 86.515 186.870 86.530 ;
        RECT 262.440 86.515 262.770 86.530 ;
        RECT 186.540 86.215 262.770 86.515 ;
        RECT 186.540 86.200 186.870 86.215 ;
        RECT 262.440 86.200 262.770 86.215 ;
        RECT 310.740 86.515 311.070 86.530 ;
        RECT 310.740 86.215 313.585 86.515 ;
        RECT 310.740 86.200 311.070 86.215 ;
        RECT 220.120 85.835 220.450 85.850 ;
        RECT 228.400 85.835 228.730 85.850 ;
        RECT 240.360 85.835 240.690 85.850 ;
        RECT 220.120 85.535 240.690 85.835 ;
        RECT 220.120 85.520 220.450 85.535 ;
        RECT 228.400 85.520 228.730 85.535 ;
        RECT 240.360 85.520 240.690 85.535 ;
        RECT 313.285 85.305 313.585 86.215 ;
        RECT 240.820 85.155 241.150 85.170 ;
        RECT 253.240 85.155 253.570 85.170 ;
        RECT 240.820 84.855 253.570 85.155 ;
        RECT 240.820 84.840 241.150 84.855 ;
        RECT 253.240 84.840 253.570 84.855 ;
        RECT 312.335 85.145 314.335 85.305 ;
        RECT 315.070 85.145 315.370 153.575 ;
        RECT 312.335 84.845 315.370 85.145 ;
        RECT 198.565 84.500 200.145 84.830 ;
        RECT 235.825 84.500 237.405 84.830 ;
        RECT 273.085 84.500 274.665 84.830 ;
        RECT 310.345 84.500 311.925 84.830 ;
        RECT 312.335 84.705 314.335 84.845 ;
        RECT 242.660 84.475 242.990 84.490 ;
        RECT 244.500 84.475 244.830 84.490 ;
        RECT 260.600 84.475 260.930 84.490 ;
        RECT 242.660 84.175 260.930 84.475 ;
        RECT 242.660 84.160 242.990 84.175 ;
        RECT 244.500 84.160 244.830 84.175 ;
        RECT 260.600 84.160 260.930 84.175 ;
        RECT 207.700 83.795 208.030 83.810 ;
        RECT 226.560 83.795 226.890 83.810 ;
        RECT 276.700 83.795 277.030 83.810 ;
        RECT 207.700 83.495 277.030 83.795 ;
        RECT 207.700 83.480 208.030 83.495 ;
        RECT 226.560 83.480 226.890 83.495 ;
        RECT 276.700 83.480 277.030 83.495 ;
        RECT 192.980 83.115 193.310 83.130 ;
        RECT 202.640 83.115 202.970 83.130 ;
        RECT 256.920 83.115 257.250 83.130 ;
        RECT 192.980 82.815 257.250 83.115 ;
        RECT 192.980 82.800 193.310 82.815 ;
        RECT 202.640 82.800 202.970 82.815 ;
        RECT 256.920 82.800 257.250 82.815 ;
        RECT 261.060 83.115 261.390 83.130 ;
        RECT 281.760 83.115 282.090 83.130 ;
        RECT 261.060 82.815 282.090 83.115 ;
        RECT 261.060 82.800 261.390 82.815 ;
        RECT 281.760 82.800 282.090 82.815 ;
        RECT 221.040 82.435 221.370 82.450 ;
        RECT 227.020 82.435 227.350 82.450 ;
        RECT 242.200 82.435 242.530 82.450 ;
        RECT 221.040 82.135 242.530 82.435 ;
        RECT 221.040 82.120 221.370 82.135 ;
        RECT 227.020 82.120 227.350 82.135 ;
        RECT 242.200 82.120 242.530 82.135 ;
        RECT 244.500 82.435 244.830 82.450 ;
        RECT 249.100 82.435 249.430 82.450 ;
        RECT 244.500 82.135 249.430 82.435 ;
        RECT 244.500 82.120 244.830 82.135 ;
        RECT 249.100 82.120 249.430 82.135 ;
        RECT 179.935 81.780 181.515 82.110 ;
        RECT 217.195 81.780 218.775 82.110 ;
        RECT 254.455 81.780 256.035 82.110 ;
        RECT 291.715 81.780 293.295 82.110 ;
        RECT 233.460 81.755 233.790 81.770 ;
        RECT 241.740 81.755 242.070 81.770 ;
        RECT 252.320 81.755 252.650 81.770 ;
        RECT 233.460 81.455 252.650 81.755 ;
        RECT 233.460 81.440 233.790 81.455 ;
        RECT 241.740 81.440 242.070 81.455 ;
        RECT 252.320 81.440 252.650 81.455 ;
        RECT 256.920 81.755 257.250 81.770 ;
        RECT 259.220 81.755 259.550 81.770 ;
        RECT 256.920 81.455 259.550 81.755 ;
        RECT 256.920 81.440 257.250 81.455 ;
        RECT 259.220 81.440 259.550 81.455 ;
        RECT 213.680 81.075 214.010 81.090 ;
        RECT 238.980 81.075 239.310 81.090 ;
        RECT 289.120 81.075 289.450 81.090 ;
        RECT 293.720 81.075 294.050 81.090 ;
        RECT 213.680 80.775 239.310 81.075 ;
        RECT 213.680 80.760 214.010 80.775 ;
        RECT 238.980 80.760 239.310 80.775 ;
        RECT 283.385 80.775 294.050 81.075 ;
        RECT 177.340 80.395 177.670 80.410 ;
        RECT 200.800 80.395 201.130 80.410 ;
        RECT 177.340 80.095 201.130 80.395 ;
        RECT 177.340 80.080 177.670 80.095 ;
        RECT 200.800 80.080 201.130 80.095 ;
        RECT 216.440 80.395 216.770 80.410 ;
        RECT 229.780 80.395 230.110 80.410 ;
        RECT 216.440 80.095 230.110 80.395 ;
        RECT 216.440 80.080 216.770 80.095 ;
        RECT 229.780 80.080 230.110 80.095 ;
        RECT 198.565 79.060 200.145 79.390 ;
        RECT 235.825 79.060 237.405 79.390 ;
        RECT 238.995 79.035 239.295 80.760 ;
        RECT 256.000 80.395 256.330 80.410 ;
        RECT 283.385 80.395 283.685 80.775 ;
        RECT 289.120 80.760 289.450 80.775 ;
        RECT 293.720 80.760 294.050 80.775 ;
        RECT 256.000 80.095 283.685 80.395 ;
        RECT 256.000 80.080 256.330 80.095 ;
        RECT 245.880 79.725 246.210 79.730 ;
        RECT 245.880 79.715 246.465 79.725 ;
        RECT 245.880 79.415 246.665 79.715 ;
        RECT 245.880 79.405 246.465 79.415 ;
        RECT 245.880 79.400 246.210 79.405 ;
        RECT 273.085 79.060 274.665 79.390 ;
        RECT 310.345 79.060 311.925 79.390 ;
        RECT 239.900 79.035 240.230 79.050 ;
        RECT 238.995 78.735 240.230 79.035 ;
        RECT 239.900 78.720 240.230 78.735 ;
        RECT 256.460 79.035 256.790 79.050 ;
        RECT 259.680 79.035 260.010 79.050 ;
        RECT 256.460 78.735 260.010 79.035 ;
        RECT 256.460 78.720 256.790 78.735 ;
        RECT 259.680 78.720 260.010 78.735 ;
        RECT 177.800 78.355 178.130 78.370 ;
        RECT 213.680 78.355 214.010 78.370 ;
        RECT 177.800 78.055 214.010 78.355 ;
        RECT 177.800 78.040 178.130 78.055 ;
        RECT 213.680 78.040 214.010 78.055 ;
        RECT 223.340 78.355 223.670 78.370 ;
        RECT 301.540 78.355 301.870 78.370 ;
        RECT 223.340 78.055 301.870 78.355 ;
        RECT 223.340 78.040 223.670 78.055 ;
        RECT 301.540 78.040 301.870 78.055 ;
        RECT 219.660 77.675 219.990 77.690 ;
        RECT 275.780 77.675 276.110 77.690 ;
        RECT 219.660 77.375 276.110 77.675 ;
        RECT 219.660 77.360 219.990 77.375 ;
        RECT 275.780 77.360 276.110 77.375 ;
        RECT 220.120 76.995 220.450 77.010 ;
        RECT 233.920 76.995 234.250 77.010 ;
        RECT 220.120 76.695 234.250 76.995 ;
        RECT 220.120 76.680 220.450 76.695 ;
        RECT 233.920 76.680 234.250 76.695 ;
        RECT 237.600 76.995 237.930 77.010 ;
        RECT 247.720 76.995 248.050 77.010 ;
        RECT 237.600 76.695 248.050 76.995 ;
        RECT 237.600 76.680 237.930 76.695 ;
        RECT 247.720 76.680 248.050 76.695 ;
        RECT 258.760 76.995 259.090 77.010 ;
        RECT 260.140 76.995 260.470 77.010 ;
        RECT 264.280 76.995 264.610 77.010 ;
        RECT 258.760 76.695 264.610 76.995 ;
        RECT 258.760 76.680 259.090 76.695 ;
        RECT 260.140 76.680 260.470 76.695 ;
        RECT 264.280 76.680 264.610 76.695 ;
        RECT 179.935 76.340 181.515 76.670 ;
        RECT 217.195 76.340 218.775 76.670 ;
        RECT 254.455 76.340 256.035 76.670 ;
        RECT 291.715 76.340 293.295 76.670 ;
        RECT 236.220 76.315 236.550 76.330 ;
        RECT 242.200 76.315 242.530 76.330 ;
        RECT 236.220 76.015 242.530 76.315 ;
        RECT 236.220 76.000 236.550 76.015 ;
        RECT 242.200 76.000 242.530 76.015 ;
        RECT 231.620 75.635 231.950 75.650 ;
        RECT 179.885 75.335 231.950 75.635 ;
        RECT 179.180 74.955 179.510 74.970 ;
        RECT 179.885 74.955 180.185 75.335 ;
        RECT 231.620 75.320 231.950 75.335 ;
        RECT 179.180 74.655 180.185 74.955 ;
        RECT 184.700 74.955 185.030 74.970 ;
        RECT 194.360 74.955 194.690 74.970 ;
        RECT 257.840 74.955 258.170 74.970 ;
        RECT 259.680 74.955 260.010 74.970 ;
        RECT 276.240 74.955 276.570 74.970 ;
        RECT 184.700 74.655 260.010 74.955 ;
        RECT 179.180 74.640 179.510 74.655 ;
        RECT 184.700 74.640 185.030 74.655 ;
        RECT 194.360 74.640 194.690 74.655 ;
        RECT 257.840 74.640 258.170 74.655 ;
        RECT 259.680 74.640 260.010 74.655 ;
        RECT 269.585 74.655 276.570 74.955 ;
        RECT 220.120 74.275 220.450 74.290 ;
        RECT 221.040 74.275 221.370 74.290 ;
        RECT 227.480 74.275 227.810 74.290 ;
        RECT 269.585 74.275 269.885 74.655 ;
        RECT 276.240 74.640 276.570 74.655 ;
        RECT 220.120 73.975 227.810 74.275 ;
        RECT 220.120 73.960 220.450 73.975 ;
        RECT 221.040 73.960 221.370 73.975 ;
        RECT 227.480 73.960 227.810 73.975 ;
        RECT 269.125 73.975 269.885 74.275 ;
        RECT 198.565 73.620 200.145 73.950 ;
        RECT 235.825 73.620 237.405 73.950 ;
        RECT 219.200 73.595 219.530 73.610 ;
        RECT 225.640 73.595 225.970 73.610 ;
        RECT 259.885 73.595 260.265 73.605 ;
        RECT 269.125 73.595 269.425 73.975 ;
        RECT 273.085 73.620 274.665 73.950 ;
        RECT 310.345 73.620 311.925 73.950 ;
        RECT 219.200 73.295 225.970 73.595 ;
        RECT 219.200 73.280 219.530 73.295 ;
        RECT 225.640 73.280 225.970 73.295 ;
        RECT 255.785 73.295 269.425 73.595 ;
        RECT 175.500 72.915 175.830 72.930 ;
        RECT 214.600 72.915 214.930 72.930 ;
        RECT 234.840 72.915 235.170 72.930 ;
        RECT 255.785 72.915 256.085 73.295 ;
        RECT 259.885 73.285 260.265 73.295 ;
        RECT 175.500 72.615 221.585 72.915 ;
        RECT 175.500 72.600 175.830 72.615 ;
        RECT 214.600 72.600 214.930 72.615 ;
        RECT 202.640 72.235 202.970 72.250 ;
        RECT 221.285 72.235 221.585 72.615 ;
        RECT 234.840 72.615 256.085 72.915 ;
        RECT 234.840 72.600 235.170 72.615 ;
        RECT 232.080 72.235 232.410 72.250 ;
        RECT 202.640 71.935 219.515 72.235 ;
        RECT 221.285 71.935 232.410 72.235 ;
        RECT 202.640 71.920 202.970 71.935 ;
        RECT 195.280 71.555 195.610 71.570 ;
        RECT 201.260 71.555 201.590 71.570 ;
        RECT 195.280 71.255 201.590 71.555 ;
        RECT 219.215 71.555 219.515 71.935 ;
        RECT 232.080 71.920 232.410 71.935 ;
        RECT 246.085 72.235 246.465 72.245 ;
        RECT 246.800 72.235 247.130 72.250 ;
        RECT 246.085 71.935 247.130 72.235 ;
        RECT 246.085 71.925 246.465 71.935 ;
        RECT 246.800 71.920 247.130 71.935 ;
        RECT 253.240 71.555 253.570 71.570 ;
        RECT 219.215 71.255 253.570 71.555 ;
        RECT 195.280 71.240 195.610 71.255 ;
        RECT 201.260 71.240 201.590 71.255 ;
        RECT 253.240 71.240 253.570 71.255 ;
        RECT 179.935 70.900 181.515 71.230 ;
        RECT 217.195 70.900 218.775 71.230 ;
        RECT 254.455 70.900 256.035 71.230 ;
        RECT 291.715 70.900 293.295 71.230 ;
        RECT 183.320 70.875 183.650 70.890 ;
        RECT 203.560 70.875 203.890 70.890 ;
        RECT 232.080 70.875 232.410 70.890 ;
        RECT 250.480 70.875 250.810 70.890 ;
        RECT 183.320 70.575 203.890 70.875 ;
        RECT 183.320 70.560 183.650 70.575 ;
        RECT 203.560 70.560 203.890 70.575 ;
        RECT 219.215 70.575 229.865 70.875 ;
        RECT 199.880 70.195 200.210 70.210 ;
        RECT 219.215 70.195 219.515 70.575 ;
        RECT 229.565 70.205 229.865 70.575 ;
        RECT 232.080 70.575 250.810 70.875 ;
        RECT 232.080 70.560 232.410 70.575 ;
        RECT 250.480 70.560 250.810 70.575 ;
        RECT 199.880 69.895 219.515 70.195 ;
        RECT 229.525 70.195 229.905 70.205 ;
        RECT 256.000 70.195 256.330 70.210 ;
        RECT 277.160 70.205 277.490 70.210 ;
        RECT 277.160 70.195 277.745 70.205 ;
        RECT 284.520 70.195 284.850 70.210 ;
        RECT 229.525 69.895 256.330 70.195 ;
        RECT 276.755 69.895 284.850 70.195 ;
        RECT 199.880 69.880 200.210 69.895 ;
        RECT 229.525 69.885 229.905 69.895 ;
        RECT 256.000 69.880 256.330 69.895 ;
        RECT 277.160 69.885 277.745 69.895 ;
        RECT 277.160 69.880 277.490 69.885 ;
        RECT 284.520 69.880 284.850 69.895 ;
        RECT 310.740 70.195 311.070 70.210 ;
        RECT 310.740 69.895 313.585 70.195 ;
        RECT 310.740 69.880 311.070 69.895 ;
        RECT 228.400 69.515 228.730 69.530 ;
        RECT 271.640 69.515 271.970 69.530 ;
        RECT 228.400 69.215 271.970 69.515 ;
        RECT 228.400 69.200 228.730 69.215 ;
        RECT 271.640 69.200 271.970 69.215 ;
        RECT 313.285 68.985 313.585 69.895 ;
        RECT 239.900 68.835 240.230 68.850 ;
        RECT 241.740 68.835 242.070 68.850 ;
        RECT 239.900 68.535 242.070 68.835 ;
        RECT 239.900 68.520 240.230 68.535 ;
        RECT 241.740 68.520 242.070 68.535 ;
        RECT 312.335 68.820 314.335 68.985 ;
        RECT 315.845 68.820 316.145 154.625 ;
        RECT 312.335 68.520 316.145 68.820 ;
        RECT 198.565 68.180 200.145 68.510 ;
        RECT 235.825 68.180 237.405 68.510 ;
        RECT 273.085 68.180 274.665 68.510 ;
        RECT 310.345 68.180 311.925 68.510 ;
        RECT 312.335 68.385 314.335 68.520 ;
        RECT 226.100 67.475 226.430 67.490 ;
        RECT 297.860 67.475 298.190 67.490 ;
        RECT 226.100 67.175 298.190 67.475 ;
        RECT 226.100 67.160 226.430 67.175 ;
        RECT 297.860 67.160 298.190 67.175 ;
        RECT 180.560 66.795 180.890 66.810 ;
        RECT 220.120 66.795 220.450 66.810 ;
        RECT 236.220 66.795 236.550 66.810 ;
        RECT 180.560 66.495 236.550 66.795 ;
        RECT 180.560 66.480 180.890 66.495 ;
        RECT 220.120 66.480 220.450 66.495 ;
        RECT 236.220 66.480 236.550 66.495 ;
        RECT 256.000 66.795 256.330 66.810 ;
        RECT 259.680 66.795 260.010 66.810 ;
        RECT 256.000 66.495 260.010 66.795 ;
        RECT 256.000 66.480 256.330 66.495 ;
        RECT 259.680 66.480 260.010 66.495 ;
        RECT 226.560 66.115 226.890 66.130 ;
        RECT 242.660 66.115 242.990 66.130 ;
        RECT 226.560 65.815 242.990 66.115 ;
        RECT 226.560 65.800 226.890 65.815 ;
        RECT 242.660 65.800 242.990 65.815 ;
        RECT 179.935 65.460 181.515 65.790 ;
        RECT 217.195 65.460 218.775 65.790 ;
        RECT 254.455 65.460 256.035 65.790 ;
        RECT 291.715 65.460 293.295 65.790 ;
        RECT 248.180 65.435 248.510 65.450 ;
        RECT 219.215 65.135 248.510 65.435 ;
        RECT 212.300 64.755 212.630 64.770 ;
        RECT 219.215 64.755 219.515 65.135 ;
        RECT 248.180 65.120 248.510 65.135 ;
        RECT 212.300 64.455 219.515 64.755 ;
        RECT 247.260 64.755 247.590 64.770 ;
        RECT 255.540 64.755 255.870 64.770 ;
        RECT 296.020 64.755 296.350 64.770 ;
        RECT 247.260 64.455 296.350 64.755 ;
        RECT 212.300 64.440 212.630 64.455 ;
        RECT 247.260 64.440 247.590 64.455 ;
        RECT 255.540 64.440 255.870 64.455 ;
        RECT 296.020 64.440 296.350 64.455 ;
        RECT 213.220 64.075 213.550 64.090 ;
        RECT 221.960 64.075 222.290 64.090 ;
        RECT 213.220 63.775 222.290 64.075 ;
        RECT 213.220 63.760 213.550 63.775 ;
        RECT 221.960 63.760 222.290 63.775 ;
        RECT 231.160 64.075 231.490 64.090 ;
        RECT 254.620 64.075 254.950 64.090 ;
        RECT 258.760 64.075 259.090 64.090 ;
        RECT 231.160 63.775 259.090 64.075 ;
        RECT 231.160 63.760 231.490 63.775 ;
        RECT 254.620 63.760 254.950 63.775 ;
        RECT 258.760 63.760 259.090 63.775 ;
        RECT 210.460 63.395 210.790 63.410 ;
        RECT 221.500 63.395 221.830 63.410 ;
        RECT 210.460 63.095 221.830 63.395 ;
        RECT 210.460 63.080 210.790 63.095 ;
        RECT 221.500 63.080 221.830 63.095 ;
        RECT 198.565 62.740 200.145 63.070 ;
        RECT 235.825 62.740 237.405 63.070 ;
        RECT 273.085 62.740 274.665 63.070 ;
        RECT 310.345 62.740 311.925 63.070 ;
        RECT 174.120 62.725 174.450 62.730 ;
        RECT 174.120 62.715 174.705 62.725 ;
        RECT 174.120 62.415 174.905 62.715 ;
        RECT 174.120 62.405 174.705 62.415 ;
        RECT 174.120 62.400 174.450 62.405 ;
        RECT 227.685 62.035 228.065 62.045 ;
        RECT 235.300 62.035 235.630 62.050 ;
        RECT 227.685 61.735 235.630 62.035 ;
        RECT 227.685 61.725 228.065 61.735 ;
        RECT 235.300 61.720 235.630 61.735 ;
        RECT 215.060 61.355 215.390 61.370 ;
        RECT 284.520 61.355 284.850 61.370 ;
        RECT 215.060 61.055 284.850 61.355 ;
        RECT 215.060 61.040 215.390 61.055 ;
        RECT 284.520 61.040 284.850 61.055 ;
        RECT 159.335 60.675 161.335 60.825 ;
        RECT 164.000 60.675 164.330 60.690 ;
        RECT 158.335 60.375 164.330 60.675 ;
        RECT 159.335 60.225 161.335 60.375 ;
        RECT 164.000 60.360 164.330 60.375 ;
        RECT 179.935 60.020 181.515 60.350 ;
        RECT 217.195 60.020 218.775 60.350 ;
        RECT 254.455 60.020 256.035 60.350 ;
        RECT 291.715 60.020 293.295 60.350 ;
        RECT 231.160 59.315 231.490 59.330 ;
        RECT 241.280 59.315 241.610 59.330 ;
        RECT 231.160 59.015 241.610 59.315 ;
        RECT 231.160 59.000 231.490 59.015 ;
        RECT 241.280 59.000 241.610 59.015 ;
        RECT 174.120 58.635 174.450 58.650 ;
        RECT 247.720 58.635 248.050 58.650 ;
        RECT 174.120 58.335 248.050 58.635 ;
        RECT 174.120 58.320 174.450 58.335 ;
        RECT 247.720 58.320 248.050 58.335 ;
        RECT 198.565 57.300 200.145 57.630 ;
        RECT 235.825 57.300 237.405 57.630 ;
        RECT 273.085 57.300 274.665 57.630 ;
        RECT 310.345 57.300 311.925 57.630 ;
        RECT 230.240 56.595 230.570 56.610 ;
        RECT 266.580 56.595 266.910 56.610 ;
        RECT 230.240 56.295 266.910 56.595 ;
        RECT 230.240 56.280 230.570 56.295 ;
        RECT 266.580 56.280 266.910 56.295 ;
        RECT 186.540 55.925 186.870 55.930 ;
        RECT 186.285 55.915 186.870 55.925 ;
        RECT 250.020 55.915 250.350 55.930 ;
        RECT 185.905 55.615 250.350 55.915 ;
        RECT 186.285 55.605 186.870 55.615 ;
        RECT 186.540 55.600 186.870 55.605 ;
        RECT 250.020 55.600 250.350 55.615 ;
        RECT 224.720 55.235 225.050 55.250 ;
        RECT 242.660 55.235 242.990 55.250 ;
        RECT 224.720 54.935 242.990 55.235 ;
        RECT 224.720 54.920 225.050 54.935 ;
        RECT 242.660 54.920 242.990 54.935 ;
        RECT 179.935 54.580 181.515 54.910 ;
        RECT 217.195 54.580 218.775 54.910 ;
        RECT 254.455 54.580 256.035 54.910 ;
        RECT 291.715 54.580 293.295 54.910 ;
        RECT 310.740 54.555 311.070 54.570 ;
        RECT 310.740 54.255 312.665 54.555 ;
        RECT 310.740 54.240 311.070 54.255 ;
        RECT 233.920 53.875 234.250 53.890 ;
        RECT 281.300 53.875 281.630 53.890 ;
        RECT 233.920 53.575 281.630 53.875 ;
        RECT 233.920 53.560 234.250 53.575 ;
        RECT 281.300 53.560 281.630 53.575 ;
        RECT 174.120 53.195 174.450 53.210 ;
        RECT 178.720 53.195 179.050 53.210 ;
        RECT 240.820 53.195 241.150 53.210 ;
        RECT 174.120 52.895 241.150 53.195 ;
        RECT 174.120 52.880 174.450 52.895 ;
        RECT 178.720 52.880 179.050 52.895 ;
        RECT 240.820 52.880 241.150 52.895 ;
        RECT 312.365 52.665 312.665 54.255 ;
        RECT 312.335 52.505 314.335 52.665 ;
        RECT 316.545 52.505 316.845 155.650 ;
        RECT 312.335 52.205 316.845 52.505 ;
        RECT 198.565 51.860 200.145 52.190 ;
        RECT 235.825 51.860 237.405 52.190 ;
        RECT 273.085 51.860 274.665 52.190 ;
        RECT 310.345 51.860 311.925 52.190 ;
        RECT 312.335 52.065 314.335 52.205 ;
        RECT 179.935 49.140 181.515 49.470 ;
        RECT 217.195 49.140 218.775 49.470 ;
        RECT 254.455 49.140 256.035 49.470 ;
        RECT 291.715 49.140 293.295 49.470 ;
        RECT 269.800 49.115 270.130 49.130 ;
        RECT 281.760 49.115 282.090 49.130 ;
        RECT 269.800 48.815 282.090 49.115 ;
        RECT 269.800 48.800 270.130 48.815 ;
        RECT 281.760 48.800 282.090 48.815 ;
        RECT 269.800 47.755 270.130 47.770 ;
        RECT 277.160 47.755 277.490 47.770 ;
        RECT 269.800 47.455 277.490 47.755 ;
        RECT 269.800 47.440 270.130 47.455 ;
        RECT 277.160 47.440 277.490 47.455 ;
        RECT 198.565 46.420 200.145 46.750 ;
        RECT 235.825 46.420 237.405 46.750 ;
        RECT 273.085 46.420 274.665 46.750 ;
        RECT 310.345 46.420 311.925 46.750 ;
        RECT 269.340 45.715 269.670 45.730 ;
        RECT 278.080 45.715 278.410 45.730 ;
        RECT 269.340 45.415 278.410 45.715 ;
        RECT 269.340 45.400 269.670 45.415 ;
        RECT 278.080 45.400 278.410 45.415 ;
        RECT 179.935 43.700 181.515 44.030 ;
        RECT 217.195 43.700 218.775 44.030 ;
        RECT 254.455 43.700 256.035 44.030 ;
        RECT 291.715 43.700 293.295 44.030 ;
        RECT 198.565 40.980 200.145 41.310 ;
        RECT 235.825 40.980 237.405 41.310 ;
        RECT 273.085 40.980 274.665 41.310 ;
        RECT 310.345 40.980 311.925 41.310 ;
        RECT 238.520 38.925 238.850 38.930 ;
        RECT 238.520 38.915 239.105 38.925 ;
        RECT 238.295 38.615 239.105 38.915 ;
        RECT 238.520 38.605 239.105 38.615 ;
        RECT 238.520 38.600 238.850 38.605 ;
        RECT 179.935 38.260 181.515 38.590 ;
        RECT 217.195 38.260 218.775 38.590 ;
        RECT 254.455 38.260 256.035 38.590 ;
        RECT 291.715 38.260 293.295 38.590 ;
        RECT 238.520 36.875 238.850 36.890 ;
        RECT 296.940 36.875 297.270 36.890 ;
        RECT 238.520 36.575 297.270 36.875 ;
        RECT 238.520 36.560 238.850 36.575 ;
        RECT 296.940 36.560 297.270 36.575 ;
        RECT 316.555 36.345 316.955 36.545 ;
        RECT 198.565 35.540 200.145 35.870 ;
        RECT 235.825 35.540 237.405 35.870 ;
        RECT 273.085 35.540 274.665 35.870 ;
        RECT 310.345 35.540 311.925 35.870 ;
        RECT 312.335 35.745 316.955 36.345 ;
        RECT 270.720 34.835 271.050 34.850 ;
        RECT 294.640 34.835 294.970 34.850 ;
        RECT 270.720 34.535 294.970 34.835 ;
        RECT 270.720 34.520 271.050 34.535 ;
        RECT 294.640 34.520 294.970 34.535 ;
        RECT 300.160 34.835 300.490 34.850 ;
        RECT 312.365 34.835 312.665 35.745 ;
        RECT 300.160 34.535 312.665 34.835 ;
        RECT 300.160 34.520 300.490 34.535 ;
        RECT 179.935 32.820 181.515 33.150 ;
        RECT 217.195 32.820 218.775 33.150 ;
        RECT 254.455 32.820 256.035 33.150 ;
        RECT 291.715 32.820 293.295 33.150 ;
        RECT 233.460 31.435 233.790 31.450 ;
        RECT 236.220 31.435 236.550 31.450 ;
        RECT 233.460 31.135 236.550 31.435 ;
        RECT 233.460 31.120 233.790 31.135 ;
        RECT 236.220 31.120 236.550 31.135 ;
        RECT 198.565 30.100 200.145 30.430 ;
        RECT 235.825 30.100 237.405 30.430 ;
        RECT 273.085 30.100 274.665 30.430 ;
        RECT 310.345 30.100 311.925 30.430 ;
        RECT 159.335 28.035 161.335 28.185 ;
        RECT 164.000 28.035 164.330 28.050 ;
        RECT 157.560 27.735 164.330 28.035 ;
        RECT 159.335 27.585 161.335 27.735 ;
        RECT 164.000 27.720 164.330 27.735 ;
        RECT 179.935 27.380 181.515 27.710 ;
        RECT 217.195 27.380 218.775 27.710 ;
        RECT 254.455 27.380 256.035 27.710 ;
        RECT 291.715 27.380 293.295 27.710 ;
        RECT 198.565 24.660 200.145 24.990 ;
        RECT 235.825 24.660 237.405 24.990 ;
        RECT 273.085 24.660 274.665 24.990 ;
        RECT 310.345 24.660 311.925 24.990 ;
        RECT 179.935 21.940 181.515 22.270 ;
        RECT 217.195 21.940 218.775 22.270 ;
        RECT 254.455 21.940 256.035 22.270 ;
        RECT 291.715 21.940 293.295 22.270 ;
        RECT 276.485 20.935 313.585 21.235 ;
        RECT 248.640 20.555 248.970 20.570 ;
        RECT 276.485 20.555 276.785 20.935 ;
        RECT 248.640 20.255 276.785 20.555 ;
        RECT 248.640 20.240 248.970 20.255 ;
        RECT 313.285 20.025 313.585 20.935 ;
        RECT 312.335 19.845 314.335 20.025 ;
        RECT 317.375 19.845 317.675 156.780 ;
        RECT 318.485 36.545 318.785 157.875 ;
        RECT 318.085 35.745 318.785 36.545 ;
        RECT 198.565 19.220 200.145 19.550 ;
        RECT 235.825 19.220 237.405 19.550 ;
        RECT 273.085 19.220 274.665 19.550 ;
        RECT 310.345 19.220 311.925 19.550 ;
        RECT 312.335 19.545 317.675 19.845 ;
        RECT 312.335 19.425 314.335 19.545 ;
        RECT 179.935 16.500 181.515 16.830 ;
        RECT 217.195 16.500 218.775 16.830 ;
        RECT 254.455 16.500 256.035 16.830 ;
        RECT 291.715 16.500 293.295 16.830 ;
        RECT 198.565 13.780 200.145 14.110 ;
        RECT 235.825 13.780 237.405 14.110 ;
        RECT 273.085 13.780 274.665 14.110 ;
        RECT 310.345 13.780 311.925 14.110 ;
      LAYER met4 ;
        RECT 23.260 224.760 23.310 225.560 ;
        RECT 23.610 224.760 23.660 225.560 ;
        RECT 45.340 224.760 45.390 225.560 ;
        RECT 45.690 224.760 45.740 225.560 ;
        RECT 65.010 225.310 65.510 225.710 ;
        RECT 125.730 225.360 126.530 225.760 ;
        RECT 59.490 224.760 59.990 225.160 ;
        RECT 67.770 224.760 68.270 225.110 ;
        RECT 129.395 225.050 130.195 225.100 ;
        RECT 75.700 224.760 75.750 224.860 ;
        RECT 76.050 224.760 76.100 224.860 ;
        RECT 78.810 224.760 78.945 224.860 ;
        RECT 15.030 224.460 15.330 224.760 ;
        RECT 17.790 224.460 18.090 224.760 ;
        RECT 20.550 224.460 20.850 224.760 ;
        RECT 26.070 224.460 26.370 224.760 ;
        RECT 28.830 224.460 29.130 224.760 ;
        RECT 31.590 224.460 31.890 224.760 ;
        RECT 34.350 224.460 34.650 224.760 ;
        RECT 37.110 224.460 37.410 224.760 ;
        RECT 39.870 224.460 40.170 224.760 ;
        RECT 42.630 224.460 42.930 224.760 ;
        RECT 48.150 224.460 48.450 224.760 ;
        RECT 50.910 224.460 51.210 224.760 ;
        RECT 53.670 224.460 53.970 224.760 ;
        RECT 56.430 224.460 56.730 224.760 ;
        RECT 3.600 224.060 56.730 224.460 ;
        RECT 61.950 224.560 62.250 224.760 ;
        RECT 67.470 224.710 68.270 224.760 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.510 70.530 224.760 ;
        RECT 70.230 224.110 71.030 224.510 ;
        RECT 1.000 220.760 1.800 221.560 ;
        RECT 3.600 220.760 5.200 224.060 ;
        RECT 72.990 223.910 73.290 224.760 ;
        RECT 75.700 224.060 76.100 224.760 ;
        RECT 78.510 224.060 78.945 224.760 ;
        RECT 83.980 224.760 84.030 224.860 ;
        RECT 84.330 224.760 84.380 224.860 ;
        RECT 83.980 224.060 84.380 224.760 ;
        RECT 86.740 224.760 86.790 224.860 ;
        RECT 87.090 224.760 87.140 224.860 ;
        RECT 86.740 224.060 87.140 224.760 ;
        RECT 92.260 224.760 92.310 224.860 ;
        RECT 92.610 224.760 92.660 224.860 ;
        RECT 128.490 224.760 130.195 225.050 ;
        RECT 92.260 224.060 92.660 224.760 ;
        RECT 95.070 224.450 95.370 224.760 ;
        RECT 97.830 224.450 98.130 224.760 ;
        RECT 100.590 224.450 100.890 224.760 ;
        RECT 103.350 224.450 103.650 224.760 ;
        RECT 106.110 224.450 106.410 224.760 ;
        RECT 108.870 224.615 109.170 224.760 ;
        RECT 72.990 223.510 73.790 223.910 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.650 106.460 224.450 ;
        RECT 108.865 224.215 109.665 224.615 ;
        RECT 6.200 221.180 109.540 222.780 ;
        RECT 111.630 221.515 111.930 224.760 ;
        RECT 114.390 222.115 114.690 224.760 ;
        RECT 117.150 222.715 117.450 224.760 ;
        RECT 119.910 223.315 120.210 224.760 ;
        RECT 122.670 223.915 122.970 224.760 ;
        RECT 128.190 224.750 130.195 224.760 ;
        RECT 129.395 224.700 130.195 224.750 ;
        RECT 122.670 223.615 149.190 223.915 ;
        RECT 119.910 223.015 145.160 223.315 ;
        RECT 117.150 222.415 141.130 222.715 ;
        RECT 114.390 221.815 137.100 222.115 ;
        RECT 136.800 221.515 137.100 221.815 ;
        RECT 140.830 221.515 141.130 222.415 ;
        RECT 144.860 221.515 145.160 223.015 ;
        RECT 148.890 221.515 149.190 223.615 ;
      LAYER met4 ;
        RECT 255.465 221.585 317.065 223.185 ;
      LAYER met4 ;
        RECT 111.630 221.215 133.120 221.515 ;
        RECT 6.200 220.760 7.800 221.180 ;
        RECT 10.550 218.590 105.040 220.190 ;
        RECT 7.800 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 103.440 211.240 105.040 218.590 ;
        RECT 106.340 219.305 109.540 221.180 ;
        RECT 132.720 220.715 133.120 221.215 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 106.340 217.705 151.230 219.305 ;
        RECT 106.340 217.515 109.540 217.705 ;
        RECT 106.415 211.240 108.015 213.740 ;
        RECT 150.830 211.240 248.550 212.040 ;
        RECT 27.080 209.940 53.660 210.740 ;
        RECT 27.080 209.640 27.570 209.940 ;
        RECT 16.115 199.365 25.725 208.975 ;
        RECT 16.115 196.975 16.715 199.365 ;
        RECT 16.115 187.365 25.725 196.975 ;
        RECT 16.115 184.975 16.715 187.365 ;
        RECT 16.115 175.365 25.725 184.975 ;
        RECT 16.115 172.975 16.715 175.365 ;
        RECT 16.115 163.365 25.725 172.975 ;
        RECT 16.115 160.975 16.715 163.365 ;
        RECT 16.115 151.365 25.725 160.975 ;
        RECT 16.115 150.210 16.715 151.365 ;
        RECT 27.080 150.970 27.565 209.640 ;
        RECT 28.915 199.365 38.525 208.975 ;
        RECT 37.925 196.975 38.525 199.365 ;
        RECT 28.915 187.365 38.525 196.975 ;
        RECT 52.860 188.465 53.660 209.940 ;
        RECT 103.440 209.640 248.550 211.240 ;
        RECT 150.830 208.840 248.550 209.640 ;
        RECT 110.530 187.540 156.765 189.140 ;
        RECT 37.925 184.975 38.525 187.365 ;
        RECT 28.915 175.365 38.525 184.975 ;
        RECT 37.925 172.975 38.525 175.365 ;
        RECT 28.915 163.365 38.525 172.975 ;
        RECT 51.950 184.940 103.750 186.540 ;
        RECT 51.950 169.890 53.550 184.940 ;
        RECT 57.020 177.390 109.070 178.990 ;
        RECT 153.565 178.210 156.765 187.540 ;
        RECT 151.155 175.010 156.765 178.210 ;
        RECT 173.605 176.770 175.205 208.840 ;
        RECT 175.565 189.425 175.895 189.755 ;
        RECT 175.580 176.155 175.880 189.425 ;
        RECT 182.005 188.745 182.335 189.075 ;
        RECT 182.020 176.835 182.320 188.745 ;
        RECT 182.005 176.505 182.335 176.835 ;
        RECT 175.565 175.825 175.895 176.155 ;
        RECT 51.950 168.290 58.420 169.890 ;
        RECT 37.925 160.975 38.525 163.365 ;
        RECT 28.915 151.365 38.525 160.975 ;
        RECT 153.565 168.200 156.765 175.010 ;
        RECT 182.860 168.200 184.460 201.730 ;
        RECT 191.205 194.865 191.535 195.195 ;
        RECT 187.525 189.425 187.855 189.755 ;
        RECT 185.685 185.345 186.015 185.675 ;
        RECT 184.765 184.665 185.095 184.995 ;
        RECT 184.780 180.235 185.080 184.665 ;
        RECT 185.700 180.235 186.000 185.345 ;
        RECT 187.540 184.995 187.840 189.425 ;
        RECT 190.285 188.065 190.615 188.395 ;
        RECT 187.525 184.665 187.855 184.995 ;
        RECT 184.765 179.905 185.095 180.235 ;
        RECT 185.685 179.905 186.015 180.235 ;
        RECT 190.300 175.475 190.600 188.065 ;
        RECT 191.220 180.235 191.520 194.865 ;
        RECT 191.205 179.905 191.535 180.235 ;
        RECT 192.115 176.770 193.715 208.840 ;
        RECT 190.285 175.145 190.615 175.475 ;
        RECT 201.370 168.200 202.970 201.730 ;
        RECT 210.625 176.770 212.225 208.840 ;
        RECT 216.965 189.425 217.295 189.755 ;
        RECT 213.285 186.705 213.615 187.035 ;
        RECT 213.300 179.555 213.600 186.705 ;
        RECT 215.125 182.625 215.455 182.955 ;
        RECT 213.285 179.225 213.615 179.555 ;
        RECT 215.140 176.155 215.440 182.625 ;
        RECT 216.980 178.875 217.280 189.425 ;
        RECT 218.805 188.745 219.135 189.075 ;
        RECT 216.965 178.545 217.295 178.875 ;
        RECT 215.125 175.825 215.455 176.155 ;
        RECT 218.820 174.795 219.120 188.745 ;
        RECT 218.805 174.465 219.135 174.795 ;
        RECT 219.880 168.200 221.480 201.730 ;
        RECT 222.485 183.305 222.815 183.635 ;
        RECT 222.500 177.515 222.800 183.305 ;
        RECT 222.485 177.185 222.815 177.515 ;
        RECT 229.135 176.770 230.735 208.840 ;
        RECT 238.390 168.200 239.990 201.730 ;
        RECT 153.565 165.000 240.760 168.200 ;
        RECT 111.685 158.165 112.085 158.565 ;
        RECT 105.385 157.765 112.085 158.165 ;
        RECT 105.385 157.365 105.785 157.765 ;
        RECT 109.415 156.565 109.815 156.965 ;
        RECT 113.085 156.565 113.485 156.965 ;
        RECT 109.415 156.165 113.485 156.565 ;
        RECT 37.925 150.210 38.525 151.365 ;
        RECT 16.115 149.410 46.630 150.210 ;
        RECT 51.575 145.090 73.495 148.290 ;
        RECT 9.490 135.030 17.100 142.640 ;
        RECT 18.455 142.175 20.750 142.975 ;
        RECT 13.385 130.025 14.185 135.030 ;
        RECT 18.455 134.695 18.935 142.175 ;
        RECT 20.350 141.375 20.750 142.175 ;
        RECT 61.980 135.495 62.780 135.895 ;
        RECT 61.980 135.095 140.370 135.495 ;
        RECT 22.615 133.320 80.925 134.120 ;
        RECT 20.650 131.810 21.050 132.210 ;
        RECT 137.945 131.810 138.345 132.210 ;
        RECT 20.650 131.410 138.345 131.810 ;
        RECT 139.120 130.025 139.520 132.990 ;
        RECT 13.385 129.625 139.520 130.025 ;
        RECT 16.805 128.710 139.520 129.110 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 128.710 ;
        RECT 139.970 125.690 140.370 135.095 ;
        RECT 140.940 131.390 142.100 132.990 ;
        RECT 140.940 125.060 141.340 131.390 ;
        RECT 131.145 124.660 141.340 125.060 ;
        RECT 103.315 121.565 118.965 123.165 ;
        RECT 109.865 107.965 118.715 109.565 ;
        RECT 63.315 103.465 74.365 105.065 ;
        RECT 105.965 103.615 118.565 105.215 ;
        RECT 131.145 98.015 131.545 124.660 ;
        RECT 153.565 124.090 156.765 165.000 ;
        RECT 142.760 122.490 156.765 124.090 ;
        RECT 153.565 114.150 156.765 122.490 ;
        RECT 139.355 113.350 156.765 114.150 ;
        RECT 245.350 113.705 248.550 208.840 ;
      LAYER met4 ;
        RECT 255.465 207.185 257.065 221.585 ;
      LAYER met4 ;
        RECT 257.065 219.185 271.465 221.585 ;
      LAYER met4 ;
        RECT 271.465 219.585 277.065 221.585 ;
      LAYER met4 ;
        RECT 277.065 219.585 279.465 221.585 ;
      LAYER met4 ;
        RECT 279.465 219.585 285.065 221.585 ;
      LAYER met4 ;
        RECT 285.065 219.585 289.465 221.585 ;
      LAYER met4 ;
        RECT 289.465 219.585 293.065 221.585 ;
      LAYER met4 ;
        RECT 293.065 219.585 297.465 221.585 ;
      LAYER met4 ;
        RECT 297.465 219.585 301.065 221.585 ;
      LAYER met4 ;
        RECT 257.065 209.585 259.465 219.185 ;
      LAYER met4 ;
        RECT 259.465 217.585 269.065 219.185 ;
        RECT 259.465 211.185 261.065 217.585 ;
      LAYER met4 ;
        RECT 261.065 211.185 267.465 217.585 ;
      LAYER met4 ;
        RECT 267.465 211.185 269.065 217.585 ;
        RECT 259.465 209.585 269.065 211.185 ;
      LAYER met4 ;
        RECT 269.065 209.585 271.465 219.185 ;
      LAYER met4 ;
        RECT 271.465 215.185 273.065 219.585 ;
      LAYER met4 ;
        RECT 273.065 217.185 279.465 219.585 ;
      LAYER met4 ;
        RECT 279.465 217.185 283.065 219.585 ;
      LAYER met4 ;
        RECT 283.065 217.185 289.465 219.585 ;
      LAYER met4 ;
        RECT 289.465 217.185 291.065 219.585 ;
      LAYER met4 ;
        RECT 291.065 219.185 299.465 219.585 ;
        RECT 291.065 217.585 295.465 219.185 ;
      LAYER met4 ;
        RECT 295.465 217.585 297.065 219.185 ;
      LAYER met4 ;
        RECT 297.065 217.585 299.465 219.185 ;
        RECT 291.065 217.185 299.465 217.585 ;
        RECT 273.065 215.585 275.465 217.185 ;
      LAYER met4 ;
        RECT 275.465 215.585 291.065 217.185 ;
      LAYER met4 ;
        RECT 291.065 215.585 293.465 217.185 ;
      LAYER met4 ;
        RECT 293.465 215.585 295.065 217.185 ;
      LAYER met4 ;
        RECT 295.065 215.585 299.465 217.185 ;
        RECT 273.065 215.185 277.465 215.585 ;
      LAYER met4 ;
        RECT 271.465 213.585 275.065 215.185 ;
      LAYER met4 ;
        RECT 275.065 213.585 277.465 215.185 ;
      LAYER met4 ;
        RECT 277.465 213.585 281.065 215.585 ;
      LAYER met4 ;
        RECT 281.065 213.585 285.465 215.585 ;
      LAYER met4 ;
        RECT 285.465 213.585 287.065 215.585 ;
      LAYER met4 ;
        RECT 287.065 213.585 289.465 215.585 ;
      LAYER met4 ;
        RECT 289.465 215.185 291.065 215.585 ;
      LAYER met4 ;
        RECT 291.065 215.185 299.465 215.585 ;
      LAYER met4 ;
        RECT 289.465 213.585 293.065 215.185 ;
      LAYER met4 ;
        RECT 293.065 213.585 299.465 215.185 ;
        RECT 257.065 207.185 271.465 209.585 ;
      LAYER met4 ;
        RECT 271.465 207.185 273.065 213.585 ;
      LAYER met4 ;
        RECT 273.065 211.185 279.465 213.585 ;
      LAYER met4 ;
        RECT 255.465 205.585 273.065 207.185 ;
      LAYER met4 ;
        RECT 273.065 205.585 275.465 211.185 ;
      LAYER met4 ;
        RECT 255.465 199.185 257.065 205.585 ;
      LAYER met4 ;
        RECT 257.065 201.585 261.465 205.585 ;
      LAYER met4 ;
        RECT 261.465 203.185 263.065 205.585 ;
      LAYER met4 ;
        RECT 263.065 203.185 265.465 205.585 ;
      LAYER met4 ;
        RECT 265.465 203.585 269.065 205.585 ;
      LAYER met4 ;
        RECT 269.065 205.185 275.465 205.585 ;
      LAYER met4 ;
        RECT 275.465 205.185 277.065 211.185 ;
      LAYER met4 ;
        RECT 277.065 207.585 279.465 211.185 ;
      LAYER met4 ;
        RECT 279.465 207.585 281.065 213.585 ;
      LAYER met4 ;
        RECT 281.065 213.185 299.465 213.585 ;
      LAYER met4 ;
        RECT 299.465 213.185 301.065 219.585 ;
      LAYER met4 ;
        RECT 301.065 219.185 315.465 221.585 ;
        RECT 281.065 207.585 283.465 213.185 ;
      LAYER met4 ;
        RECT 283.465 211.185 285.065 213.185 ;
      LAYER met4 ;
        RECT 285.065 211.585 295.465 213.185 ;
      LAYER met4 ;
        RECT 295.465 211.585 301.065 213.185 ;
      LAYER met4 ;
        RECT 285.065 211.185 297.465 211.585 ;
      LAYER met4 ;
        RECT 283.465 209.585 287.065 211.185 ;
      LAYER met4 ;
        RECT 287.065 209.585 289.465 211.185 ;
      LAYER met4 ;
        RECT 289.465 209.585 295.065 211.185 ;
      LAYER met4 ;
        RECT 295.065 209.585 297.465 211.185 ;
      LAYER met4 ;
        RECT 297.465 209.585 301.065 211.585 ;
      LAYER met4 ;
        RECT 301.065 209.585 303.465 219.185 ;
      LAYER met4 ;
        RECT 303.465 217.585 313.065 219.185 ;
        RECT 303.465 211.185 305.065 217.585 ;
      LAYER met4 ;
        RECT 305.065 211.185 311.465 217.585 ;
      LAYER met4 ;
        RECT 311.465 211.185 313.065 217.585 ;
        RECT 303.465 209.585 313.065 211.185 ;
      LAYER met4 ;
        RECT 313.065 209.585 315.465 219.185 ;
      LAYER met4 ;
        RECT 283.465 207.585 285.065 209.585 ;
      LAYER met4 ;
        RECT 285.065 209.185 291.465 209.585 ;
        RECT 285.065 207.585 287.465 209.185 ;
        RECT 277.065 207.185 287.465 207.585 ;
      LAYER met4 ;
        RECT 287.465 207.185 289.065 209.185 ;
      LAYER met4 ;
        RECT 289.065 207.585 291.465 209.185 ;
      LAYER met4 ;
        RECT 291.465 207.585 293.065 209.585 ;
      LAYER met4 ;
        RECT 293.065 209.185 299.465 209.585 ;
        RECT 293.065 207.585 295.465 209.185 ;
        RECT 277.065 205.585 281.465 207.185 ;
      LAYER met4 ;
        RECT 281.465 205.585 283.065 207.185 ;
      LAYER met4 ;
        RECT 283.065 205.585 285.465 207.185 ;
      LAYER met4 ;
        RECT 285.465 205.585 289.065 207.185 ;
      LAYER met4 ;
        RECT 289.065 205.585 295.465 207.585 ;
      LAYER met4 ;
        RECT 295.465 205.585 297.065 209.185 ;
      LAYER met4 ;
        RECT 297.065 205.585 299.465 209.185 ;
      LAYER met4 ;
        RECT 299.465 207.185 301.065 209.585 ;
      LAYER met4 ;
        RECT 301.065 207.185 315.465 209.585 ;
      LAYER met4 ;
        RECT 315.465 207.185 317.065 221.585 ;
        RECT 299.465 205.585 317.065 207.185 ;
      LAYER met4 ;
        RECT 277.065 205.185 287.465 205.585 ;
      LAYER met4 ;
        RECT 287.465 205.185 289.065 205.585 ;
      LAYER met4 ;
        RECT 289.065 205.185 299.465 205.585 ;
      LAYER met4 ;
        RECT 299.465 205.185 301.065 205.585 ;
      LAYER met4 ;
        RECT 269.065 203.585 273.465 205.185 ;
      LAYER met4 ;
        RECT 273.465 203.585 279.065 205.185 ;
      LAYER met4 ;
        RECT 279.065 203.585 283.465 205.185 ;
      LAYER met4 ;
        RECT 283.465 203.585 285.065 205.185 ;
      LAYER met4 ;
        RECT 285.065 203.585 287.465 205.185 ;
      LAYER met4 ;
        RECT 287.465 203.585 295.065 205.185 ;
      LAYER met4 ;
        RECT 295.065 203.585 297.465 205.185 ;
      LAYER met4 ;
        RECT 297.465 203.585 301.065 205.185 ;
      LAYER met4 ;
        RECT 301.065 203.585 307.465 205.585 ;
      LAYER met4 ;
        RECT 307.465 203.585 309.065 205.585 ;
      LAYER met4 ;
        RECT 309.065 203.585 313.465 205.585 ;
      LAYER met4 ;
        RECT 313.465 203.585 317.065 205.585 ;
        RECT 265.465 203.185 267.065 203.585 ;
      LAYER met4 ;
        RECT 267.065 203.185 277.465 203.585 ;
      LAYER met4 ;
        RECT 261.465 201.585 267.065 203.185 ;
      LAYER met4 ;
        RECT 267.065 201.585 269.465 203.185 ;
      LAYER met4 ;
        RECT 269.465 201.585 271.065 203.185 ;
      LAYER met4 ;
        RECT 271.065 201.585 277.465 203.185 ;
        RECT 257.065 201.185 277.465 201.585 ;
      LAYER met4 ;
        RECT 277.465 201.185 279.065 203.585 ;
      LAYER met4 ;
        RECT 279.065 203.185 287.465 203.585 ;
      LAYER met4 ;
        RECT 287.465 203.185 289.065 203.585 ;
      LAYER met4 ;
        RECT 289.065 203.185 297.465 203.585 ;
      LAYER met4 ;
        RECT 297.465 203.185 299.065 203.585 ;
      LAYER met4 ;
        RECT 299.065 203.185 315.465 203.585 ;
        RECT 279.065 201.585 285.465 203.185 ;
      LAYER met4 ;
        RECT 285.465 201.585 289.065 203.185 ;
      LAYER met4 ;
        RECT 289.065 201.585 295.465 203.185 ;
      LAYER met4 ;
        RECT 295.465 201.585 299.065 203.185 ;
      LAYER met4 ;
        RECT 299.065 201.585 303.465 203.185 ;
      LAYER met4 ;
        RECT 303.465 201.585 307.065 203.185 ;
      LAYER met4 ;
        RECT 257.065 199.185 271.465 201.185 ;
      LAYER met4 ;
        RECT 271.465 199.185 273.065 201.185 ;
      LAYER met4 ;
        RECT 273.065 199.585 275.465 201.185 ;
      LAYER met4 ;
        RECT 275.465 199.585 279.065 201.185 ;
      LAYER met4 ;
        RECT 279.065 199.585 287.465 201.585 ;
      LAYER met4 ;
        RECT 287.465 201.185 289.065 201.585 ;
      LAYER met4 ;
        RECT 289.065 201.185 305.465 201.585 ;
      LAYER met4 ;
        RECT 287.465 199.585 291.065 201.185 ;
      LAYER met4 ;
        RECT 291.065 199.585 299.465 201.185 ;
      LAYER met4 ;
        RECT 299.465 199.585 301.065 201.185 ;
      LAYER met4 ;
        RECT 301.065 199.585 305.465 201.185 ;
        RECT 273.065 199.185 287.465 199.585 ;
      LAYER met4 ;
        RECT 287.465 199.185 289.065 199.585 ;
      LAYER met4 ;
        RECT 289.065 199.185 305.465 199.585 ;
      LAYER met4 ;
        RECT 305.465 199.185 307.065 201.585 ;
      LAYER met4 ;
        RECT 307.065 201.185 315.465 203.185 ;
      LAYER met4 ;
        RECT 315.465 201.185 317.065 203.585 ;
      LAYER met4 ;
        RECT 307.065 199.185 313.465 201.185 ;
      LAYER met4 ;
        RECT 255.465 195.185 259.065 199.185 ;
      LAYER met4 ;
        RECT 259.065 197.585 261.465 199.185 ;
        POLYGON 261.465 199.185 261.770 199.185 261.465 198.880 ;
      LAYER met4 ;
        RECT 261.770 198.880 273.065 199.185 ;
        RECT 261.465 197.585 273.065 198.880 ;
      LAYER met4 ;
        RECT 273.065 197.585 285.465 199.185 ;
      LAYER met4 ;
        RECT 285.465 197.585 289.065 199.185 ;
      LAYER met4 ;
        RECT 289.065 197.585 291.465 199.185 ;
      LAYER met4 ;
        RECT 291.465 197.585 293.065 199.185 ;
      LAYER met4 ;
        RECT 293.065 197.585 301.465 199.185 ;
      LAYER met4 ;
        RECT 301.465 197.585 309.065 199.185 ;
      LAYER met4 ;
        RECT 309.065 197.585 313.465 199.185 ;
      LAYER met4 ;
        RECT 313.465 197.585 317.065 201.185 ;
      LAYER met4 ;
        RECT 259.065 195.585 265.465 197.585 ;
      LAYER met4 ;
        RECT 265.465 195.585 267.065 197.585 ;
      LAYER met4 ;
        RECT 267.065 197.185 287.465 197.585 ;
      LAYER met4 ;
        RECT 287.465 197.185 289.065 197.585 ;
      LAYER met4 ;
        RECT 289.065 197.185 303.465 197.585 ;
        RECT 267.065 195.585 275.465 197.185 ;
        RECT 259.065 195.185 275.465 195.585 ;
      LAYER met4 ;
        RECT 275.465 195.185 277.065 197.185 ;
      LAYER met4 ;
        RECT 277.065 195.185 281.465 197.185 ;
      LAYER met4 ;
        RECT 281.465 195.585 285.065 197.185 ;
      LAYER met4 ;
        RECT 285.065 195.585 287.465 197.185 ;
      LAYER met4 ;
        RECT 255.465 193.585 263.065 195.185 ;
      LAYER met4 ;
        RECT 263.065 193.585 269.465 195.185 ;
      LAYER met4 ;
        RECT 269.465 193.585 273.065 195.185 ;
      LAYER met4 ;
        RECT 273.065 193.585 275.465 195.185 ;
      LAYER met4 ;
        RECT 255.465 191.585 259.065 193.585 ;
      LAYER met4 ;
        RECT 259.065 193.185 275.465 193.585 ;
        RECT 259.065 191.585 263.465 193.185 ;
      LAYER met4 ;
        RECT 263.465 191.585 269.065 193.185 ;
      LAYER met4 ;
        RECT 269.065 191.585 275.465 193.185 ;
      LAYER met4 ;
        RECT 255.465 189.185 257.065 191.585 ;
      LAYER met4 ;
        RECT 257.065 191.185 263.465 191.585 ;
        RECT 257.065 189.585 259.465 191.185 ;
      LAYER met4 ;
        RECT 259.465 189.585 261.065 191.185 ;
      LAYER met4 ;
        RECT 261.065 189.585 263.465 191.185 ;
      LAYER met4 ;
        RECT 263.465 189.585 267.065 191.585 ;
      LAYER met4 ;
        RECT 267.065 191.185 275.465 191.585 ;
      LAYER met4 ;
        RECT 275.465 191.185 279.065 195.185 ;
      LAYER met4 ;
        RECT 267.065 189.585 269.465 191.185 ;
      LAYER met4 ;
        RECT 269.465 189.585 271.065 191.185 ;
      LAYER met4 ;
        RECT 271.065 189.585 273.465 191.185 ;
      LAYER met4 ;
        RECT 273.465 189.585 279.065 191.185 ;
      LAYER met4 ;
        RECT 279.065 189.585 281.465 195.185 ;
      LAYER met4 ;
        RECT 281.465 191.185 283.065 195.585 ;
      LAYER met4 ;
        RECT 283.065 191.585 287.465 195.585 ;
      LAYER met4 ;
        RECT 287.465 191.585 291.065 197.185 ;
      LAYER met4 ;
        RECT 291.065 191.585 293.465 197.185 ;
      LAYER met4 ;
        RECT 293.465 193.185 295.065 197.185 ;
      LAYER met4 ;
        RECT 295.065 195.185 303.465 197.185 ;
      LAYER met4 ;
        RECT 303.465 195.185 307.065 197.585 ;
      LAYER met4 ;
        RECT 307.065 197.185 315.465 197.585 ;
        RECT 295.065 193.185 299.465 195.185 ;
      LAYER met4 ;
        RECT 299.465 193.585 307.065 195.185 ;
        RECT 299.465 193.185 301.065 193.585 ;
        RECT 293.465 191.585 301.065 193.185 ;
      LAYER met4 ;
        RECT 301.065 191.585 303.465 193.585 ;
      LAYER met4 ;
        RECT 303.465 191.585 307.065 193.585 ;
      LAYER met4 ;
        RECT 307.065 191.585 309.465 197.185 ;
      LAYER met4 ;
        RECT 309.465 195.185 311.065 197.185 ;
      LAYER met4 ;
        RECT 311.065 195.185 315.465 197.185 ;
      LAYER met4 ;
        RECT 315.465 195.185 317.065 197.585 ;
        RECT 309.465 193.585 317.065 195.185 ;
      LAYER met4 ;
        RECT 283.065 191.185 297.465 191.585 ;
      LAYER met4 ;
        RECT 281.465 189.585 287.065 191.185 ;
      LAYER met4 ;
        RECT 257.065 189.185 263.465 189.585 ;
      LAYER met4 ;
        RECT 263.465 189.185 265.065 189.585 ;
      LAYER met4 ;
        RECT 265.065 189.185 273.465 189.585 ;
      LAYER met4 ;
        RECT 255.465 185.585 259.065 189.185 ;
      LAYER met4 ;
        RECT 259.065 185.585 261.465 189.185 ;
      LAYER met4 ;
        RECT 261.465 187.890 265.065 189.185 ;
        RECT 261.465 187.585 264.760 187.890 ;
        POLYGON 264.760 187.890 265.065 187.890 264.760 187.585 ;
      LAYER met4 ;
        RECT 265.065 187.585 267.465 189.185 ;
      LAYER met4 ;
        RECT 267.465 187.585 269.065 189.185 ;
      LAYER met4 ;
        RECT 269.065 187.585 273.465 189.185 ;
      LAYER met4 ;
        RECT 261.465 185.585 263.065 187.585 ;
      LAYER met4 ;
        RECT 263.065 187.185 273.465 187.585 ;
      LAYER met4 ;
        RECT 273.465 187.185 275.065 189.585 ;
      LAYER met4 ;
        RECT 275.065 187.585 277.465 189.585 ;
      LAYER met4 ;
        RECT 277.465 189.185 279.065 189.585 ;
      LAYER met4 ;
        RECT 279.065 189.185 285.465 189.585 ;
      LAYER met4 ;
        RECT 277.465 187.585 281.065 189.185 ;
      LAYER met4 ;
        RECT 281.065 187.585 285.465 189.185 ;
      LAYER met4 ;
        RECT 285.465 187.585 287.065 189.585 ;
      LAYER met4 ;
        RECT 287.065 189.185 297.465 191.185 ;
        RECT 287.065 187.585 289.465 189.185 ;
        RECT 263.065 185.585 269.465 187.185 ;
      LAYER met4 ;
        RECT 269.465 185.585 275.065 187.185 ;
      LAYER met4 ;
        RECT 275.065 185.585 279.465 187.585 ;
      LAYER met4 ;
        RECT 279.465 185.585 281.065 187.585 ;
      LAYER met4 ;
        RECT 281.065 187.185 289.465 187.585 ;
      LAYER met4 ;
        RECT 289.465 187.185 291.065 189.185 ;
      LAYER met4 ;
        RECT 291.065 187.585 293.465 189.185 ;
      LAYER met4 ;
        RECT 293.465 187.585 295.065 189.185 ;
      LAYER met4 ;
        RECT 295.065 187.585 297.465 189.185 ;
        RECT 291.065 187.185 297.465 187.585 ;
      LAYER met4 ;
        RECT 297.465 187.185 299.065 191.585 ;
      LAYER met4 ;
        RECT 299.065 189.185 303.465 191.585 ;
      LAYER met4 ;
        RECT 303.465 189.185 305.065 191.585 ;
      LAYER met4 ;
        RECT 305.065 191.185 309.465 191.585 ;
      LAYER met4 ;
        RECT 309.465 191.185 311.065 193.585 ;
      LAYER met4 ;
        RECT 311.065 191.185 315.465 193.585 ;
      LAYER met4 ;
        RECT 315.465 191.185 317.065 193.585 ;
      LAYER met4 ;
        RECT 305.065 189.585 307.465 191.185 ;
      LAYER met4 ;
        RECT 307.465 189.585 317.065 191.185 ;
      LAYER met4 ;
        RECT 305.065 189.185 309.465 189.585 ;
        RECT 299.065 187.585 301.465 189.185 ;
      LAYER met4 ;
        RECT 301.465 187.585 307.065 189.185 ;
      LAYER met4 ;
        RECT 307.065 187.585 309.465 189.185 ;
      LAYER met4 ;
        RECT 309.465 187.585 313.065 189.585 ;
      LAYER met4 ;
        RECT 313.065 187.585 315.465 189.585 ;
        RECT 281.065 185.585 287.465 187.185 ;
      LAYER met4 ;
        RECT 287.465 185.585 293.065 187.185 ;
      LAYER met4 ;
        RECT 293.065 185.585 295.465 187.185 ;
      LAYER met4 ;
        RECT 255.465 183.185 257.065 185.585 ;
      LAYER met4 ;
        RECT 257.065 185.185 273.465 185.585 ;
      LAYER met4 ;
        RECT 273.465 185.185 275.065 185.585 ;
      LAYER met4 ;
        RECT 275.065 185.185 287.465 185.585 ;
        RECT 257.065 183.185 259.465 185.185 ;
      LAYER met4 ;
        RECT 259.465 183.185 261.065 185.185 ;
      LAYER met4 ;
        RECT 261.065 183.185 263.465 185.185 ;
      LAYER met4 ;
        RECT 263.465 183.185 265.065 185.185 ;
      LAYER met4 ;
        RECT 265.065 183.185 273.465 185.185 ;
      LAYER met4 ;
        RECT 273.465 183.585 277.065 185.185 ;
      LAYER met4 ;
        RECT 277.065 183.585 283.465 185.185 ;
      LAYER met4 ;
        RECT 255.465 181.585 265.065 183.185 ;
      LAYER met4 ;
        RECT 265.065 181.585 267.465 183.185 ;
      LAYER met4 ;
        RECT 267.465 181.585 271.065 183.185 ;
      LAYER met4 ;
        RECT 271.065 181.585 273.465 183.185 ;
      LAYER met4 ;
        RECT 255.465 179.185 257.065 181.585 ;
      LAYER met4 ;
        RECT 257.065 179.185 259.465 181.585 ;
      LAYER met4 ;
        RECT 259.465 179.185 265.065 181.585 ;
      LAYER met4 ;
        RECT 265.065 181.185 273.465 181.585 ;
      LAYER met4 ;
        RECT 273.465 181.185 275.065 183.585 ;
      LAYER met4 ;
        RECT 275.065 183.185 283.465 183.585 ;
        RECT 275.065 181.185 279.465 183.185 ;
      LAYER met4 ;
        RECT 279.465 181.185 281.065 183.185 ;
      LAYER met4 ;
        RECT 281.065 181.185 283.465 183.185 ;
      LAYER met4 ;
        RECT 283.465 181.185 285.065 185.185 ;
      LAYER met4 ;
        RECT 285.065 183.585 287.465 185.185 ;
      LAYER met4 ;
        RECT 287.465 183.585 289.065 185.585 ;
      LAYER met4 ;
        RECT 289.065 183.585 295.465 185.585 ;
      LAYER met4 ;
        RECT 295.465 185.185 299.065 187.185 ;
      LAYER met4 ;
        RECT 299.065 185.585 303.465 187.585 ;
      LAYER met4 ;
        RECT 303.465 185.585 307.065 187.585 ;
      LAYER met4 ;
        RECT 307.065 185.585 315.465 187.585 ;
        RECT 299.065 185.185 315.465 185.585 ;
      LAYER met4 ;
        RECT 295.465 183.585 303.065 185.185 ;
      LAYER met4 ;
        RECT 303.065 183.585 307.465 185.185 ;
        RECT 285.065 183.185 299.465 183.585 ;
        RECT 285.065 181.585 293.465 183.185 ;
      LAYER met4 ;
        RECT 293.465 181.585 295.065 183.185 ;
      LAYER met4 ;
        RECT 295.065 181.585 299.465 183.185 ;
      LAYER met4 ;
        RECT 299.465 181.585 301.065 183.585 ;
      LAYER met4 ;
        RECT 301.065 183.185 307.465 183.585 ;
      LAYER met4 ;
        RECT 307.465 183.185 311.065 185.185 ;
      LAYER met4 ;
        RECT 311.065 183.185 315.465 185.185 ;
      LAYER met4 ;
        RECT 315.465 183.185 317.065 189.585 ;
      LAYER met4 ;
        RECT 301.065 181.585 303.465 183.185 ;
      LAYER met4 ;
        RECT 303.465 181.585 305.065 183.185 ;
      LAYER met4 ;
        RECT 305.065 181.585 307.465 183.185 ;
      LAYER met4 ;
        RECT 307.465 181.585 317.065 183.185 ;
      LAYER met4 ;
        RECT 285.065 181.185 307.465 181.585 ;
        RECT 265.065 179.185 271.465 181.185 ;
      LAYER met4 ;
        RECT 271.465 179.585 275.065 181.185 ;
      LAYER met4 ;
        RECT 275.065 179.585 277.465 181.185 ;
      LAYER met4 ;
        RECT 277.465 179.890 293.065 181.185 ;
      LAYER met4 ;
        POLYGON 277.465 179.890 277.770 179.585 277.465 179.585 ;
      LAYER met4 ;
        RECT 277.770 179.585 293.065 179.890 ;
        RECT 271.465 179.185 273.065 179.585 ;
        RECT 255.465 177.585 273.065 179.185 ;
        RECT 255.465 163.185 257.065 177.585 ;
      LAYER met4 ;
        RECT 257.065 175.185 271.465 177.585 ;
      LAYER met4 ;
        RECT 271.465 175.185 273.065 177.585 ;
      LAYER met4 ;
        RECT 273.065 177.185 281.465 179.585 ;
      LAYER met4 ;
        RECT 281.465 177.185 285.065 179.585 ;
      LAYER met4 ;
        RECT 285.065 177.185 287.465 179.585 ;
      LAYER met4 ;
        RECT 287.465 179.185 293.065 179.585 ;
      LAYER met4 ;
        RECT 293.065 179.185 307.465 181.185 ;
      LAYER met4 ;
        RECT 287.465 177.585 295.065 179.185 ;
        RECT 287.465 177.185 289.065 177.585 ;
      LAYER met4 ;
        RECT 273.065 175.585 277.465 177.185 ;
      LAYER met4 ;
        RECT 277.465 175.585 289.065 177.185 ;
      LAYER met4 ;
        RECT 289.065 175.585 293.465 177.585 ;
      LAYER met4 ;
        RECT 293.465 177.185 295.065 177.585 ;
      LAYER met4 ;
        RECT 295.065 177.185 299.465 179.185 ;
      LAYER met4 ;
        RECT 299.465 177.585 305.065 179.185 ;
      LAYER met4 ;
        RECT 305.065 177.585 307.465 179.185 ;
      LAYER met4 ;
        RECT 307.465 177.585 309.065 181.585 ;
      LAYER met4 ;
        RECT 309.065 177.585 315.465 181.585 ;
      LAYER met4 ;
        RECT 293.465 175.585 297.065 177.185 ;
      LAYER met4 ;
        RECT 273.065 175.185 279.465 175.585 ;
        RECT 257.065 165.585 259.465 175.185 ;
      LAYER met4 ;
        RECT 259.465 173.585 269.065 175.185 ;
        RECT 259.465 167.185 261.065 173.585 ;
      LAYER met4 ;
        RECT 261.065 167.185 267.465 173.585 ;
      LAYER met4 ;
        RECT 267.465 167.185 269.065 173.585 ;
        RECT 259.465 165.585 269.065 167.185 ;
      LAYER met4 ;
        RECT 269.065 165.585 271.465 175.185 ;
      LAYER met4 ;
        RECT 271.465 173.585 277.065 175.185 ;
      LAYER met4 ;
        RECT 277.065 173.585 279.465 175.185 ;
      LAYER met4 ;
        RECT 279.465 173.585 285.065 175.585 ;
      LAYER met4 ;
        RECT 285.065 175.185 295.465 175.585 ;
      LAYER met4 ;
        RECT 271.465 171.585 275.065 173.585 ;
      LAYER met4 ;
        RECT 275.065 173.185 279.465 173.585 ;
      LAYER met4 ;
        RECT 279.465 173.185 281.065 173.585 ;
      LAYER met4 ;
        RECT 275.065 171.585 277.465 173.185 ;
      LAYER met4 ;
        RECT 277.465 171.585 281.065 173.185 ;
      LAYER met4 ;
        RECT 281.065 171.585 283.465 173.585 ;
      LAYER met4 ;
        RECT 283.465 173.185 285.065 173.585 ;
      LAYER met4 ;
        RECT 285.065 173.185 289.465 175.185 ;
      LAYER met4 ;
        RECT 289.465 173.585 293.065 175.185 ;
      LAYER met4 ;
        RECT 293.065 173.585 295.465 175.185 ;
      LAYER met4 ;
        RECT 289.465 173.185 291.065 173.585 ;
      LAYER met4 ;
        RECT 291.065 173.185 295.465 173.585 ;
      LAYER met4 ;
        RECT 295.465 173.185 297.065 175.585 ;
      LAYER met4 ;
        RECT 297.065 173.585 299.465 177.185 ;
      LAYER met4 ;
        RECT 299.465 175.185 301.065 177.585 ;
      LAYER met4 ;
        RECT 301.065 175.185 303.465 177.585 ;
      LAYER met4 ;
        RECT 303.465 175.185 305.065 177.585 ;
      LAYER met4 ;
        RECT 305.065 177.185 315.465 177.585 ;
      LAYER met4 ;
        RECT 315.465 177.185 317.065 181.585 ;
      LAYER met4 ;
        RECT 305.065 175.585 309.465 177.185 ;
      LAYER met4 ;
        RECT 309.465 175.585 311.065 177.185 ;
      LAYER met4 ;
        RECT 311.065 175.585 313.465 177.185 ;
        RECT 305.065 175.185 313.465 175.585 ;
      LAYER met4 ;
        RECT 313.465 175.185 317.065 177.185 ;
        RECT 299.465 173.585 305.065 175.185 ;
      LAYER met4 ;
        RECT 305.065 173.585 307.465 175.185 ;
      LAYER met4 ;
        RECT 283.465 171.585 291.065 173.185 ;
      LAYER met4 ;
        RECT 291.065 171.585 293.465 173.185 ;
      LAYER met4 ;
        RECT 293.465 171.890 297.065 173.185 ;
      LAYER met4 ;
        POLYGON 293.465 171.890 293.770 171.585 293.465 171.585 ;
      LAYER met4 ;
        RECT 293.770 171.585 297.065 171.890 ;
        RECT 271.465 169.185 273.065 171.585 ;
      LAYER met4 ;
        RECT 273.065 171.185 283.465 171.585 ;
        RECT 273.065 169.585 275.465 171.185 ;
      LAYER met4 ;
        RECT 275.465 169.585 277.065 171.185 ;
      LAYER met4 ;
        RECT 277.065 169.585 283.465 171.185 ;
        RECT 273.065 169.185 283.465 169.585 ;
      LAYER met4 ;
        RECT 271.465 167.585 275.065 169.185 ;
      LAYER met4 ;
        RECT 275.065 167.585 279.465 169.185 ;
        RECT 257.065 163.185 271.465 165.585 ;
      LAYER met4 ;
        RECT 271.465 163.185 273.065 167.585 ;
      LAYER met4 ;
        RECT 273.065 167.185 279.465 167.585 ;
      LAYER met4 ;
        RECT 279.465 167.185 281.065 169.185 ;
      LAYER met4 ;
        RECT 281.065 167.585 283.465 169.185 ;
      LAYER met4 ;
        RECT 283.465 167.585 289.065 171.585 ;
      LAYER met4 ;
        RECT 289.065 169.585 295.465 171.585 ;
      LAYER met4 ;
        RECT 295.465 171.185 297.065 171.585 ;
      LAYER met4 ;
        RECT 297.065 171.185 307.465 173.585 ;
      LAYER met4 ;
        RECT 307.465 173.185 309.065 175.185 ;
      LAYER met4 ;
        RECT 309.065 173.585 311.465 175.185 ;
      LAYER met4 ;
        RECT 311.465 173.585 317.065 175.185 ;
      LAYER met4 ;
        RECT 309.065 173.185 315.465 173.585 ;
      LAYER met4 ;
        RECT 295.465 169.585 301.065 171.185 ;
      LAYER met4 ;
        RECT 301.065 169.585 307.465 171.185 ;
      LAYER met4 ;
        RECT 307.465 169.585 311.065 173.185 ;
      LAYER met4 ;
        RECT 311.065 171.185 315.465 173.185 ;
      LAYER met4 ;
        RECT 315.465 171.185 317.065 173.585 ;
      LAYER met4 ;
        RECT 311.065 169.585 313.465 171.185 ;
      LAYER met4 ;
        RECT 313.465 169.585 317.065 171.185 ;
      LAYER met4 ;
        RECT 289.065 169.185 297.465 169.585 ;
        RECT 289.065 167.585 293.465 169.185 ;
        RECT 273.065 165.585 275.465 167.185 ;
      LAYER met4 ;
        RECT 275.465 165.585 281.065 167.185 ;
      LAYER met4 ;
        RECT 281.065 165.585 293.465 167.585 ;
      LAYER met4 ;
        RECT 293.465 167.185 295.065 169.185 ;
      LAYER met4 ;
        RECT 295.065 167.585 297.465 169.185 ;
      LAYER met4 ;
        RECT 297.465 167.585 299.065 169.585 ;
      LAYER met4 ;
        RECT 299.065 169.185 315.465 169.585 ;
        RECT 299.065 167.585 301.465 169.185 ;
        RECT 295.065 167.185 301.465 167.585 ;
        RECT 273.065 163.185 277.465 165.585 ;
      LAYER met4 ;
        RECT 277.465 163.185 279.065 165.585 ;
      LAYER met4 ;
        RECT 279.065 165.185 293.465 165.585 ;
        RECT 279.065 163.185 281.465 165.185 ;
      LAYER met4 ;
        RECT 281.465 163.185 283.065 165.185 ;
      LAYER met4 ;
        RECT 283.065 163.185 287.465 165.185 ;
      LAYER met4 ;
        RECT 287.465 163.185 289.065 165.185 ;
      LAYER met4 ;
        RECT 289.065 163.185 293.465 165.185 ;
      LAYER met4 ;
        RECT 293.465 163.185 297.065 167.185 ;
      LAYER met4 ;
        RECT 297.065 165.585 301.465 167.185 ;
      LAYER met4 ;
        RECT 301.465 165.585 305.065 169.185 ;
      LAYER met4 ;
        RECT 305.065 167.585 311.465 169.185 ;
      LAYER met4 ;
        RECT 311.465 167.585 313.065 169.185 ;
      LAYER met4 ;
        RECT 313.065 167.585 315.465 169.185 ;
        RECT 305.065 167.185 315.465 167.585 ;
      LAYER met4 ;
        RECT 315.465 167.185 317.065 169.585 ;
      LAYER met4 ;
        RECT 305.065 165.585 307.465 167.185 ;
      LAYER met4 ;
        RECT 307.465 165.585 311.065 167.185 ;
      LAYER met4 ;
        RECT 297.065 165.185 309.465 165.585 ;
        RECT 297.065 163.185 305.465 165.185 ;
      LAYER met4 ;
        RECT 305.465 163.185 307.065 165.185 ;
      LAYER met4 ;
        RECT 307.065 163.185 309.465 165.185 ;
      LAYER met4 ;
        RECT 309.465 163.185 311.065 165.585 ;
      LAYER met4 ;
        RECT 311.065 163.185 313.465 167.185 ;
      LAYER met4 ;
        RECT 313.465 163.185 317.065 167.185 ;
        RECT 255.465 161.585 317.065 163.185 ;
      LAYER met4 ;
        RECT 100.115 96.415 132.145 98.015 ;
        RECT 97.165 93.265 124.815 94.865 ;
        RECT 43.135 78.605 52.745 82.655 ;
        RECT 56.135 78.605 65.745 82.655 ;
        RECT 69.135 78.605 78.745 82.655 ;
        RECT 82.135 78.605 91.745 82.655 ;
        RECT 95.135 78.605 104.745 82.655 ;
        RECT 130.545 78.605 132.145 96.415 ;
        RECT 38.470 77.005 132.145 78.605 ;
        RECT 38.470 63.590 39.745 77.005 ;
        RECT 43.135 73.045 52.745 77.005 ;
        RECT 56.135 73.045 65.745 77.005 ;
        RECT 69.135 73.045 78.745 77.005 ;
        RECT 82.135 73.045 91.745 77.005 ;
        RECT 95.135 73.045 104.745 77.005 ;
        RECT 42.800 71.180 108.800 71.690 ;
        RECT 133.525 71.180 135.125 110.315 ;
        RECT 42.800 69.580 135.125 71.180 ;
        RECT 42.800 69.190 108.800 69.580 ;
        RECT 43.135 63.590 52.745 67.835 ;
        RECT 56.135 63.590 65.745 67.835 ;
        RECT 69.135 63.590 78.745 67.835 ;
        RECT 82.135 63.590 91.745 67.835 ;
        RECT 95.135 63.590 104.745 67.835 ;
        RECT 38.470 61.990 104.745 63.590 ;
        RECT 43.135 58.225 52.745 61.990 ;
        RECT 56.135 58.225 65.745 61.990 ;
        RECT 69.135 58.225 78.745 61.990 ;
        RECT 82.135 58.225 91.745 61.990 ;
        RECT 95.135 58.225 104.745 61.990 ;
        RECT 12.915 45.565 92.315 47.165 ;
        RECT 65.765 42.615 117.715 44.215 ;
        RECT 68.865 40.015 120.815 41.615 ;
        RECT 72.095 9.265 82.535 10.865 ;
        RECT 153.565 8.890 156.765 113.350 ;
        RECT 179.925 110.505 293.305 113.705 ;
        RECT 174.350 101.160 174.680 101.490 ;
        RECT 174.365 62.730 174.665 101.160 ;
        RECT 174.350 62.400 174.680 62.730 ;
        RECT 179.925 13.705 181.525 110.505 ;
        RECT 186.310 104.560 186.640 104.890 ;
        RECT 186.325 55.930 186.625 104.560 ;
        RECT 186.310 55.600 186.640 55.930 ;
        RECT 198.555 8.890 200.155 106.665 ;
        RECT 208.390 99.800 208.720 100.130 ;
        RECT 208.405 87.210 208.705 99.800 ;
        RECT 208.390 86.880 208.720 87.210 ;
        RECT 217.185 13.705 218.785 110.505 ;
        RECT 229.550 101.160 229.880 101.490 ;
        RECT 221.270 94.360 221.600 94.690 ;
        RECT 227.710 94.360 228.040 94.690 ;
        RECT 221.285 92.650 221.585 94.360 ;
        RECT 221.270 92.320 221.600 92.650 ;
        RECT 227.725 62.050 228.025 94.360 ;
        RECT 229.565 70.210 229.865 101.160 ;
        RECT 229.550 69.880 229.880 70.210 ;
        RECT 227.710 61.720 228.040 62.050 ;
        RECT 235.815 8.890 237.415 106.665 ;
        RECT 238.750 101.840 239.080 102.170 ;
        RECT 238.765 38.930 239.065 101.840 ;
        RECT 246.110 79.400 246.440 79.730 ;
        RECT 246.125 72.250 246.425 79.400 ;
        RECT 246.110 71.920 246.440 72.250 ;
        RECT 238.750 38.600 239.080 38.930 ;
        RECT 254.445 13.705 256.045 110.505 ;
        RECT 259.910 101.160 260.240 101.490 ;
        RECT 259.925 73.610 260.225 101.160 ;
        RECT 260.830 97.080 261.160 97.410 ;
        RECT 260.845 87.890 261.145 97.080 ;
        RECT 260.830 87.560 261.160 87.890 ;
        RECT 259.910 73.280 260.240 73.610 ;
        RECT 273.075 8.890 274.675 106.665 ;
        RECT 277.390 101.160 277.720 101.490 ;
        RECT 277.405 70.210 277.705 101.160 ;
        RECT 277.390 69.880 277.720 70.210 ;
        RECT 291.705 13.705 293.305 110.505 ;
        RECT 310.335 8.890 311.935 106.665 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.160 5.690 311.935 8.890 ;
        RECT 97.530 1.000 98.430 2.125 ;
        RECT 116.850 1.750 132.465 2.650 ;
        RECT 136.170 1.750 152.360 2.650 ;
        RECT 116.850 1.000 117.750 1.750 ;
        RECT 136.170 1.000 137.070 1.750 ;
  END
END tt_um_cw_vref
END LIBRARY

