VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_simon
  CLASS BLOCK ;
  FOREIGN tt_um_urish_simon ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.450 2.480 62.050 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.320 2.480 100.920 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.190 2.480 139.790 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.150 2.480 58.750 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.020 2.480 97.620 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.890 2.480 136.490 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 110.520 144.130 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 110.520 146.890 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 141.070 110.520 141.370 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 138.310 110.520 138.610 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 110.520 135.850 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 110.520 133.090 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 110.520 130.330 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 127.270 110.520 127.570 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 110.520 124.810 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 110.520 122.050 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 118.990 110.520 119.290 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 110.520 116.530 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 110.520 113.770 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 110.520 111.010 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 110.520 108.250 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 110.520 105.490 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 110.520 102.730 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 110.520 99.970 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 110.520 97.210 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 110.520 50.290 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 110.520 47.530 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 110.520 44.770 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 110.520 42.010 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 110.520 39.250 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 110.520 36.490 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 110.520 33.730 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 110.520 30.970 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 110.520 72.370 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 110.520 69.610 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 110.520 66.850 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 110.520 64.090 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.030 110.520 61.330 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 58.270 110.520 58.570 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 110.520 55.810 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 110.520 53.050 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 110.520 94.450 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 110.520 91.690 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 110.520 88.930 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 110.520 86.170 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 110.520 83.410 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 110.520 80.650 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 110.520 77.890 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 110.520 75.130 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 2.635 158.430 108.990 ;
      LAYER li1 ;
        RECT 2.760 2.635 158.240 108.885 ;
      LAYER met1 ;
        RECT 2.760 1.060 158.540 110.120 ;
      LAYER met2 ;
        RECT 3.780 1.030 156.760 110.685 ;
      LAYER met3 ;
        RECT 6.505 2.555 156.335 110.665 ;
      LAYER met4 ;
        RECT 31.370 110.120 33.030 110.665 ;
        RECT 34.130 110.120 35.790 110.665 ;
        RECT 36.890 110.120 38.550 110.665 ;
        RECT 39.650 110.120 41.310 110.665 ;
        RECT 42.410 110.120 44.070 110.665 ;
        RECT 45.170 110.120 46.830 110.665 ;
        RECT 47.930 110.120 49.590 110.665 ;
        RECT 50.690 110.120 52.350 110.665 ;
        RECT 53.450 110.120 55.110 110.665 ;
        RECT 56.210 110.120 57.870 110.665 ;
        RECT 58.970 110.120 60.630 110.665 ;
        RECT 61.730 110.120 63.390 110.665 ;
        RECT 64.490 110.120 66.150 110.665 ;
        RECT 67.250 110.120 68.910 110.665 ;
        RECT 70.010 110.120 71.670 110.665 ;
        RECT 72.770 110.120 74.430 110.665 ;
        RECT 75.530 110.120 77.190 110.665 ;
        RECT 78.290 110.120 79.950 110.665 ;
        RECT 81.050 110.120 82.710 110.665 ;
        RECT 83.810 110.120 85.470 110.665 ;
        RECT 86.570 110.120 88.230 110.665 ;
        RECT 89.330 110.120 90.990 110.665 ;
        RECT 92.090 110.120 93.750 110.665 ;
        RECT 94.850 110.120 96.510 110.665 ;
        RECT 97.610 110.120 99.270 110.665 ;
        RECT 100.370 110.120 102.030 110.665 ;
        RECT 103.130 110.120 104.790 110.665 ;
        RECT 105.890 110.120 107.550 110.665 ;
        RECT 108.650 110.120 110.310 110.665 ;
        RECT 111.410 110.120 113.070 110.665 ;
        RECT 114.170 110.120 115.830 110.665 ;
        RECT 116.930 110.120 118.590 110.665 ;
        RECT 119.690 110.120 121.350 110.665 ;
        RECT 122.450 110.120 124.110 110.665 ;
        RECT 125.210 110.120 126.870 110.665 ;
        RECT 127.970 110.120 129.630 110.665 ;
        RECT 130.730 110.120 132.390 110.665 ;
        RECT 133.490 110.120 135.150 110.665 ;
        RECT 136.250 110.120 137.910 110.665 ;
        RECT 139.010 110.120 140.670 110.665 ;
        RECT 141.770 110.120 143.430 110.665 ;
        RECT 144.530 110.120 146.190 110.665 ;
        RECT 147.290 110.120 148.745 110.665 ;
        RECT 30.655 109.440 148.745 110.120 ;
        RECT 30.655 18.535 56.750 109.440 ;
        RECT 59.150 18.535 60.050 109.440 ;
        RECT 62.450 18.535 95.620 109.440 ;
        RECT 98.020 18.535 98.920 109.440 ;
        RECT 101.320 18.535 134.490 109.440 ;
        RECT 136.890 18.535 137.790 109.440 ;
        RECT 140.190 18.535 148.745 109.440 ;
  END
END tt_um_urish_simon
END LIBRARY

